`timescale 1ns / 1ps
module test;
reg clk, rst;
reg in_valid;
reg [15:0] in_index;
wire out_valid;
wire [15:0] out_index;
initial begin
clk = 1'b1;
rst = 1'b1;
in_valid = 0;
in_index = 0;
#1
rst = 1'b0;
#1
rst = 1'b1;
#1
in_valid = 1;
end
always #5 clk = ~clk;
always @ (posedge clk) begin
    if (in_valid == 1) begin
        if (in_index < 1440 - 4)
       in_index <= in_index + 4;
        else
        in_valid <= 0;
    end
end
wire [1440 * 10 - 1: 0] L = {10'd21, 10'd42, -10'd48, 10'd43, 10'd9, 10'd26, -10'd25, 10'd38, 10'd35, 10'd47, 10'd50, 10'd6, -10'd19, -10'd40, -10'd38, 10'd42, -10'd51, -10'd35, 10'd29, 10'd15, 10'd22, 10'd31, 10'd31, -10'd48, -10'd40, -10'd59, -10'd43, -10'd40, -10'd6, 10'd52, -10'd34, -10'd10, 10'd26, 10'd10, 10'd29, -10'd41, -10'd11, 10'd77, -10'd14, -10'd11, -10'd26, 10'd57, -10'd34, 10'd16, -10'd13, -10'd17, 10'd45, 10'd41, 10'd15, -10'd8, -10'd28, -10'd46, 10'd12, 10'd26, -10'd50, 10'd42, -10'd61, 10'd28, 10'd39, -10'd53, 10'd45, -10'd31, -10'd39, 10'd54, -10'd49, -10'd62, -10'd27, 10'd52, -10'd23, -10'd14, 10'd43, 10'd24, 10'd42, 10'd83, -10'd53, 10'd27, 10'd21, -10'd50, -10'd24, 10'd39, -10'd29, 10'd8, 10'd22, -10'd34, 10'd26, -10'd31, 10'd2, -10'd38, -10'd19, -10'd38, 10'd58, 10'd49, 10'd42, -10'd12, -10'd29, 10'd24, 10'd25, 10'd24, 10'd62, -10'd44, 10'd51, 10'd24, 10'd35, -10'd19, -10'd46, -10'd43, 10'd59, -10'd41, -10'd33, 10'd57, -10'd28, -10'd102, -10'd45, 10'd14, -10'd55, -10'd31, -10'd17, 10'd76, -10'd30, -10'd57, -10'd45, -10'd35, 10'd54, 10'd56, -10'd32, -10'd35, 10'd45, 10'd27, -10'd49, 10'd43, -10'd68, 10'd14, 10'd46, -10'd37, 10'd32, -10'd56, -10'd39, -10'd20, 10'd36, -10'd25, -10'd55, 10'd19, -10'd46, -10'd19, -10'd47, 10'd11, 10'd47, 10'd23, 10'd41, -10'd26, -10'd34, 10'd41, -10'd62, -10'd36, -10'd41, 10'd55, -10'd35, -10'd23, 10'd33, -10'd5, 10'd35, -10'd14, 10'd47, -10'd47, 10'd19, -10'd19, -10'd20, -10'd1, 10'd25, 10'd46, 10'd53, 10'd29, -10'd10, -10'd45, -10'd68, 10'd24, 10'd42, -10'd41, -10'd16, 10'd41, -10'd30, -10'd31, -10'd38, -10'd45, 10'd38, 10'd67, -10'd46, -10'd53, 10'd21, -10'd54, -10'd42, -10'd36, 10'd43, 10'd29, -10'd45, -10'd33, -10'd59, 10'd27, 10'd64, 10'd34, -10'd56, -10'd27, 10'd45, 10'd13, -10'd27, -10'd22, -10'd56, -10'd72, 10'd46, -10'd50, 10'd31, -10'd33, 10'd56, -10'd30, -10'd38, 10'd28, 10'd59, -10'd52, -10'd63, -10'd46, -10'd30, 10'd28, -10'd8, 10'd16, -10'd43, -10'd5, 10'd46, -10'd37, 10'd50, -10'd43, -10'd58, -10'd13, 10'd29, 10'd45, 10'd22, -10'd16, -10'd16, -10'd51, 10'd52, 10'd61, 10'd18, 10'd33, 10'd69, -10'd54, -10'd68, -10'd50, 10'd40, -10'd37, -10'd30, -10'd63, 10'd54, -10'd32, -10'd59, -10'd11, 10'd78, -10'd27, 10'd35, 10'd54, 10'd1, 10'd38, 10'd20, 10'd67, 10'd23, -10'd29, 10'd11, 10'd29, -10'd16, 10'd38, -10'd41, 10'd6, -10'd22, 10'd16, 10'd17, 10'd35, 10'd46, 10'd46, -10'd52, 10'd59, 10'd54, -10'd29, 10'd9, -10'd65, -10'd29, -10'd30, -10'd68, -10'd53, -10'd14, -10'd20, -10'd3, 10'd29, 10'd55, 10'd43, -10'd40, -10'd44, 10'd27, -10'd43, -10'd44, 10'd25, 10'd14, -10'd48, -10'd58, 10'd71, 10'd44, -10'd26, 10'd28, -10'd35, -10'd21, 10'd27, -10'd24, -10'd1, 10'd42, -10'd46, -10'd56, -10'd59, 10'd27, -10'd43, 10'd63, 10'd28, -10'd71, -10'd43, 10'd39, 10'd81, 10'd18, -10'd4, -10'd57, 10'd59, -10'd6, -10'd28, 10'd38, -10'd37, 10'd25, -10'd47, -10'd36, -10'd34, -10'd13, 10'd32, -10'd42, 10'd38, -10'd37, -10'd76, -10'd41, -10'd32, 10'd30, 10'd38, 10'd76, -10'd13, -10'd23, -10'd22, -10'd16, 10'd40, 10'd68, -10'd31, 10'd25, 10'd16, 10'd68, -10'd37, 10'd36, 10'd28, 10'd38, 10'd53, 10'd2, -10'd35, 10'd36, 10'd51, -10'd45, 10'd70, 10'd33, 10'd28, -10'd34, -10'd51, 10'd44, 10'd24, 10'd23, -10'd42, 10'd28, 10'd4, -10'd13, 10'd22, 10'd43, 10'd44, 10'd9, -10'd36, 10'd39, -10'd46, 10'd49, 10'd44, -10'd20, -10'd62, -10'd20, 10'd23, 10'd35, 10'd22, 10'd42, -10'd19, 10'd42, 10'd42, -10'd60, 10'd7, 10'd29, -10'd47, 10'd12, -10'd22, -10'd24, -10'd25, 10'd40, 10'd55, 10'd41, -10'd46, -10'd22, 10'd63, 10'd26, 10'd39, -10'd41, 10'd13, 10'd47, -10'd38, -10'd67, -10'd31, -10'd33, -10'd70, 10'd50, -10'd38, 10'd38, -10'd55, -10'd18, -10'd48, -10'd42, 10'd7, 10'd68, 10'd15, 10'd48, -10'd30, 10'd65, -10'd23, 10'd54, -10'd63, 10'd34, 10'd45, -10'd49, -10'd47, -10'd7, 10'd22, -10'd20, -10'd31, 10'd58, 10'd53, -10'd35, -10'd38, 10'd50, -10'd29, -10'd37, 10'd21, 10'd29, -10'd70, 10'd29, -10'd61, 10'd42, 10'd48, 10'd45, -10'd41, 10'd53, 10'd43, 10'd36, 10'd56, -10'd11, -10'd56, -10'd20, 10'd29, -10'd22, 10'd52, -10'd35, -10'd45, 10'd64, -10'd58, -10'd12, -10'd48, 10'd30, -10'd48, -10'd25, 10'd39, 10'd29, 10'd40, -10'd29, 10'd20, -10'd55, 10'd35, 10'd52, 10'd16, 10'd21, 10'd64, -10'd34, 10'd24, 10'd55, -10'd31, -10'd55, -10'd19, 10'd30, -10'd10, 10'd43, 10'd54, 10'd12, 10'd41, -10'd46, 10'd18, 10'd41, -10'd63, -10'd53, 10'd2, -10'd33, 10'd43, -10'd45, -10'd15, 10'd56, 10'd28, 10'd63, -10'd40, -10'd27, -10'd34, -10'd12, 10'd10, 10'd30, -10'd61, -10'd27, 10'd13, -10'd39, -10'd34, 10'd32, 10'd30, 10'd56, -10'd28, -10'd37, -10'd16, -10'd45, 10'd42, -10'd31, 10'd57, 10'd48, -10'd46, -10'd32, 10'd37, 10'd21, 10'd52, -10'd32, -10'd79, 10'd6, 10'd55, 10'd24, -10'd29, -10'd32, -10'd35, 10'd60, 10'd22, -10'd45, -10'd20, -10'd11, -10'd48, 10'd32, 10'd64, -10'd34, -10'd46, 10'd35, -10'd46, 10'd43, -10'd29, 10'd31, -10'd13, -10'd8, -10'd19, -10'd43, 10'd37, 10'd34, -10'd40, -10'd64, 10'd31, 10'd38, 10'd55, -10'd60, -10'd23, -10'd27, -10'd46, -10'd41, -10'd33, -10'd47, 10'd51, 10'd45, -10'd42, 10'd36, -10'd19, 10'd7, 10'd30, -10'd0, 10'd22, -10'd48, -10'd45, -10'd13, 10'd35, -10'd22, -10'd56, 10'd45, 10'd27, 10'd60, -10'd66, 10'd52, -10'd52, -10'd69, -10'd31, -10'd47, 10'd54, -10'd36, -10'd42, 10'd30, -10'd0, 10'd58, -10'd27, -10'd18, -10'd28, 10'd46, -10'd55, 10'd2, 10'd20, -10'd18, -10'd50, 10'd43, 10'd50, 10'd5, 10'd6, -10'd20, -10'd50, 10'd31, -10'd57, 10'd23, -10'd28, 10'd17, 10'd19, 10'd47, -10'd13, -10'd53, 10'd26, 10'd35, 10'd32, 10'd17, -10'd14, 10'd52, 10'd42, 10'd50, -10'd28, -10'd20, 10'd65, 10'd76, 10'd29, 10'd13, -10'd37, -10'd49, 10'd35, -10'd28, 10'd40, 10'd46, -10'd54, -10'd36, 10'd26, -10'd17, -10'd42, -10'd41, 10'd37, -10'd31, 10'd56, -10'd35, -10'd43, 10'd53, -10'd27, 10'd27, -10'd54, -10'd35, 10'd77, 10'd44, 10'd30, 10'd8, -10'd56, -10'd74, 10'd41, -10'd50, -10'd52, 10'd38, 10'd48, 10'd46, -10'd34, -10'd45, 10'd33, -10'd50, -10'd20, -10'd56, -10'd46, 10'd69, -10'd4, 10'd40, 10'd70, -10'd30, 10'd42, -10'd78, 10'd68, -10'd35, 10'd68, 10'd32, -10'd20, -10'd47, 10'd28, -10'd44, -10'd48, 10'd62, 10'd31, 10'd57, -10'd23, 10'd30, 10'd27, 10'd38, 10'd63, -10'd2, -10'd16, -10'd18, 10'd58, 10'd54, 10'd48, -10'd43, -10'd72, -10'd40, 10'd53, -10'd43, 10'd42, -10'd53, 10'd15, -10'd41, -10'd5, 10'd35, -10'd1, 10'd25, 10'd39, -10'd42, -10'd7, 10'd30, -10'd59, 10'd21, 10'd42, 10'd24, 10'd29, 10'd49, 10'd41, -10'd6, 10'd32, -10'd33, -10'd48, 10'd54, 10'd35, 10'd63, 10'd48, 10'd24, -10'd38, 10'd20, 10'd44, -10'd14, -10'd25, -10'd35, 10'd73, 10'd43, 10'd33, 10'd15, -10'd33, 10'd65, -10'd44, 10'd39, -10'd54, 10'd50, 10'd42, 10'd26, 10'd39, -10'd5, 10'd11, -10'd42, -10'd42, 10'd44, 10'd37, 10'd3, -10'd48, -10'd6, 10'd27, 10'd29, 10'd9, -10'd13, 10'd57, 10'd29, -10'd11, 10'd30, -10'd39, 10'd18, 10'd25, 10'd60, 10'd62, -10'd53, 10'd32, -10'd79, -10'd64, 10'd41, 10'd14, 10'd38, -10'd50, 10'd31, -10'd31, -10'd56, -10'd54, 10'd37, -10'd14, 10'd55, 10'd24, -10'd38, -10'd35, 10'd29, 10'd41, 10'd47, 10'd29, 10'd34, 10'd43, -10'd0, -10'd40, -10'd59, 10'd12, -10'd54, -10'd35, -10'd25, -10'd85, -10'd59, 10'd0, 10'd12, -10'd79, -10'd8, 10'd10, -10'd48, -10'd49, -10'd42, -10'd24, 10'd27, -10'd13, -10'd49, -10'd26, 10'd37, -10'd59, -10'd35, 10'd11, -10'd11, 10'd47, 10'd55, -10'd28, -10'd48, 10'd34, 10'd40, -10'd25, 10'd20, 10'd55, -10'd63, -10'd20, -10'd36, -10'd34, 10'd90, 10'd42, -10'd46, -10'd33, -10'd37, 10'd53, 10'd46, -10'd16, -10'd27, 10'd57, -10'd39, 10'd35, 10'd23, -10'd26, -10'd35, 10'd23, -10'd24, 10'd42, 10'd48, -10'd22, -10'd26, 10'd48, 10'd53, -10'd15, -10'd51, -10'd39, -10'd41, 10'd47, -10'd42, 10'd30, 10'd43, -10'd3, 10'd51, 10'd5, -10'd45, 10'd25, 10'd5, -10'd41, -10'd31, 10'd30, -10'd42, -10'd36, -10'd57, 10'd22, -10'd53, 10'd31, -10'd21, -10'd17, 10'd3, -10'd24, 10'd51, -10'd43, -10'd44, 10'd37, 10'd60, 10'd16, 10'd76, -10'd14, 10'd55, -10'd28, 10'd13, -10'd68, -10'd51, -10'd34, -10'd48, 10'd25, 10'd27, -10'd36, 10'd5, 10'd38, 10'd42, 10'd66, -10'd16, 10'd33, 10'd33, -10'd25, 10'd13, -10'd67, 10'd52, -10'd1, -10'd36, -10'd9, -10'd19, -10'd5, 10'd21, -10'd36, 10'd50, -10'd44, 10'd31, 10'd36, -10'd34, -10'd44, 10'd18, 10'd69, 10'd35, -10'd23, 10'd45, -10'd43, -10'd9, -10'd21, -10'd31, 10'd45, 10'd40, -10'd18, 10'd21, 10'd34, 10'd35, 10'd46, 10'd32, 10'd25, -10'd48, 10'd16, 10'd29, 10'd26, 10'd37, -10'd22, -10'd48, -10'd16, -10'd38, 10'd28, -10'd44, 10'd38, 10'd6, 10'd41, -10'd28, -10'd35, -10'd1, -10'd13, 10'd32, 10'd23, 10'd27, 10'd41, 10'd68, -10'd53, 10'd29, -10'd28, 10'd59, 10'd11, 10'd48, -10'd7, 10'd29, 10'd71, -10'd37, -10'd28, 10'd29, -10'd63, -10'd9, -10'd30, -10'd31, -10'd58, -10'd42, 10'd45, 10'd46, -10'd36, 10'd25, -10'd24, 10'd46, 10'd39, 10'd11, 10'd34, -10'd28, 10'd19, -10'd23, 10'd31, -10'd48, 10'd55, 10'd5, 10'd62, 10'd32, -10'd39, -10'd36, 10'd7, -10'd43, -10'd47, 10'd28, 10'd43, -10'd16, 10'd28, -10'd33, -10'd51, 10'd43, -10'd50, 10'd17, -10'd14, -10'd35, -10'd23, -10'd49, -10'd36, -10'd27, 10'd5, 10'd66, -10'd22, -10'd26, -10'd21, -10'd23, 10'd29, 10'd9, -10'd55, -10'd24, -10'd16, -10'd66, 10'd28, 10'd29, -10'd35, -10'd27, 10'd43, -10'd67, 10'd40, -10'd42, -10'd31, 10'd33, -10'd47, -10'd23, -10'd35, -10'd31, 10'd32, 10'd38, -10'd40, 10'd15, 10'd26, 10'd31, -10'd33, -10'd22, -10'd26, 10'd31, -10'd17, -10'd28, 10'd21, -10'd44, 10'd20, 10'd23, -10'd61, -10'd30, -10'd23, 10'd46, -10'd47, -10'd44, -10'd1, -10'd51, 10'd73, 10'd39, 10'd22, -10'd39, 10'd13, 10'd53, -10'd12, -10'd59, 10'd1, -10'd75, -10'd20, -10'd55, 10'd37, -10'd28, 10'd24, 10'd73, 10'd32, -10'd25, -10'd60, -10'd24, 10'd27, 10'd36, 10'd53, -10'd38, 10'd30, -10'd45, -10'd44, -10'd18, -10'd35, -10'd66, -10'd48, -10'd55, 10'd69, -10'd31, -10'd19, 10'd7, -10'd28, 10'd47, 10'd33, 10'd23, 10'd35, 10'd38, -10'd23, 10'd6, 10'd4, 10'd46, -10'd31, 10'd40, 10'd25, -10'd65, 10'd31, -10'd30, -10'd35, -10'd30, -10'd32, -10'd27, -10'd60, 10'd3, -10'd36, -10'd46, -10'd27, 10'd47, -10'd65, -10'd16, 10'd35, -10'd2, -10'd85, 10'd35, -10'd54, -10'd25, -10'd52, 10'd21, -10'd28, -10'd30, -10'd4, 10'd62, 10'd12, -10'd22, 10'd24, 10'd59, 10'd19, -10'd2, -10'd47, 10'd33, 10'd14, 10'd67, -10'd19, -10'd49, -10'd61, 10'd40, 10'd64, 10'd28, 10'd66, -10'd14, -10'd16, -10'd56, -10'd23, -10'd6, -10'd56, -10'd13, -10'd32, 10'd42, 10'd46, -10'd25, -10'd37, -10'd1, 10'd26, 10'd33, -10'd56, 10'd13, 10'd12, 10'd45, 10'd24, 10'd46, -10'd24, -10'd65, -10'd43, 10'd37, 10'd15, 10'd33, -10'd67, 10'd53, -10'd27, -10'd66, -10'd14, -10'd53, -10'd56, -10'd26, -10'd33, 10'd9, -10'd26, 10'd46, 10'd16, -10'd63, 10'd32, -10'd28, -10'd21, 10'd33, -10'd36, -10'd6, -10'd31, 10'd58, 10'd34, -10'd40, 10'd36, -10'd53, -10'd48, 10'd59, 10'd2, 10'd46, -10'd49, -10'd18, 10'd35, 10'd71, -10'd13, -10'd74, -10'd32, 10'd40, 10'd26, -10'd15, 10'd19, -10'd6, -10'd59, -10'd37, -10'd13, 10'd63, 10'd48, 10'd21, -10'd51, 10'd53, 10'd43, -10'd37, -10'd29, 10'd58, 10'd20, 10'd27, 10'd29, -10'd21, -10'd0, 10'd66, 10'd57, -10'd60, -10'd35, 10'd10, -10'd20, -10'd7, 10'd63, 10'd53, -10'd21, 10'd36, 10'd9, -10'd14, 10'd60, -10'd36, -10'd3, 10'd5, -10'd24, -10'd66, 10'd16, -10'd22, -10'd49, 10'd57, 10'd61, -10'd34, -10'd48, 10'd3, 10'd20, -10'd7, 10'd23, -10'd22, -10'd43, 10'd2, -10'd56, -10'd46, 10'd28, 10'd40, -10'd26, 10'd14, -10'd25, -10'd46, 10'd36, 10'd69, -10'd36, -10'd34, -10'd45, -10'd73, 10'd55, 10'd6, -10'd33, 10'd12, 10'd43, 10'd52, 10'd41, 10'd43, -10'd15, 10'd43, -10'd26, 10'd35, -10'd47, -10'd42, -10'd70, -10'd19, 10'd50, -10'd38, 10'd24, 10'd67, -10'd32, 10'd41, -10'd39, 10'd19, -10'd29, -10'd35, 10'd55, 10'd12, 10'd11, -10'd24, -10'd59, -10'd56, -10'd41, 10'd34, 10'd14, 10'd68, 10'd16, -10'd9, 10'd37, 10'd5, 10'd51, 10'd35, -10'd12, 10'd25, -10'd20, -10'd46, 10'd35, 10'd20, 10'd36, 10'd32, -10'd2, 10'd44, -10'd29, 10'd54, 10'd33, -10'd38, 10'd40, 10'd65, -10'd48, -10'd6, -10'd64, -10'd21, -10'd20, 10'd39, -10'd42, -10'd19, 10'd23, -10'd34, -10'd7, -10'd33, 10'd41, 10'd82, 10'd42, 10'd37, 10'd38, 10'd50, 10'd42, 10'd27, 10'd17, 10'd23, -10'd65, -10'd43, 10'd43, 10'd62, 10'd18, -10'd28, 10'd34, -10'd11, -10'd31, 10'd13, 10'd38, -10'd7, 10'd54, -10'd34, 10'd45, 10'd26, 10'd33, -10'd69, 10'd23, -10'd52, 10'd29, -10'd47, -10'd61, 10'd79, -10'd30, -10'd43, -10'd8, 10'd30, 10'd33, 10'd32, -10'd44, 10'd50, -10'd17, 10'd25, -10'd57};
wire done;
wire [1439:0] Bit;
wire [1439:0] Check_Bit;
assign Check_Bit[0] = (Bit[0] == 1) ? 1 : 0;
assign Check_Bit[1] = (Bit[1] == 0) ? 1 : 0;
assign Check_Bit[2] = (Bit[2] == 1) ? 1 : 0;
assign Check_Bit[3] = (Bit[3] == 0) ? 1 : 0;
assign Check_Bit[4] = (Bit[4] == 1) ? 1 : 0;
assign Check_Bit[5] = (Bit[5] == 0) ? 1 : 0;
assign Check_Bit[6] = (Bit[6] == 0) ? 1 : 0;
assign Check_Bit[7] = (Bit[7] == 0) ? 1 : 0;
assign Check_Bit[8] = (Bit[8] == 0) ? 1 : 0;
assign Check_Bit[9] = (Bit[9] == 1) ? 1 : 0;
assign Check_Bit[10] = (Bit[10] == 1) ? 1 : 0;
assign Check_Bit[11] = (Bit[11] == 0) ? 1 : 0;
assign Check_Bit[12] = (Bit[12] == 1) ? 1 : 0;
assign Check_Bit[13] = (Bit[13] == 1) ? 1 : 0;
assign Check_Bit[14] = (Bit[14] == 0) ? 1 : 0;
assign Check_Bit[15] = (Bit[15] == 1) ? 1 : 0;
assign Check_Bit[16] = (Bit[16] == 0) ? 1 : 0;
assign Check_Bit[17] = (Bit[17] == 1) ? 1 : 0;
assign Check_Bit[18] = (Bit[18] == 0) ? 1 : 0;
assign Check_Bit[19] = (Bit[19] == 0) ? 1 : 0;
assign Check_Bit[20] = (Bit[20] == 0) ? 1 : 0;
assign Check_Bit[21] = (Bit[21] == 1) ? 1 : 0;
assign Check_Bit[22] = (Bit[22] == 0) ? 1 : 0;
assign Check_Bit[23] = (Bit[23] == 1) ? 1 : 0;
assign Check_Bit[24] = (Bit[24] == 0) ? 1 : 0;
assign Check_Bit[25] = (Bit[25] == 0) ? 1 : 0;
assign Check_Bit[26] = (Bit[26] == 1) ? 1 : 0;
assign Check_Bit[27] = (Bit[27] == 1) ? 1 : 0;
assign Check_Bit[28] = (Bit[28] == 0) ? 1 : 0;
assign Check_Bit[29] = (Bit[29] == 1) ? 1 : 0;
assign Check_Bit[30] = (Bit[30] == 0) ? 1 : 0;
assign Check_Bit[31] = (Bit[31] == 0) ? 1 : 0;
assign Check_Bit[32] = (Bit[32] == 0) ? 1 : 0;
assign Check_Bit[33] = (Bit[33] == 1) ? 1 : 0;
assign Check_Bit[34] = (Bit[34] == 1) ? 1 : 0;
assign Check_Bit[35] = (Bit[35] == 0) ? 1 : 0;
assign Check_Bit[36] = (Bit[36] == 0) ? 1 : 0;
assign Check_Bit[37] = (Bit[37] == 0) ? 1 : 0;
assign Check_Bit[38] = (Bit[38] == 0) ? 1 : 0;
assign Check_Bit[39] = (Bit[39] == 0) ? 1 : 0;
assign Check_Bit[40] = (Bit[40] == 0) ? 1 : 0;
assign Check_Bit[41] = (Bit[41] == 0) ? 1 : 0;
assign Check_Bit[42] = (Bit[42] == 0) ? 1 : 0;
assign Check_Bit[43] = (Bit[43] == 0) ? 1 : 0;
assign Check_Bit[44] = (Bit[44] == 0) ? 1 : 0;
assign Check_Bit[45] = (Bit[45] == 1) ? 1 : 0;
assign Check_Bit[46] = (Bit[46] == 1) ? 1 : 0;
assign Check_Bit[47] = (Bit[47] == 1) ? 1 : 0;
assign Check_Bit[48] = (Bit[48] == 0) ? 1 : 0;
assign Check_Bit[49] = (Bit[49] == 1) ? 1 : 0;
assign Check_Bit[50] = (Bit[50] == 1) ? 1 : 0;
assign Check_Bit[51] = (Bit[51] == 0) ? 1 : 0;
assign Check_Bit[52] = (Bit[52] == 1) ? 1 : 0;
assign Check_Bit[53] = (Bit[53] == 1) ? 1 : 0;
assign Check_Bit[54] = (Bit[54] == 1) ? 1 : 0;
assign Check_Bit[55] = (Bit[55] == 0) ? 1 : 0;
assign Check_Bit[56] = (Bit[56] == 1) ? 1 : 0;
assign Check_Bit[57] = (Bit[57] == 0) ? 1 : 0;
assign Check_Bit[58] = (Bit[58] == 0) ? 1 : 0;
assign Check_Bit[59] = (Bit[59] == 1) ? 1 : 0;
assign Check_Bit[60] = (Bit[60] == 0) ? 1 : 0;
assign Check_Bit[61] = (Bit[61] == 0) ? 1 : 0;
assign Check_Bit[62] = (Bit[62] == 1) ? 1 : 0;
assign Check_Bit[63] = (Bit[63] == 0) ? 1 : 0;
assign Check_Bit[64] = (Bit[64] == 0) ? 1 : 0;
assign Check_Bit[65] = (Bit[65] == 0) ? 1 : 0;
assign Check_Bit[66] = (Bit[66] == 0) ? 1 : 0;
assign Check_Bit[67] = (Bit[67] == 0) ? 1 : 0;
assign Check_Bit[68] = (Bit[68] == 0) ? 1 : 0;
assign Check_Bit[69] = (Bit[69] == 1) ? 1 : 0;
assign Check_Bit[70] = (Bit[70] == 1) ? 1 : 0;
assign Check_Bit[71] = (Bit[71] == 0) ? 1 : 0;
assign Check_Bit[72] = (Bit[72] == 1) ? 1 : 0;
assign Check_Bit[73] = (Bit[73] == 0) ? 1 : 0;
assign Check_Bit[74] = (Bit[74] == 0) ? 1 : 0;
assign Check_Bit[75] = (Bit[75] == 1) ? 1 : 0;
assign Check_Bit[76] = (Bit[76] == 0) ? 1 : 0;
assign Check_Bit[77] = (Bit[77] == 1) ? 1 : 0;
assign Check_Bit[78] = (Bit[78] == 0) ? 1 : 0;
assign Check_Bit[79] = (Bit[79] == 0) ? 1 : 0;
assign Check_Bit[80] = (Bit[80] == 0) ? 1 : 0;
assign Check_Bit[81] = (Bit[81] == 0) ? 1 : 0;
assign Check_Bit[82] = (Bit[82] == 1) ? 1 : 0;
assign Check_Bit[83] = (Bit[83] == 1) ? 1 : 0;
assign Check_Bit[84] = (Bit[84] == 1) ? 1 : 0;
assign Check_Bit[85] = (Bit[85] == 1) ? 1 : 0;
assign Check_Bit[86] = (Bit[86] == 0) ? 1 : 0;
assign Check_Bit[87] = (Bit[87] == 0) ? 1 : 0;
assign Check_Bit[88] = (Bit[88] == 0) ? 1 : 0;
assign Check_Bit[89] = (Bit[89] == 1) ? 1 : 0;
assign Check_Bit[90] = (Bit[90] == 1) ? 1 : 0;
assign Check_Bit[91] = (Bit[91] == 0) ? 1 : 0;
assign Check_Bit[92] = (Bit[92] == 1) ? 1 : 0;
assign Check_Bit[93] = (Bit[93] == 0) ? 1 : 0;
assign Check_Bit[94] = (Bit[94] == 1) ? 1 : 0;
assign Check_Bit[95] = (Bit[95] == 0) ? 1 : 0;
assign Check_Bit[96] = (Bit[96] == 0) ? 1 : 0;
assign Check_Bit[97] = (Bit[97] == 1) ? 1 : 0;
assign Check_Bit[98] = (Bit[98] == 0) ? 1 : 0;
assign Check_Bit[99] = (Bit[99] == 1) ? 1 : 0;
assign Check_Bit[100] = (Bit[100] == 1) ? 1 : 0;
assign Check_Bit[101] = (Bit[101] == 1) ? 1 : 0;
assign Check_Bit[102] = (Bit[102] == 1) ? 1 : 0;
assign Check_Bit[103] = (Bit[103] == 0) ? 1 : 0;
assign Check_Bit[104] = (Bit[104] == 1) ? 1 : 0;
assign Check_Bit[105] = (Bit[105] == 0) ? 1 : 0;
assign Check_Bit[106] = (Bit[106] == 1) ? 1 : 0;
assign Check_Bit[107] = (Bit[107] == 0) ? 1 : 0;
assign Check_Bit[108] = (Bit[108] == 0) ? 1 : 0;
assign Check_Bit[109] = (Bit[109] == 0) ? 1 : 0;
assign Check_Bit[110] = (Bit[110] == 0) ? 1 : 0;
assign Check_Bit[111] = (Bit[111] == 0) ? 1 : 0;
assign Check_Bit[112] = (Bit[112] == 1) ? 1 : 0;
assign Check_Bit[113] = (Bit[113] == 0) ? 1 : 0;
assign Check_Bit[114] = (Bit[114] == 0) ? 1 : 0;
assign Check_Bit[115] = (Bit[115] == 1) ? 1 : 0;
assign Check_Bit[116] = (Bit[116] == 1) ? 1 : 0;
assign Check_Bit[117] = (Bit[117] == 1) ? 1 : 0;
assign Check_Bit[118] = (Bit[118] == 1) ? 1 : 0;
assign Check_Bit[119] = (Bit[119] == 0) ? 1 : 0;
assign Check_Bit[120] = (Bit[120] == 0) ? 1 : 0;
assign Check_Bit[121] = (Bit[121] == 1) ? 1 : 0;
assign Check_Bit[122] = (Bit[122] == 1) ? 1 : 0;
assign Check_Bit[123] = (Bit[123] == 0) ? 1 : 0;
assign Check_Bit[124] = (Bit[124] == 1) ? 1 : 0;
assign Check_Bit[125] = (Bit[125] == 0) ? 1 : 0;
assign Check_Bit[126] = (Bit[126] == 0) ? 1 : 0;
assign Check_Bit[127] = (Bit[127] == 1) ? 1 : 0;
assign Check_Bit[128] = (Bit[128] == 1) ? 1 : 0;
assign Check_Bit[129] = (Bit[129] == 0) ? 1 : 0;
assign Check_Bit[130] = (Bit[130] == 1) ? 1 : 0;
assign Check_Bit[131] = (Bit[131] == 1) ? 1 : 0;
assign Check_Bit[132] = (Bit[132] == 0) ? 1 : 0;
assign Check_Bit[133] = (Bit[133] == 1) ? 1 : 0;
assign Check_Bit[134] = (Bit[134] == 0) ? 1 : 0;
assign Check_Bit[135] = (Bit[135] == 1) ? 1 : 0;
assign Check_Bit[136] = (Bit[136] == 1) ? 1 : 0;
assign Check_Bit[137] = (Bit[137] == 1) ? 1 : 0;
assign Check_Bit[138] = (Bit[138] == 0) ? 1 : 0;
assign Check_Bit[139] = (Bit[139] == 0) ? 1 : 0;
assign Check_Bit[140] = (Bit[140] == 1) ? 1 : 0;
assign Check_Bit[141] = (Bit[141] == 1) ? 1 : 0;
assign Check_Bit[142] = (Bit[142] == 0) ? 1 : 0;
assign Check_Bit[143] = (Bit[143] == 1) ? 1 : 0;
assign Check_Bit[144] = (Bit[144] == 1) ? 1 : 0;
assign Check_Bit[145] = (Bit[145] == 0) ? 1 : 0;
assign Check_Bit[146] = (Bit[146] == 0) ? 1 : 0;
assign Check_Bit[147] = (Bit[147] == 1) ? 1 : 0;
assign Check_Bit[148] = (Bit[148] == 0) ? 1 : 0;
assign Check_Bit[149] = (Bit[149] == 1) ? 1 : 0;
assign Check_Bit[150] = (Bit[150] == 0) ? 1 : 0;
assign Check_Bit[151] = (Bit[151] == 0) ? 1 : 0;
assign Check_Bit[152] = (Bit[152] == 1) ? 1 : 0;
assign Check_Bit[153] = (Bit[153] == 0) ? 1 : 0;
assign Check_Bit[154] = (Bit[154] == 0) ? 1 : 0;
assign Check_Bit[155] = (Bit[155] == 1) ? 1 : 0;
assign Check_Bit[156] = (Bit[156] == 1) ? 1 : 0;
assign Check_Bit[157] = (Bit[157] == 0) ? 1 : 0;
assign Check_Bit[158] = (Bit[158] == 1) ? 1 : 0;
assign Check_Bit[159] = (Bit[159] == 1) ? 1 : 0;
assign Check_Bit[160] = (Bit[160] == 0) ? 1 : 0;
assign Check_Bit[161] = (Bit[161] == 0) ? 1 : 0;
assign Check_Bit[162] = (Bit[162] == 0) ? 1 : 0;
assign Check_Bit[163] = (Bit[163] == 1) ? 1 : 0;
assign Check_Bit[164] = (Bit[164] == 0) ? 1 : 0;
assign Check_Bit[165] = (Bit[165] == 0) ? 1 : 0;
assign Check_Bit[166] = (Bit[166] == 0) ? 1 : 0;
assign Check_Bit[167] = (Bit[167] == 0) ? 1 : 0;
assign Check_Bit[168] = (Bit[168] == 1) ? 1 : 0;
assign Check_Bit[169] = (Bit[169] == 1) ? 1 : 0;
assign Check_Bit[170] = (Bit[170] == 0) ? 1 : 0;
assign Check_Bit[171] = (Bit[171] == 0) ? 1 : 0;
assign Check_Bit[172] = (Bit[172] == 1) ? 1 : 0;
assign Check_Bit[173] = (Bit[173] == 0) ? 1 : 0;
assign Check_Bit[174] = (Bit[174] == 0) ? 1 : 0;
assign Check_Bit[175] = (Bit[175] == 0) ? 1 : 0;
assign Check_Bit[176] = (Bit[176] == 1) ? 1 : 0;
assign Check_Bit[177] = (Bit[177] == 1) ? 1 : 0;
assign Check_Bit[178] = (Bit[178] == 1) ? 1 : 0;
assign Check_Bit[179] = (Bit[179] == 0) ? 1 : 0;
assign Check_Bit[180] = (Bit[180] == 0) ? 1 : 0;
assign Check_Bit[181] = (Bit[181] == 1) ? 1 : 0;
assign Check_Bit[182] = (Bit[182] == 0) ? 1 : 0;
assign Check_Bit[183] = (Bit[183] == 0) ? 1 : 0;
assign Check_Bit[184] = (Bit[184] == 1) ? 1 : 0;
assign Check_Bit[185] = (Bit[185] == 1) ? 1 : 0;
assign Check_Bit[186] = (Bit[186] == 1) ? 1 : 0;
assign Check_Bit[187] = (Bit[187] == 0) ? 1 : 0;
assign Check_Bit[188] = (Bit[188] == 0) ? 1 : 0;
assign Check_Bit[189] = (Bit[189] == 1) ? 1 : 0;
assign Check_Bit[190] = (Bit[190] == 1) ? 1 : 0;
assign Check_Bit[191] = (Bit[191] == 0) ? 1 : 0;
assign Check_Bit[192] = (Bit[192] == 1) ? 1 : 0;
assign Check_Bit[193] = (Bit[193] == 0) ? 1 : 0;
assign Check_Bit[194] = (Bit[194] == 1) ? 1 : 0;
assign Check_Bit[195] = (Bit[195] == 1) ? 1 : 0;
assign Check_Bit[196] = (Bit[196] == 0) ? 1 : 0;
assign Check_Bit[197] = (Bit[197] == 1) ? 1 : 0;
assign Check_Bit[198] = (Bit[198] == 0) ? 1 : 0;
assign Check_Bit[199] = (Bit[199] == 0) ? 1 : 0;
assign Check_Bit[200] = (Bit[200] == 1) ? 1 : 0;
assign Check_Bit[201] = (Bit[201] == 1) ? 1 : 0;
assign Check_Bit[202] = (Bit[202] == 1) ? 1 : 0;
assign Check_Bit[203] = (Bit[203] == 0) ? 1 : 0;
assign Check_Bit[204] = (Bit[204] == 1) ? 1 : 0;
assign Check_Bit[205] = (Bit[205] == 1) ? 1 : 0;
assign Check_Bit[206] = (Bit[206] == 0) ? 1 : 0;
assign Check_Bit[207] = (Bit[207] == 1) ? 1 : 0;
assign Check_Bit[208] = (Bit[208] == 0) ? 1 : 0;
assign Check_Bit[209] = (Bit[209] == 0) ? 1 : 0;
assign Check_Bit[210] = (Bit[210] == 1) ? 1 : 0;
assign Check_Bit[211] = (Bit[211] == 0) ? 1 : 0;
assign Check_Bit[212] = (Bit[212] == 1) ? 1 : 0;
assign Check_Bit[213] = (Bit[213] == 1) ? 1 : 0;
assign Check_Bit[214] = (Bit[214] == 1) ? 1 : 0;
assign Check_Bit[215] = (Bit[215] == 1) ? 1 : 0;
assign Check_Bit[216] = (Bit[216] == 1) ? 1 : 0;
assign Check_Bit[217] = (Bit[217] == 1) ? 1 : 0;
assign Check_Bit[218] = (Bit[218] == 1) ? 1 : 0;
assign Check_Bit[219] = (Bit[219] == 0) ? 1 : 0;
assign Check_Bit[220] = (Bit[220] == 1) ? 1 : 0;
assign Check_Bit[221] = (Bit[221] == 0) ? 1 : 0;
assign Check_Bit[222] = (Bit[222] == 0) ? 1 : 0;
assign Check_Bit[223] = (Bit[223] == 0) ? 1 : 0;
assign Check_Bit[224] = (Bit[224] == 1) ? 1 : 0;
assign Check_Bit[225] = (Bit[225] == 1) ? 1 : 0;
assign Check_Bit[226] = (Bit[226] == 1) ? 1 : 0;
assign Check_Bit[227] = (Bit[227] == 0) ? 1 : 0;
assign Check_Bit[228] = (Bit[228] == 0) ? 1 : 0;
assign Check_Bit[229] = (Bit[229] == 0) ? 1 : 0;
assign Check_Bit[230] = (Bit[230] == 0) ? 1 : 0;
assign Check_Bit[231] = (Bit[231] == 0) ? 1 : 0;
assign Check_Bit[232] = (Bit[232] == 1) ? 1 : 0;
assign Check_Bit[233] = (Bit[233] == 0) ? 1 : 0;
assign Check_Bit[234] = (Bit[234] == 0) ? 1 : 0;
assign Check_Bit[235] = (Bit[235] == 1) ? 1 : 0;
assign Check_Bit[236] = (Bit[236] == 1) ? 1 : 0;
assign Check_Bit[237] = (Bit[237] == 1) ? 1 : 0;
assign Check_Bit[238] = (Bit[238] == 0) ? 1 : 0;
assign Check_Bit[239] = (Bit[239] == 0) ? 1 : 0;
assign Check_Bit[240] = (Bit[240] == 1) ? 1 : 0;
assign Check_Bit[241] = (Bit[241] == 1) ? 1 : 0;
assign Check_Bit[242] = (Bit[242] == 1) ? 1 : 0;
assign Check_Bit[243] = (Bit[243] == 1) ? 1 : 0;
assign Check_Bit[244] = (Bit[244] == 1) ? 1 : 0;
assign Check_Bit[245] = (Bit[245] == 1) ? 1 : 0;
assign Check_Bit[246] = (Bit[246] == 1) ? 1 : 0;
assign Check_Bit[247] = (Bit[247] == 1) ? 1 : 0;
assign Check_Bit[248] = (Bit[248] == 0) ? 1 : 0;
assign Check_Bit[249] = (Bit[249] == 0) ? 1 : 0;
assign Check_Bit[250] = (Bit[250] == 0) ? 1 : 0;
assign Check_Bit[251] = (Bit[251] == 0) ? 1 : 0;
assign Check_Bit[252] = (Bit[252] == 1) ? 1 : 0;
assign Check_Bit[253] = (Bit[253] == 1) ? 1 : 0;
assign Check_Bit[254] = (Bit[254] == 1) ? 1 : 0;
assign Check_Bit[255] = (Bit[255] == 0) ? 1 : 0;
assign Check_Bit[256] = (Bit[256] == 0) ? 1 : 0;
assign Check_Bit[257] = (Bit[257] == 0) ? 1 : 0;
assign Check_Bit[258] = (Bit[258] == 1) ? 1 : 0;
assign Check_Bit[259] = (Bit[259] == 1) ? 1 : 0;
assign Check_Bit[260] = (Bit[260] == 0) ? 1 : 0;
assign Check_Bit[261] = (Bit[261] == 0) ? 1 : 0;
assign Check_Bit[262] = (Bit[262] == 0) ? 1 : 0;
assign Check_Bit[263] = (Bit[263] == 1) ? 1 : 0;
assign Check_Bit[264] = (Bit[264] == 0) ? 1 : 0;
assign Check_Bit[265] = (Bit[265] == 0) ? 1 : 0;
assign Check_Bit[266] = (Bit[266] == 0) ? 1 : 0;
assign Check_Bit[267] = (Bit[267] == 1) ? 1 : 0;
assign Check_Bit[268] = (Bit[268] == 1) ? 1 : 0;
assign Check_Bit[269] = (Bit[269] == 0) ? 1 : 0;
assign Check_Bit[270] = (Bit[270] == 1) ? 1 : 0;
assign Check_Bit[271] = (Bit[271] == 1) ? 1 : 0;
assign Check_Bit[272] = (Bit[272] == 1) ? 1 : 0;
assign Check_Bit[273] = (Bit[273] == 0) ? 1 : 0;
assign Check_Bit[274] = (Bit[274] == 1) ? 1 : 0;
assign Check_Bit[275] = (Bit[275] == 0) ? 1 : 0;
assign Check_Bit[276] = (Bit[276] == 0) ? 1 : 0;
assign Check_Bit[277] = (Bit[277] == 1) ? 1 : 0;
assign Check_Bit[278] = (Bit[278] == 1) ? 1 : 0;
assign Check_Bit[279] = (Bit[279] == 0) ? 1 : 0;
assign Check_Bit[280] = (Bit[280] == 1) ? 1 : 0;
assign Check_Bit[281] = (Bit[281] == 1) ? 1 : 0;
assign Check_Bit[282] = (Bit[282] == 1) ? 1 : 0;
assign Check_Bit[283] = (Bit[283] == 1) ? 1 : 0;
assign Check_Bit[284] = (Bit[284] == 1) ? 1 : 0;
assign Check_Bit[285] = (Bit[285] == 1) ? 1 : 0;
assign Check_Bit[286] = (Bit[286] == 1) ? 1 : 0;
assign Check_Bit[287] = (Bit[287] == 1) ? 1 : 0;
assign Check_Bit[288] = (Bit[288] == 1) ? 1 : 0;
assign Check_Bit[289] = (Bit[289] == 1) ? 1 : 0;
assign Check_Bit[290] = (Bit[290] == 0) ? 1 : 0;
assign Check_Bit[291] = (Bit[291] == 1) ? 1 : 0;
assign Check_Bit[292] = (Bit[292] == 0) ? 1 : 0;
assign Check_Bit[293] = (Bit[293] == 0) ? 1 : 0;
assign Check_Bit[294] = (Bit[294] == 1) ? 1 : 0;
assign Check_Bit[295] = (Bit[295] == 0) ? 1 : 0;
assign Check_Bit[296] = (Bit[296] == 1) ? 1 : 0;
assign Check_Bit[297] = (Bit[297] == 0) ? 1 : 0;
assign Check_Bit[298] = (Bit[298] == 1) ? 1 : 0;
assign Check_Bit[299] = (Bit[299] == 0) ? 1 : 0;
assign Check_Bit[300] = (Bit[300] == 0) ? 1 : 0;
assign Check_Bit[301] = (Bit[301] == 0) ? 1 : 0;
assign Check_Bit[302] = (Bit[302] == 0) ? 1 : 0;
assign Check_Bit[303] = (Bit[303] == 0) ? 1 : 0;
assign Check_Bit[304] = (Bit[304] == 1) ? 1 : 0;
assign Check_Bit[305] = (Bit[305] == 0) ? 1 : 0;
assign Check_Bit[306] = (Bit[306] == 1) ? 1 : 0;
assign Check_Bit[307] = (Bit[307] == 1) ? 1 : 0;
assign Check_Bit[308] = (Bit[308] == 0) ? 1 : 0;
assign Check_Bit[309] = (Bit[309] == 1) ? 1 : 0;
assign Check_Bit[310] = (Bit[310] == 1) ? 1 : 0;
assign Check_Bit[311] = (Bit[311] == 1) ? 1 : 0;
assign Check_Bit[312] = (Bit[312] == 1) ? 1 : 0;
assign Check_Bit[313] = (Bit[313] == 1) ? 1 : 0;
assign Check_Bit[314] = (Bit[314] == 1) ? 1 : 0;
assign Check_Bit[315] = (Bit[315] == 1) ? 1 : 0;
assign Check_Bit[316] = (Bit[316] == 0) ? 1 : 0;
assign Check_Bit[317] = (Bit[317] == 1) ? 1 : 0;
assign Check_Bit[318] = (Bit[318] == 0) ? 1 : 0;
assign Check_Bit[319] = (Bit[319] == 0) ? 1 : 0;
assign Check_Bit[320] = (Bit[320] == 0) ? 1 : 0;
assign Check_Bit[321] = (Bit[321] == 1) ? 1 : 0;
assign Check_Bit[322] = (Bit[322] == 1) ? 1 : 0;
assign Check_Bit[323] = (Bit[323] == 1) ? 1 : 0;
assign Check_Bit[324] = (Bit[324] == 0) ? 1 : 0;
assign Check_Bit[325] = (Bit[325] == 0) ? 1 : 0;
assign Check_Bit[326] = (Bit[326] == 0) ? 1 : 0;
assign Check_Bit[327] = (Bit[327] == 1) ? 1 : 0;
assign Check_Bit[328] = (Bit[328] == 0) ? 1 : 0;
assign Check_Bit[329] = (Bit[329] == 1) ? 1 : 0;
assign Check_Bit[330] = (Bit[330] == 1) ? 1 : 0;
assign Check_Bit[331] = (Bit[331] == 1) ? 1 : 0;
assign Check_Bit[332] = (Bit[332] == 0) ? 1 : 0;
assign Check_Bit[333] = (Bit[333] == 1) ? 1 : 0;
assign Check_Bit[334] = (Bit[334] == 1) ? 1 : 0;
assign Check_Bit[335] = (Bit[335] == 0) ? 1 : 0;
assign Check_Bit[336] = (Bit[336] == 0) ? 1 : 0;
assign Check_Bit[337] = (Bit[337] == 1) ? 1 : 0;
assign Check_Bit[338] = (Bit[338] == 0) ? 1 : 0;
assign Check_Bit[339] = (Bit[339] == 0) ? 1 : 0;
assign Check_Bit[340] = (Bit[340] == 0) ? 1 : 0;
assign Check_Bit[341] = (Bit[341] == 1) ? 1 : 0;
assign Check_Bit[342] = (Bit[342] == 1) ? 1 : 0;
assign Check_Bit[343] = (Bit[343] == 1) ? 1 : 0;
assign Check_Bit[344] = (Bit[344] == 1) ? 1 : 0;
assign Check_Bit[345] = (Bit[345] == 0) ? 1 : 0;
assign Check_Bit[346] = (Bit[346] == 1) ? 1 : 0;
assign Check_Bit[347] = (Bit[347] == 1) ? 1 : 0;
assign Check_Bit[348] = (Bit[348] == 1) ? 1 : 0;
assign Check_Bit[349] = (Bit[349] == 0) ? 1 : 0;
assign Check_Bit[350] = (Bit[350] == 0) ? 1 : 0;
assign Check_Bit[351] = (Bit[351] == 1) ? 1 : 0;
assign Check_Bit[352] = (Bit[352] == 0) ? 1 : 0;
assign Check_Bit[353] = (Bit[353] == 1) ? 1 : 0;
assign Check_Bit[354] = (Bit[354] == 1) ? 1 : 0;
assign Check_Bit[355] = (Bit[355] == 0) ? 1 : 0;
assign Check_Bit[356] = (Bit[356] == 1) ? 1 : 0;
assign Check_Bit[357] = (Bit[357] == 1) ? 1 : 0;
assign Check_Bit[358] = (Bit[358] == 1) ? 1 : 0;
assign Check_Bit[359] = (Bit[359] == 0) ? 1 : 0;
assign Check_Bit[360] = (Bit[360] == 0) ? 1 : 0;
assign Check_Bit[361] = (Bit[361] == 0) ? 1 : 0;
assign Check_Bit[362] = (Bit[362] == 1) ? 1 : 0;
assign Check_Bit[363] = (Bit[363] == 0) ? 1 : 0;
assign Check_Bit[364] = (Bit[364] == 0) ? 1 : 0;
assign Check_Bit[365] = (Bit[365] == 1) ? 1 : 0;
assign Check_Bit[366] = (Bit[366] == 1) ? 1 : 0;
assign Check_Bit[367] = (Bit[367] == 1) ? 1 : 0;
assign Check_Bit[368] = (Bit[368] == 1) ? 1 : 0;
assign Check_Bit[369] = (Bit[369] == 0) ? 1 : 0;
assign Check_Bit[370] = (Bit[370] == 1) ? 1 : 0;
assign Check_Bit[371] = (Bit[371] == 1) ? 1 : 0;
assign Check_Bit[372] = (Bit[372] == 0) ? 1 : 0;
assign Check_Bit[373] = (Bit[373] == 1) ? 1 : 0;
assign Check_Bit[374] = (Bit[374] == 0) ? 1 : 0;
assign Check_Bit[375] = (Bit[375] == 1) ? 1 : 0;
assign Check_Bit[376] = (Bit[376] == 1) ? 1 : 0;
assign Check_Bit[377] = (Bit[377] == 0) ? 1 : 0;
assign Check_Bit[378] = (Bit[378] == 0) ? 1 : 0;
assign Check_Bit[379] = (Bit[379] == 1) ? 1 : 0;
assign Check_Bit[380] = (Bit[380] == 1) ? 1 : 0;
assign Check_Bit[381] = (Bit[381] == 1) ? 1 : 0;
assign Check_Bit[382] = (Bit[382] == 1) ? 1 : 0;
assign Check_Bit[383] = (Bit[383] == 0) ? 1 : 0;
assign Check_Bit[384] = (Bit[384] == 0) ? 1 : 0;
assign Check_Bit[385] = (Bit[385] == 1) ? 1 : 0;
assign Check_Bit[386] = (Bit[386] == 1) ? 1 : 0;
assign Check_Bit[387] = (Bit[387] == 1) ? 1 : 0;
assign Check_Bit[388] = (Bit[388] == 1) ? 1 : 0;
assign Check_Bit[389] = (Bit[389] == 0) ? 1 : 0;
assign Check_Bit[390] = (Bit[390] == 0) ? 1 : 0;
assign Check_Bit[391] = (Bit[391] == 1) ? 1 : 0;
assign Check_Bit[392] = (Bit[392] == 1) ? 1 : 0;
assign Check_Bit[393] = (Bit[393] == 1) ? 1 : 0;
assign Check_Bit[394] = (Bit[394] == 1) ? 1 : 0;
assign Check_Bit[395] = (Bit[395] == 1) ? 1 : 0;
assign Check_Bit[396] = (Bit[396] == 1) ? 1 : 0;
assign Check_Bit[397] = (Bit[397] == 0) ? 1 : 0;
assign Check_Bit[398] = (Bit[398] == 1) ? 1 : 0;
assign Check_Bit[399] = (Bit[399] == 0) ? 1 : 0;
assign Check_Bit[400] = (Bit[400] == 1) ? 1 : 0;
assign Check_Bit[401] = (Bit[401] == 1) ? 1 : 0;
assign Check_Bit[402] = (Bit[402] == 0) ? 1 : 0;
assign Check_Bit[403] = (Bit[403] == 1) ? 1 : 0;
assign Check_Bit[404] = (Bit[404] == 0) ? 1 : 0;
assign Check_Bit[405] = (Bit[405] == 0) ? 1 : 0;
assign Check_Bit[406] = (Bit[406] == 1) ? 1 : 0;
assign Check_Bit[407] = (Bit[407] == 1) ? 1 : 0;
assign Check_Bit[408] = (Bit[408] == 1) ? 1 : 0;
assign Check_Bit[409] = (Bit[409] == 1) ? 1 : 0;
assign Check_Bit[410] = (Bit[410] == 1) ? 1 : 0;
assign Check_Bit[411] = (Bit[411] == 0) ? 1 : 0;
assign Check_Bit[412] = (Bit[412] == 0) ? 1 : 0;
assign Check_Bit[413] = (Bit[413] == 0) ? 1 : 0;
assign Check_Bit[414] = (Bit[414] == 0) ? 1 : 0;
assign Check_Bit[415] = (Bit[415] == 1) ? 1 : 0;
assign Check_Bit[416] = (Bit[416] == 0) ? 1 : 0;
assign Check_Bit[417] = (Bit[417] == 1) ? 1 : 0;
assign Check_Bit[418] = (Bit[418] == 0) ? 1 : 0;
assign Check_Bit[419] = (Bit[419] == 1) ? 1 : 0;
assign Check_Bit[420] = (Bit[420] == 0) ? 1 : 0;
assign Check_Bit[421] = (Bit[421] == 0) ? 1 : 0;
assign Check_Bit[422] = (Bit[422] == 0) ? 1 : 0;
assign Check_Bit[423] = (Bit[423] == 0) ? 1 : 0;
assign Check_Bit[424] = (Bit[424] == 1) ? 1 : 0;
assign Check_Bit[425] = (Bit[425] == 0) ? 1 : 0;
assign Check_Bit[426] = (Bit[426] == 1) ? 1 : 0;
assign Check_Bit[427] = (Bit[427] == 0) ? 1 : 0;
assign Check_Bit[428] = (Bit[428] == 0) ? 1 : 0;
assign Check_Bit[429] = (Bit[429] == 1) ? 1 : 0;
assign Check_Bit[430] = (Bit[430] == 1) ? 1 : 0;
assign Check_Bit[431] = (Bit[431] == 1) ? 1 : 0;
assign Check_Bit[432] = (Bit[432] == 1) ? 1 : 0;
assign Check_Bit[433] = (Bit[433] == 1) ? 1 : 0;
assign Check_Bit[434] = (Bit[434] == 1) ? 1 : 0;
assign Check_Bit[435] = (Bit[435] == 0) ? 1 : 0;
assign Check_Bit[436] = (Bit[436] == 1) ? 1 : 0;
assign Check_Bit[437] = (Bit[437] == 1) ? 1 : 0;
assign Check_Bit[438] = (Bit[438] == 0) ? 1 : 0;
assign Check_Bit[439] = (Bit[439] == 0) ? 1 : 0;
assign Check_Bit[440] = (Bit[440] == 0) ? 1 : 0;
assign Check_Bit[441] = (Bit[441] == 0) ? 1 : 0;
assign Check_Bit[442] = (Bit[442] == 0) ? 1 : 0;
assign Check_Bit[443] = (Bit[443] == 0) ? 1 : 0;
assign Check_Bit[444] = (Bit[444] == 1) ? 1 : 0;
assign Check_Bit[445] = (Bit[445] == 0) ? 1 : 0;
assign Check_Bit[446] = (Bit[446] == 1) ? 1 : 0;
assign Check_Bit[447] = (Bit[447] == 0) ? 1 : 0;
assign Check_Bit[448] = (Bit[448] == 0) ? 1 : 0;
assign Check_Bit[449] = (Bit[449] == 0) ? 1 : 0;
assign Check_Bit[450] = (Bit[450] == 0) ? 1 : 0;
assign Check_Bit[451] = (Bit[451] == 0) ? 1 : 0;
assign Check_Bit[452] = (Bit[452] == 1) ? 1 : 0;
assign Check_Bit[453] = (Bit[453] == 1) ? 1 : 0;
assign Check_Bit[454] = (Bit[454] == 1) ? 1 : 0;
assign Check_Bit[455] = (Bit[455] == 1) ? 1 : 0;
assign Check_Bit[456] = (Bit[456] == 0) ? 1 : 0;
assign Check_Bit[457] = (Bit[457] == 0) ? 1 : 0;
assign Check_Bit[458] = (Bit[458] == 0) ? 1 : 0;
assign Check_Bit[459] = (Bit[459] == 1) ? 1 : 0;
assign Check_Bit[460] = (Bit[460] == 0) ? 1 : 0;
assign Check_Bit[461] = (Bit[461] == 1) ? 1 : 0;
assign Check_Bit[462] = (Bit[462] == 0) ? 1 : 0;
assign Check_Bit[463] = (Bit[463] == 1) ? 1 : 0;
assign Check_Bit[464] = (Bit[464] == 1) ? 1 : 0;
assign Check_Bit[465] = (Bit[465] == 0) ? 1 : 0;
assign Check_Bit[466] = (Bit[466] == 0) ? 1 : 0;
assign Check_Bit[467] = (Bit[467] == 0) ? 1 : 0;
assign Check_Bit[468] = (Bit[468] == 0) ? 1 : 0;
assign Check_Bit[469] = (Bit[469] == 1) ? 1 : 0;
assign Check_Bit[470] = (Bit[470] == 0) ? 1 : 0;
assign Check_Bit[471] = (Bit[471] == 0) ? 1 : 0;
assign Check_Bit[472] = (Bit[472] == 0) ? 1 : 0;
assign Check_Bit[473] = (Bit[473] == 0) ? 1 : 0;
assign Check_Bit[474] = (Bit[474] == 0) ? 1 : 0;
assign Check_Bit[475] = (Bit[475] == 0) ? 1 : 0;
assign Check_Bit[476] = (Bit[476] == 1) ? 1 : 0;
assign Check_Bit[477] = (Bit[477] == 0) ? 1 : 0;
assign Check_Bit[478] = (Bit[478] == 0) ? 1 : 0;
assign Check_Bit[479] = (Bit[479] == 1) ? 1 : 0;
assign Check_Bit[480] = (Bit[480] == 1) ? 1 : 0;
assign Check_Bit[481] = (Bit[481] == 1) ? 1 : 0;
assign Check_Bit[482] = (Bit[482] == 1) ? 1 : 0;
assign Check_Bit[483] = (Bit[483] == 0) ? 1 : 0;
assign Check_Bit[484] = (Bit[484] == 1) ? 1 : 0;
assign Check_Bit[485] = (Bit[485] == 0) ? 1 : 0;
assign Check_Bit[486] = (Bit[486] == 0) ? 1 : 0;
assign Check_Bit[487] = (Bit[487] == 0) ? 1 : 0;
assign Check_Bit[488] = (Bit[488] == 1) ? 1 : 0;
assign Check_Bit[489] = (Bit[489] == 1) ? 1 : 0;
assign Check_Bit[490] = (Bit[490] == 0) ? 1 : 0;
assign Check_Bit[491] = (Bit[491] == 0) ? 1 : 0;
assign Check_Bit[492] = (Bit[492] == 1) ? 1 : 0;
assign Check_Bit[493] = (Bit[493] == 0) ? 1 : 0;
assign Check_Bit[494] = (Bit[494] == 1) ? 1 : 0;
assign Check_Bit[495] = (Bit[495] == 0) ? 1 : 0;
assign Check_Bit[496] = (Bit[496] == 1) ? 1 : 0;
assign Check_Bit[497] = (Bit[497] == 1) ? 1 : 0;
assign Check_Bit[498] = (Bit[498] == 1) ? 1 : 0;
assign Check_Bit[499] = (Bit[499] == 1) ? 1 : 0;
assign Check_Bit[500] = (Bit[500] == 1) ? 1 : 0;
assign Check_Bit[501] = (Bit[501] == 0) ? 1 : 0;
assign Check_Bit[502] = (Bit[502] == 1) ? 1 : 0;
assign Check_Bit[503] = (Bit[503] == 0) ? 1 : 0;
assign Check_Bit[504] = (Bit[504] == 1) ? 1 : 0;
assign Check_Bit[505] = (Bit[505] == 0) ? 1 : 0;
assign Check_Bit[506] = (Bit[506] == 0) ? 1 : 0;
assign Check_Bit[507] = (Bit[507] == 1) ? 1 : 0;
assign Check_Bit[508] = (Bit[508] == 0) ? 1 : 0;
assign Check_Bit[509] = (Bit[509] == 0) ? 1 : 0;
assign Check_Bit[510] = (Bit[510] == 0) ? 1 : 0;
assign Check_Bit[511] = (Bit[511] == 1) ? 1 : 0;
assign Check_Bit[512] = (Bit[512] == 1) ? 1 : 0;
assign Check_Bit[513] = (Bit[513] == 0) ? 1 : 0;
assign Check_Bit[514] = (Bit[514] == 0) ? 1 : 0;
assign Check_Bit[515] = (Bit[515] == 1) ? 1 : 0;
assign Check_Bit[516] = (Bit[516] == 1) ? 1 : 0;
assign Check_Bit[517] = (Bit[517] == 1) ? 1 : 0;
assign Check_Bit[518] = (Bit[518] == 1) ? 1 : 0;
assign Check_Bit[519] = (Bit[519] == 0) ? 1 : 0;
assign Check_Bit[520] = (Bit[520] == 1) ? 1 : 0;
assign Check_Bit[521] = (Bit[521] == 0) ? 1 : 0;
assign Check_Bit[522] = (Bit[522] == 1) ? 1 : 0;
assign Check_Bit[523] = (Bit[523] == 0) ? 1 : 0;
assign Check_Bit[524] = (Bit[524] == 0) ? 1 : 0;
assign Check_Bit[525] = (Bit[525] == 0) ? 1 : 0;
assign Check_Bit[526] = (Bit[526] == 0) ? 1 : 0;
assign Check_Bit[527] = (Bit[527] == 1) ? 1 : 0;
assign Check_Bit[528] = (Bit[528] == 1) ? 1 : 0;
assign Check_Bit[529] = (Bit[529] == 0) ? 1 : 0;
assign Check_Bit[530] = (Bit[530] == 1) ? 1 : 0;
assign Check_Bit[531] = (Bit[531] == 0) ? 1 : 0;
assign Check_Bit[532] = (Bit[532] == 1) ? 1 : 0;
assign Check_Bit[533] = (Bit[533] == 1) ? 1 : 0;
assign Check_Bit[534] = (Bit[534] == 0) ? 1 : 0;
assign Check_Bit[535] = (Bit[535] == 1) ? 1 : 0;
assign Check_Bit[536] = (Bit[536] == 0) ? 1 : 0;
assign Check_Bit[537] = (Bit[537] == 1) ? 1 : 0;
assign Check_Bit[538] = (Bit[538] == 1) ? 1 : 0;
assign Check_Bit[539] = (Bit[539] == 1) ? 1 : 0;
assign Check_Bit[540] = (Bit[540] == 0) ? 1 : 0;
assign Check_Bit[541] = (Bit[541] == 1) ? 1 : 0;
assign Check_Bit[542] = (Bit[542] == 1) ? 1 : 0;
assign Check_Bit[543] = (Bit[543] == 0) ? 1 : 0;
assign Check_Bit[544] = (Bit[544] == 0) ? 1 : 0;
assign Check_Bit[545] = (Bit[545] == 1) ? 1 : 0;
assign Check_Bit[546] = (Bit[546] == 0) ? 1 : 0;
assign Check_Bit[547] = (Bit[547] == 0) ? 1 : 0;
assign Check_Bit[548] = (Bit[548] == 0) ? 1 : 0;
assign Check_Bit[549] = (Bit[549] == 0) ? 1 : 0;
assign Check_Bit[550] = (Bit[550] == 0) ? 1 : 0;
assign Check_Bit[551] = (Bit[551] == 1) ? 1 : 0;
assign Check_Bit[552] = (Bit[552] == 0) ? 1 : 0;
assign Check_Bit[553] = (Bit[553] == 1) ? 1 : 0;
assign Check_Bit[554] = (Bit[554] == 1) ? 1 : 0;
assign Check_Bit[555] = (Bit[555] == 1) ? 1 : 0;
assign Check_Bit[556] = (Bit[556] == 1) ? 1 : 0;
assign Check_Bit[557] = (Bit[557] == 0) ? 1 : 0;
assign Check_Bit[558] = (Bit[558] == 0) ? 1 : 0;
assign Check_Bit[559] = (Bit[559] == 1) ? 1 : 0;
assign Check_Bit[560] = (Bit[560] == 1) ? 1 : 0;
assign Check_Bit[561] = (Bit[561] == 0) ? 1 : 0;
assign Check_Bit[562] = (Bit[562] == 0) ? 1 : 0;
assign Check_Bit[563] = (Bit[563] == 1) ? 1 : 0;
assign Check_Bit[564] = (Bit[564] == 0) ? 1 : 0;
assign Check_Bit[565] = (Bit[565] == 1) ? 1 : 0;
assign Check_Bit[566] = (Bit[566] == 1) ? 1 : 0;
assign Check_Bit[567] = (Bit[567] == 0) ? 1 : 0;
assign Check_Bit[568] = (Bit[568] == 0) ? 1 : 0;
assign Check_Bit[569] = (Bit[569] == 1) ? 1 : 0;
assign Check_Bit[570] = (Bit[570] == 0) ? 1 : 0;
assign Check_Bit[571] = (Bit[571] == 1) ? 1 : 0;
assign Check_Bit[572] = (Bit[572] == 1) ? 1 : 0;
assign Check_Bit[573] = (Bit[573] == 0) ? 1 : 0;
assign Check_Bit[574] = (Bit[574] == 0) ? 1 : 0;
assign Check_Bit[575] = (Bit[575] == 1) ? 1 : 0;
assign Check_Bit[576] = (Bit[576] == 1) ? 1 : 0;
assign Check_Bit[577] = (Bit[577] == 1) ? 1 : 0;
assign Check_Bit[578] = (Bit[578] == 0) ? 1 : 0;
assign Check_Bit[579] = (Bit[579] == 0) ? 1 : 0;
assign Check_Bit[580] = (Bit[580] == 1) ? 1 : 0;
assign Check_Bit[581] = (Bit[581] == 1) ? 1 : 0;
assign Check_Bit[582] = (Bit[582] == 1) ? 1 : 0;
assign Check_Bit[583] = (Bit[583] == 1) ? 1 : 0;
assign Check_Bit[584] = (Bit[584] == 0) ? 1 : 0;
assign Check_Bit[585] = (Bit[585] == 0) ? 1 : 0;
assign Check_Bit[586] = (Bit[586] == 1) ? 1 : 0;
assign Check_Bit[587] = (Bit[587] == 0) ? 1 : 0;
assign Check_Bit[588] = (Bit[588] == 0) ? 1 : 0;
assign Check_Bit[589] = (Bit[589] == 1) ? 1 : 0;
assign Check_Bit[590] = (Bit[590] == 1) ? 1 : 0;
assign Check_Bit[591] = (Bit[591] == 0) ? 1 : 0;
assign Check_Bit[592] = (Bit[592] == 0) ? 1 : 0;
assign Check_Bit[593] = (Bit[593] == 1) ? 1 : 0;
assign Check_Bit[594] = (Bit[594] == 0) ? 1 : 0;
assign Check_Bit[595] = (Bit[595] == 1) ? 1 : 0;
assign Check_Bit[596] = (Bit[596] == 1) ? 1 : 0;
assign Check_Bit[597] = (Bit[597] == 0) ? 1 : 0;
assign Check_Bit[598] = (Bit[598] == 1) ? 1 : 0;
assign Check_Bit[599] = (Bit[599] == 1) ? 1 : 0;
assign Check_Bit[600] = (Bit[600] == 1) ? 1 : 0;
assign Check_Bit[601] = (Bit[601] == 0) ? 1 : 0;
assign Check_Bit[602] = (Bit[602] == 1) ? 1 : 0;
assign Check_Bit[603] = (Bit[603] == 1) ? 1 : 0;
assign Check_Bit[604] = (Bit[604] == 1) ? 1 : 0;
assign Check_Bit[605] = (Bit[605] == 1) ? 1 : 0;
assign Check_Bit[606] = (Bit[606] == 0) ? 1 : 0;
assign Check_Bit[607] = (Bit[607] == 1) ? 1 : 0;
assign Check_Bit[608] = (Bit[608] == 1) ? 1 : 0;
assign Check_Bit[609] = (Bit[609] == 0) ? 1 : 0;
assign Check_Bit[610] = (Bit[610] == 0) ? 1 : 0;
assign Check_Bit[611] = (Bit[611] == 1) ? 1 : 0;
assign Check_Bit[612] = (Bit[612] == 1) ? 1 : 0;
assign Check_Bit[613] = (Bit[613] == 1) ? 1 : 0;
assign Check_Bit[614] = (Bit[614] == 1) ? 1 : 0;
assign Check_Bit[615] = (Bit[615] == 1) ? 1 : 0;
assign Check_Bit[616] = (Bit[616] == 0) ? 1 : 0;
assign Check_Bit[617] = (Bit[617] == 1) ? 1 : 0;
assign Check_Bit[618] = (Bit[618] == 1) ? 1 : 0;
assign Check_Bit[619] = (Bit[619] == 0) ? 1 : 0;
assign Check_Bit[620] = (Bit[620] == 0) ? 1 : 0;
assign Check_Bit[621] = (Bit[621] == 0) ? 1 : 0;
assign Check_Bit[622] = (Bit[622] == 0) ? 1 : 0;
assign Check_Bit[623] = (Bit[623] == 0) ? 1 : 0;
assign Check_Bit[624] = (Bit[624] == 0) ? 1 : 0;
assign Check_Bit[625] = (Bit[625] == 0) ? 1 : 0;
assign Check_Bit[626] = (Bit[626] == 1) ? 1 : 0;
assign Check_Bit[627] = (Bit[627] == 1) ? 1 : 0;
assign Check_Bit[628] = (Bit[628] == 0) ? 1 : 0;
assign Check_Bit[629] = (Bit[629] == 0) ? 1 : 0;
assign Check_Bit[630] = (Bit[630] == 1) ? 1 : 0;
assign Check_Bit[631] = (Bit[631] == 0) ? 1 : 0;
assign Check_Bit[632] = (Bit[632] == 1) ? 1 : 0;
assign Check_Bit[633] = (Bit[633] == 1) ? 1 : 0;
assign Check_Bit[634] = (Bit[634] == 1) ? 1 : 0;
assign Check_Bit[635] = (Bit[635] == 0) ? 1 : 0;
assign Check_Bit[636] = (Bit[636] == 1) ? 1 : 0;
assign Check_Bit[637] = (Bit[637] == 0) ? 1 : 0;
assign Check_Bit[638] = (Bit[638] == 0) ? 1 : 0;
assign Check_Bit[639] = (Bit[639] == 0) ? 1 : 0;
assign Check_Bit[640] = (Bit[640] == 1) ? 1 : 0;
assign Check_Bit[641] = (Bit[641] == 1) ? 1 : 0;
assign Check_Bit[642] = (Bit[642] == 0) ? 1 : 0;
assign Check_Bit[643] = (Bit[643] == 1) ? 1 : 0;
assign Check_Bit[644] = (Bit[644] == 0) ? 1 : 0;
assign Check_Bit[645] = (Bit[645] == 0) ? 1 : 0;
assign Check_Bit[646] = (Bit[646] == 0) ? 1 : 0;
assign Check_Bit[647] = (Bit[647] == 0) ? 1 : 0;
assign Check_Bit[648] = (Bit[648] == 1) ? 1 : 0;
assign Check_Bit[649] = (Bit[649] == 0) ? 1 : 0;
assign Check_Bit[650] = (Bit[650] == 1) ? 1 : 0;
assign Check_Bit[651] = (Bit[651] == 0) ? 1 : 0;
assign Check_Bit[652] = (Bit[652] == 0) ? 1 : 0;
assign Check_Bit[653] = (Bit[653] == 1) ? 1 : 0;
assign Check_Bit[654] = (Bit[654] == 1) ? 1 : 0;
assign Check_Bit[655] = (Bit[655] == 0) ? 1 : 0;
assign Check_Bit[656] = (Bit[656] == 0) ? 1 : 0;
assign Check_Bit[657] = (Bit[657] == 1) ? 1 : 0;
assign Check_Bit[658] = (Bit[658] == 1) ? 1 : 0;
assign Check_Bit[659] = (Bit[659] == 0) ? 1 : 0;
assign Check_Bit[660] = (Bit[660] == 0) ? 1 : 0;
assign Check_Bit[661] = (Bit[661] == 0) ? 1 : 0;
assign Check_Bit[662] = (Bit[662] == 1) ? 1 : 0;
assign Check_Bit[663] = (Bit[663] == 1) ? 1 : 0;
assign Check_Bit[664] = (Bit[664] == 0) ? 1 : 0;
assign Check_Bit[665] = (Bit[665] == 1) ? 1 : 0;
assign Check_Bit[666] = (Bit[666] == 0) ? 1 : 0;
assign Check_Bit[667] = (Bit[667] == 0) ? 1 : 0;
assign Check_Bit[668] = (Bit[668] == 0) ? 1 : 0;
assign Check_Bit[669] = (Bit[669] == 0) ? 1 : 0;
assign Check_Bit[670] = (Bit[670] == 1) ? 1 : 0;
assign Check_Bit[671] = (Bit[671] == 0) ? 1 : 0;
assign Check_Bit[672] = (Bit[672] == 1) ? 1 : 0;
assign Check_Bit[673] = (Bit[673] == 0) ? 1 : 0;
assign Check_Bit[674] = (Bit[674] == 1) ? 1 : 0;
assign Check_Bit[675] = (Bit[675] == 0) ? 1 : 0;
assign Check_Bit[676] = (Bit[676] == 0) ? 1 : 0;
assign Check_Bit[677] = (Bit[677] == 0) ? 1 : 0;
assign Check_Bit[678] = (Bit[678] == 0) ? 1 : 0;
assign Check_Bit[679] = (Bit[679] == 1) ? 1 : 0;
assign Check_Bit[680] = (Bit[680] == 1) ? 1 : 0;
assign Check_Bit[681] = (Bit[681] == 1) ? 1 : 0;
assign Check_Bit[682] = (Bit[682] == 0) ? 1 : 0;
assign Check_Bit[683] = (Bit[683] == 0) ? 1 : 0;
assign Check_Bit[684] = (Bit[684] == 1) ? 1 : 0;
assign Check_Bit[685] = (Bit[685] == 0) ? 1 : 0;
assign Check_Bit[686] = (Bit[686] == 0) ? 1 : 0;
assign Check_Bit[687] = (Bit[687] == 0) ? 1 : 0;
assign Check_Bit[688] = (Bit[688] == 0) ? 1 : 0;
assign Check_Bit[689] = (Bit[689] == 0) ? 1 : 0;
assign Check_Bit[690] = (Bit[690] == 1) ? 1 : 0;
assign Check_Bit[691] = (Bit[691] == 1) ? 1 : 0;
assign Check_Bit[692] = (Bit[692] == 0) ? 1 : 0;
assign Check_Bit[693] = (Bit[693] == 1) ? 1 : 0;
assign Check_Bit[694] = (Bit[694] == 0) ? 1 : 0;
assign Check_Bit[695] = (Bit[695] == 0) ? 1 : 0;
assign Check_Bit[696] = (Bit[696] == 0) ? 1 : 0;
assign Check_Bit[697] = (Bit[697] == 0) ? 1 : 0;
assign Check_Bit[698] = (Bit[698] == 0) ? 1 : 0;
assign Check_Bit[699] = (Bit[699] == 0) ? 1 : 0;
assign Check_Bit[700] = (Bit[700] == 1) ? 1 : 0;
assign Check_Bit[701] = (Bit[701] == 0) ? 1 : 0;
assign Check_Bit[702] = (Bit[702] == 1) ? 1 : 0;
assign Check_Bit[703] = (Bit[703] == 1) ? 1 : 0;
assign Check_Bit[704] = (Bit[704] == 0) ? 1 : 0;
assign Check_Bit[705] = (Bit[705] == 0) ? 1 : 0;
assign Check_Bit[706] = (Bit[706] == 0) ? 1 : 0;
assign Check_Bit[707] = (Bit[707] == 0) ? 1 : 0;
assign Check_Bit[708] = (Bit[708] == 1) ? 1 : 0;
assign Check_Bit[709] = (Bit[709] == 1) ? 1 : 0;
assign Check_Bit[710] = (Bit[710] == 0) ? 1 : 0;
assign Check_Bit[711] = (Bit[711] == 1) ? 1 : 0;
assign Check_Bit[712] = (Bit[712] == 0) ? 1 : 0;
assign Check_Bit[713] = (Bit[713] == 1) ? 1 : 0;
assign Check_Bit[714] = (Bit[714] == 0) ? 1 : 0;
assign Check_Bit[715] = (Bit[715] == 1) ? 1 : 0;
assign Check_Bit[716] = (Bit[716] == 1) ? 1 : 0;
assign Check_Bit[717] = (Bit[717] == 1) ? 1 : 0;
assign Check_Bit[718] = (Bit[718] == 0) ? 1 : 0;
assign Check_Bit[719] = (Bit[719] == 0) ? 1 : 0;
assign Check_Bit[720] = (Bit[720] == 0) ? 1 : 0;
assign Check_Bit[721] = (Bit[721] == 1) ? 1 : 0;
assign Check_Bit[722] = (Bit[722] == 1) ? 1 : 0;
assign Check_Bit[723] = (Bit[723] == 1) ? 1 : 0;
assign Check_Bit[724] = (Bit[724] == 0) ? 1 : 0;
assign Check_Bit[725] = (Bit[725] == 0) ? 1 : 0;
assign Check_Bit[726] = (Bit[726] == 0) ? 1 : 0;
assign Check_Bit[727] = (Bit[727] == 0) ? 1 : 0;
assign Check_Bit[728] = (Bit[728] == 1) ? 1 : 0;
assign Check_Bit[729] = (Bit[729] == 0) ? 1 : 0;
assign Check_Bit[730] = (Bit[730] == 0) ? 1 : 0;
assign Check_Bit[731] = (Bit[731] == 0) ? 1 : 0;
assign Check_Bit[732] = (Bit[732] == 1) ? 1 : 0;
assign Check_Bit[733] = (Bit[733] == 1) ? 1 : 0;
assign Check_Bit[734] = (Bit[734] == 0) ? 1 : 0;
assign Check_Bit[735] = (Bit[735] == 1) ? 1 : 0;
assign Check_Bit[736] = (Bit[736] == 1) ? 1 : 0;
assign Check_Bit[737] = (Bit[737] == 0) ? 1 : 0;
assign Check_Bit[738] = (Bit[738] == 0) ? 1 : 0;
assign Check_Bit[739] = (Bit[739] == 1) ? 1 : 0;
assign Check_Bit[740] = (Bit[740] == 0) ? 1 : 0;
assign Check_Bit[741] = (Bit[741] == 1) ? 1 : 0;
assign Check_Bit[742] = (Bit[742] == 0) ? 1 : 0;
assign Check_Bit[743] = (Bit[743] == 1) ? 1 : 0;
assign Check_Bit[744] = (Bit[744] == 0) ? 1 : 0;
assign Check_Bit[745] = (Bit[745] == 0) ? 1 : 0;
assign Check_Bit[746] = (Bit[746] == 1) ? 1 : 0;
assign Check_Bit[747] = (Bit[747] == 0) ? 1 : 0;
assign Check_Bit[748] = (Bit[748] == 1) ? 1 : 0;
assign Check_Bit[749] = (Bit[749] == 1) ? 1 : 0;
assign Check_Bit[750] = (Bit[750] == 1) ? 1 : 0;
assign Check_Bit[751] = (Bit[751] == 1) ? 1 : 0;
assign Check_Bit[752] = (Bit[752] == 0) ? 1 : 0;
assign Check_Bit[753] = (Bit[753] == 1) ? 1 : 0;
assign Check_Bit[754] = (Bit[754] == 1) ? 1 : 0;
assign Check_Bit[755] = (Bit[755] == 0) ? 1 : 0;
assign Check_Bit[756] = (Bit[756] == 0) ? 1 : 0;
assign Check_Bit[757] = (Bit[757] == 0) ? 1 : 0;
assign Check_Bit[758] = (Bit[758] == 1) ? 1 : 0;
assign Check_Bit[759] = (Bit[759] == 1) ? 1 : 0;
assign Check_Bit[760] = (Bit[760] == 0) ? 1 : 0;
assign Check_Bit[761] = (Bit[761] == 1) ? 1 : 0;
assign Check_Bit[762] = (Bit[762] == 1) ? 1 : 0;
assign Check_Bit[763] = (Bit[763] == 0) ? 1 : 0;
assign Check_Bit[764] = (Bit[764] == 0) ? 1 : 0;
assign Check_Bit[765] = (Bit[765] == 0) ? 1 : 0;
assign Check_Bit[766] = (Bit[766] == 0) ? 1 : 0;
assign Check_Bit[767] = (Bit[767] == 1) ? 1 : 0;
assign Check_Bit[768] = (Bit[768] == 1) ? 1 : 0;
assign Check_Bit[769] = (Bit[769] == 0) ? 1 : 0;
assign Check_Bit[770] = (Bit[770] == 1) ? 1 : 0;
assign Check_Bit[771] = (Bit[771] == 0) ? 1 : 0;
assign Check_Bit[772] = (Bit[772] == 1) ? 1 : 0;
assign Check_Bit[773] = (Bit[773] == 1) ? 1 : 0;
assign Check_Bit[774] = (Bit[774] == 0) ? 1 : 0;
assign Check_Bit[775] = (Bit[775] == 1) ? 1 : 0;
assign Check_Bit[776] = (Bit[776] == 0) ? 1 : 0;
assign Check_Bit[777] = (Bit[777] == 1) ? 1 : 0;
assign Check_Bit[778] = (Bit[778] == 1) ? 1 : 0;
assign Check_Bit[779] = (Bit[779] == 1) ? 1 : 0;
assign Check_Bit[780] = (Bit[780] == 0) ? 1 : 0;
assign Check_Bit[781] = (Bit[781] == 1) ? 1 : 0;
assign Check_Bit[782] = (Bit[782] == 1) ? 1 : 0;
assign Check_Bit[783] = (Bit[783] == 0) ? 1 : 0;
assign Check_Bit[784] = (Bit[784] == 0) ? 1 : 0;
assign Check_Bit[785] = (Bit[785] == 1) ? 1 : 0;
assign Check_Bit[786] = (Bit[786] == 0) ? 1 : 0;
assign Check_Bit[787] = (Bit[787] == 1) ? 1 : 0;
assign Check_Bit[788] = (Bit[788] == 1) ? 1 : 0;
assign Check_Bit[789] = (Bit[789] == 0) ? 1 : 0;
assign Check_Bit[790] = (Bit[790] == 0) ? 1 : 0;
assign Check_Bit[791] = (Bit[791] == 0) ? 1 : 0;
assign Check_Bit[792] = (Bit[792] == 0) ? 1 : 0;
assign Check_Bit[793] = (Bit[793] == 1) ? 1 : 0;
assign Check_Bit[794] = (Bit[794] == 1) ? 1 : 0;
assign Check_Bit[795] = (Bit[795] == 0) ? 1 : 0;
assign Check_Bit[796] = (Bit[796] == 0) ? 1 : 0;
assign Check_Bit[797] = (Bit[797] == 0) ? 1 : 0;
assign Check_Bit[798] = (Bit[798] == 1) ? 1 : 0;
assign Check_Bit[799] = (Bit[799] == 0) ? 1 : 0;
assign Check_Bit[800] = (Bit[800] == 0) ? 1 : 0;
assign Check_Bit[801] = (Bit[801] == 0) ? 1 : 0;
assign Check_Bit[802] = (Bit[802] == 0) ? 1 : 0;
assign Check_Bit[803] = (Bit[803] == 1) ? 1 : 0;
assign Check_Bit[804] = (Bit[804] == 1) ? 1 : 0;
assign Check_Bit[805] = (Bit[805] == 0) ? 1 : 0;
assign Check_Bit[806] = (Bit[806] == 0) ? 1 : 0;
assign Check_Bit[807] = (Bit[807] == 0) ? 1 : 0;
assign Check_Bit[808] = (Bit[808] == 1) ? 1 : 0;
assign Check_Bit[809] = (Bit[809] == 0) ? 1 : 0;
assign Check_Bit[810] = (Bit[810] == 1) ? 1 : 0;
assign Check_Bit[811] = (Bit[811] == 0) ? 1 : 0;
assign Check_Bit[812] = (Bit[812] == 1) ? 1 : 0;
assign Check_Bit[813] = (Bit[813] == 1) ? 1 : 0;
assign Check_Bit[814] = (Bit[814] == 1) ? 1 : 0;
assign Check_Bit[815] = (Bit[815] == 0) ? 1 : 0;
assign Check_Bit[816] = (Bit[816] == 0) ? 1 : 0;
assign Check_Bit[817] = (Bit[817] == 0) ? 1 : 0;
assign Check_Bit[818] = (Bit[818] == 1) ? 1 : 0;
assign Check_Bit[819] = (Bit[819] == 1) ? 1 : 0;
assign Check_Bit[820] = (Bit[820] == 0) ? 1 : 0;
assign Check_Bit[821] = (Bit[821] == 0) ? 1 : 0;
assign Check_Bit[822] = (Bit[822] == 1) ? 1 : 0;
assign Check_Bit[823] = (Bit[823] == 0) ? 1 : 0;
assign Check_Bit[824] = (Bit[824] == 1) ? 1 : 0;
assign Check_Bit[825] = (Bit[825] == 1) ? 1 : 0;
assign Check_Bit[826] = (Bit[826] == 1) ? 1 : 0;
assign Check_Bit[827] = (Bit[827] == 0) ? 1 : 0;
assign Check_Bit[828] = (Bit[828] == 0) ? 1 : 0;
assign Check_Bit[829] = (Bit[829] == 0) ? 1 : 0;
assign Check_Bit[830] = (Bit[830] == 1) ? 1 : 0;
assign Check_Bit[831] = (Bit[831] == 1) ? 1 : 0;
assign Check_Bit[832] = (Bit[832] == 0) ? 1 : 0;
assign Check_Bit[833] = (Bit[833] == 1) ? 1 : 0;
assign Check_Bit[834] = (Bit[834] == 1) ? 1 : 0;
assign Check_Bit[835] = (Bit[835] == 1) ? 1 : 0;
assign Check_Bit[836] = (Bit[836] == 1) ? 1 : 0;
assign Check_Bit[837] = (Bit[837] == 0) ? 1 : 0;
assign Check_Bit[838] = (Bit[838] == 1) ? 1 : 0;
assign Check_Bit[839] = (Bit[839] == 0) ? 1 : 0;
assign Check_Bit[840] = (Bit[840] == 0) ? 1 : 0;
assign Check_Bit[841] = (Bit[841] == 0) ? 1 : 0;
assign Check_Bit[842] = (Bit[842] == 1) ? 1 : 0;
assign Check_Bit[843] = (Bit[843] == 1) ? 1 : 0;
assign Check_Bit[844] = (Bit[844] == 0) ? 1 : 0;
assign Check_Bit[845] = (Bit[845] == 1) ? 1 : 0;
assign Check_Bit[846] = (Bit[846] == 1) ? 1 : 0;
assign Check_Bit[847] = (Bit[847] == 1) ? 1 : 0;
assign Check_Bit[848] = (Bit[848] == 0) ? 1 : 0;
assign Check_Bit[849] = (Bit[849] == 1) ? 1 : 0;
assign Check_Bit[850] = (Bit[850] == 0) ? 1 : 0;
assign Check_Bit[851] = (Bit[851] == 0) ? 1 : 0;
assign Check_Bit[852] = (Bit[852] == 1) ? 1 : 0;
assign Check_Bit[853] = (Bit[853] == 0) ? 1 : 0;
assign Check_Bit[854] = (Bit[854] == 1) ? 1 : 0;
assign Check_Bit[855] = (Bit[855] == 0) ? 1 : 0;
assign Check_Bit[856] = (Bit[856] == 0) ? 1 : 0;
assign Check_Bit[857] = (Bit[857] == 1) ? 1 : 0;
assign Check_Bit[858] = (Bit[858] == 1) ? 1 : 0;
assign Check_Bit[859] = (Bit[859] == 1) ? 1 : 0;
assign Check_Bit[860] = (Bit[860] == 1) ? 1 : 0;
assign Check_Bit[861] = (Bit[861] == 1) ? 1 : 0;
assign Check_Bit[862] = (Bit[862] == 1) ? 1 : 0;
assign Check_Bit[863] = (Bit[863] == 1) ? 1 : 0;
assign Check_Bit[864] = (Bit[864] == 0) ? 1 : 0;
assign Check_Bit[865] = (Bit[865] == 0) ? 1 : 0;
assign Check_Bit[866] = (Bit[866] == 0) ? 1 : 0;
assign Check_Bit[867] = (Bit[867] == 1) ? 1 : 0;
assign Check_Bit[868] = (Bit[868] == 1) ? 1 : 0;
assign Check_Bit[869] = (Bit[869] == 0) ? 1 : 0;
assign Check_Bit[870] = (Bit[870] == 0) ? 1 : 0;
assign Check_Bit[871] = (Bit[871] == 1) ? 1 : 0;
assign Check_Bit[872] = (Bit[872] == 1) ? 1 : 0;
assign Check_Bit[873] = (Bit[873] == 1) ? 1 : 0;
assign Check_Bit[874] = (Bit[874] == 1) ? 1 : 0;
assign Check_Bit[875] = (Bit[875] == 0) ? 1 : 0;
assign Check_Bit[876] = (Bit[876] == 1) ? 1 : 0;
assign Check_Bit[877] = (Bit[877] == 0) ? 1 : 0;
assign Check_Bit[878] = (Bit[878] == 1) ? 1 : 0;
assign Check_Bit[879] = (Bit[879] == 0) ? 1 : 0;
assign Check_Bit[880] = (Bit[880] == 1) ? 1 : 0;
assign Check_Bit[881] = (Bit[881] == 1) ? 1 : 0;
assign Check_Bit[882] = (Bit[882] == 0) ? 1 : 0;
assign Check_Bit[883] = (Bit[883] == 0) ? 1 : 0;
assign Check_Bit[884] = (Bit[884] == 1) ? 1 : 0;
assign Check_Bit[885] = (Bit[885] == 1) ? 1 : 0;
assign Check_Bit[886] = (Bit[886] == 1) ? 1 : 0;
assign Check_Bit[887] = (Bit[887] == 1) ? 1 : 0;
assign Check_Bit[888] = (Bit[888] == 0) ? 1 : 0;
assign Check_Bit[889] = (Bit[889] == 0) ? 1 : 0;
assign Check_Bit[890] = (Bit[890] == 1) ? 1 : 0;
assign Check_Bit[891] = (Bit[891] == 1) ? 1 : 0;
assign Check_Bit[892] = (Bit[892] == 1) ? 1 : 0;
assign Check_Bit[893] = (Bit[893] == 0) ? 1 : 0;
assign Check_Bit[894] = (Bit[894] == 0) ? 1 : 0;
assign Check_Bit[895] = (Bit[895] == 1) ? 1 : 0;
assign Check_Bit[896] = (Bit[896] == 1) ? 1 : 0;
assign Check_Bit[897] = (Bit[897] == 1) ? 1 : 0;
assign Check_Bit[898] = (Bit[898] == 0) ? 1 : 0;
assign Check_Bit[899] = (Bit[899] == 0) ? 1 : 0;
assign Check_Bit[900] = (Bit[900] == 0) ? 1 : 0;
assign Check_Bit[901] = (Bit[901] == 1) ? 1 : 0;
assign Check_Bit[902] = (Bit[902] == 1) ? 1 : 0;
assign Check_Bit[903] = (Bit[903] == 0) ? 1 : 0;
assign Check_Bit[904] = (Bit[904] == 0) ? 1 : 0;
assign Check_Bit[905] = (Bit[905] == 1) ? 1 : 0;
assign Check_Bit[906] = (Bit[906] == 0) ? 1 : 0;
assign Check_Bit[907] = (Bit[907] == 1) ? 1 : 0;
assign Check_Bit[908] = (Bit[908] == 1) ? 1 : 0;
assign Check_Bit[909] = (Bit[909] == 1) ? 1 : 0;
assign Check_Bit[910] = (Bit[910] == 1) ? 1 : 0;
assign Check_Bit[911] = (Bit[911] == 0) ? 1 : 0;
assign Check_Bit[912] = (Bit[912] == 0) ? 1 : 0;
assign Check_Bit[913] = (Bit[913] == 0) ? 1 : 0;
assign Check_Bit[914] = (Bit[914] == 1) ? 1 : 0;
assign Check_Bit[915] = (Bit[915] == 1) ? 1 : 0;
assign Check_Bit[916] = (Bit[916] == 0) ? 1 : 0;
assign Check_Bit[917] = (Bit[917] == 1) ? 1 : 0;
assign Check_Bit[918] = (Bit[918] == 1) ? 1 : 0;
assign Check_Bit[919] = (Bit[919] == 0) ? 1 : 0;
assign Check_Bit[920] = (Bit[920] == 0) ? 1 : 0;
assign Check_Bit[921] = (Bit[921] == 1) ? 1 : 0;
assign Check_Bit[922] = (Bit[922] == 1) ? 1 : 0;
assign Check_Bit[923] = (Bit[923] == 1) ? 1 : 0;
assign Check_Bit[924] = (Bit[924] == 1) ? 1 : 0;
assign Check_Bit[925] = (Bit[925] == 0) ? 1 : 0;
assign Check_Bit[926] = (Bit[926] == 0) ? 1 : 0;
assign Check_Bit[927] = (Bit[927] == 0) ? 1 : 0;
assign Check_Bit[928] = (Bit[928] == 1) ? 1 : 0;
assign Check_Bit[929] = (Bit[929] == 1) ? 1 : 0;
assign Check_Bit[930] = (Bit[930] == 0) ? 1 : 0;
assign Check_Bit[931] = (Bit[931] == 1) ? 1 : 0;
assign Check_Bit[932] = (Bit[932] == 1) ? 1 : 0;
assign Check_Bit[933] = (Bit[933] == 1) ? 1 : 0;
assign Check_Bit[934] = (Bit[934] == 1) ? 1 : 0;
assign Check_Bit[935] = (Bit[935] == 0) ? 1 : 0;
assign Check_Bit[936] = (Bit[936] == 0) ? 1 : 0;
assign Check_Bit[937] = (Bit[937] == 1) ? 1 : 0;
assign Check_Bit[938] = (Bit[938] == 0) ? 1 : 0;
assign Check_Bit[939] = (Bit[939] == 0) ? 1 : 0;
assign Check_Bit[940] = (Bit[940] == 0) ? 1 : 0;
assign Check_Bit[941] = (Bit[941] == 0) ? 1 : 0;
assign Check_Bit[942] = (Bit[942] == 1) ? 1 : 0;
assign Check_Bit[943] = (Bit[943] == 0) ? 1 : 0;
assign Check_Bit[944] = (Bit[944] == 1) ? 1 : 0;
assign Check_Bit[945] = (Bit[945] == 1) ? 1 : 0;
assign Check_Bit[946] = (Bit[946] == 1) ? 1 : 0;
assign Check_Bit[947] = (Bit[947] == 0) ? 1 : 0;
assign Check_Bit[948] = (Bit[948] == 0) ? 1 : 0;
assign Check_Bit[949] = (Bit[949] == 1) ? 1 : 0;
assign Check_Bit[950] = (Bit[950] == 0) ? 1 : 0;
assign Check_Bit[951] = (Bit[951] == 0) ? 1 : 0;
assign Check_Bit[952] = (Bit[952] == 0) ? 1 : 0;
assign Check_Bit[953] = (Bit[953] == 0) ? 1 : 0;
assign Check_Bit[954] = (Bit[954] == 0) ? 1 : 0;
assign Check_Bit[955] = (Bit[955] == 1) ? 1 : 0;
assign Check_Bit[956] = (Bit[956] == 0) ? 1 : 0;
assign Check_Bit[957] = (Bit[957] == 1) ? 1 : 0;
assign Check_Bit[958] = (Bit[958] == 0) ? 1 : 0;
assign Check_Bit[959] = (Bit[959] == 0) ? 1 : 0;
assign Check_Bit[960] = (Bit[960] == 0) ? 1 : 0;
assign Check_Bit[961] = (Bit[961] == 1) ? 1 : 0;
assign Check_Bit[962] = (Bit[962] == 1) ? 1 : 0;
assign Check_Bit[963] = (Bit[963] == 0) ? 1 : 0;
assign Check_Bit[964] = (Bit[964] == 1) ? 1 : 0;
assign Check_Bit[965] = (Bit[965] == 1) ? 1 : 0;
assign Check_Bit[966] = (Bit[966] == 1) ? 1 : 0;
assign Check_Bit[967] = (Bit[967] == 0) ? 1 : 0;
assign Check_Bit[968] = (Bit[968] == 1) ? 1 : 0;
assign Check_Bit[969] = (Bit[969] == 1) ? 1 : 0;
assign Check_Bit[970] = (Bit[970] == 0) ? 1 : 0;
assign Check_Bit[971] = (Bit[971] == 1) ? 1 : 0;
assign Check_Bit[972] = (Bit[972] == 0) ? 1 : 0;
assign Check_Bit[973] = (Bit[973] == 1) ? 1 : 0;
assign Check_Bit[974] = (Bit[974] == 1) ? 1 : 0;
assign Check_Bit[975] = (Bit[975] == 1) ? 1 : 0;
assign Check_Bit[976] = (Bit[976] == 0) ? 1 : 0;
assign Check_Bit[977] = (Bit[977] == 0) ? 1 : 0;
assign Check_Bit[978] = (Bit[978] == 0) ? 1 : 0;
assign Check_Bit[979] = (Bit[979] == 0) ? 1 : 0;
assign Check_Bit[980] = (Bit[980] == 1) ? 1 : 0;
assign Check_Bit[981] = (Bit[981] == 0) ? 1 : 0;
assign Check_Bit[982] = (Bit[982] == 0) ? 1 : 0;
assign Check_Bit[983] = (Bit[983] == 0) ? 1 : 0;
assign Check_Bit[984] = (Bit[984] == 1) ? 1 : 0;
assign Check_Bit[985] = (Bit[985] == 0) ? 1 : 0;
assign Check_Bit[986] = (Bit[986] == 1) ? 1 : 0;
assign Check_Bit[987] = (Bit[987] == 0) ? 1 : 0;
assign Check_Bit[988] = (Bit[988] == 0) ? 1 : 0;
assign Check_Bit[989] = (Bit[989] == 1) ? 1 : 0;
assign Check_Bit[990] = (Bit[990] == 1) ? 1 : 0;
assign Check_Bit[991] = (Bit[991] == 0) ? 1 : 0;
assign Check_Bit[992] = (Bit[992] == 1) ? 1 : 0;
assign Check_Bit[993] = (Bit[993] == 1) ? 1 : 0;
assign Check_Bit[994] = (Bit[994] == 0) ? 1 : 0;
assign Check_Bit[995] = (Bit[995] == 0) ? 1 : 0;
assign Check_Bit[996] = (Bit[996] == 1) ? 1 : 0;
assign Check_Bit[997] = (Bit[997] == 1) ? 1 : 0;
assign Check_Bit[998] = (Bit[998] == 0) ? 1 : 0;
assign Check_Bit[999] = (Bit[999] == 1) ? 1 : 0;
assign Check_Bit[1000] = (Bit[1000] == 1) ? 1 : 0;
assign Check_Bit[1001] = (Bit[1001] == 1) ? 1 : 0;
assign Check_Bit[1002] = (Bit[1002] == 0) ? 1 : 0;
assign Check_Bit[1003] = (Bit[1003] == 0) ? 1 : 0;
assign Check_Bit[1004] = (Bit[1004] == 1) ? 1 : 0;
assign Check_Bit[1005] = (Bit[1005] == 0) ? 1 : 0;
assign Check_Bit[1006] = (Bit[1006] == 1) ? 1 : 0;
assign Check_Bit[1007] = (Bit[1007] == 0) ? 1 : 0;
assign Check_Bit[1008] = (Bit[1008] == 1) ? 1 : 0;
assign Check_Bit[1009] = (Bit[1009] == 0) ? 1 : 0;
assign Check_Bit[1010] = (Bit[1010] == 0) ? 1 : 0;
assign Check_Bit[1011] = (Bit[1011] == 0) ? 1 : 0;
assign Check_Bit[1012] = (Bit[1012] == 1) ? 1 : 0;
assign Check_Bit[1013] = (Bit[1013] == 1) ? 1 : 0;
assign Check_Bit[1014] = (Bit[1014] == 1) ? 1 : 0;
assign Check_Bit[1015] = (Bit[1015] == 1) ? 1 : 0;
assign Check_Bit[1016] = (Bit[1016] == 1) ? 1 : 0;
assign Check_Bit[1017] = (Bit[1017] == 0) ? 1 : 0;
assign Check_Bit[1018] = (Bit[1018] == 1) ? 1 : 0;
assign Check_Bit[1019] = (Bit[1019] == 0) ? 1 : 0;
assign Check_Bit[1020] = (Bit[1020] == 1) ? 1 : 0;
assign Check_Bit[1021] = (Bit[1021] == 1) ? 1 : 0;
assign Check_Bit[1022] = (Bit[1022] == 1) ? 1 : 0;
assign Check_Bit[1023] = (Bit[1023] == 1) ? 1 : 0;
assign Check_Bit[1024] = (Bit[1024] == 1) ? 1 : 0;
assign Check_Bit[1025] = (Bit[1025] == 0) ? 1 : 0;
assign Check_Bit[1026] = (Bit[1026] == 0) ? 1 : 0;
assign Check_Bit[1027] = (Bit[1027] == 1) ? 1 : 0;
assign Check_Bit[1028] = (Bit[1028] == 0) ? 1 : 0;
assign Check_Bit[1029] = (Bit[1029] == 0) ? 1 : 0;
assign Check_Bit[1030] = (Bit[1030] == 0) ? 1 : 0;
assign Check_Bit[1031] = (Bit[1031] == 1) ? 1 : 0;
assign Check_Bit[1032] = (Bit[1032] == 1) ? 1 : 0;
assign Check_Bit[1033] = (Bit[1033] == 0) ? 1 : 0;
assign Check_Bit[1034] = (Bit[1034] == 0) ? 1 : 0;
assign Check_Bit[1035] = (Bit[1035] == 0) ? 1 : 0;
assign Check_Bit[1036] = (Bit[1036] == 1) ? 1 : 0;
assign Check_Bit[1037] = (Bit[1037] == 1) ? 1 : 0;
assign Check_Bit[1038] = (Bit[1038] == 1) ? 1 : 0;
assign Check_Bit[1039] = (Bit[1039] == 0) ? 1 : 0;
assign Check_Bit[1040] = (Bit[1040] == 1) ? 1 : 0;
assign Check_Bit[1041] = (Bit[1041] == 0) ? 1 : 0;
assign Check_Bit[1042] = (Bit[1042] == 0) ? 1 : 0;
assign Check_Bit[1043] = (Bit[1043] == 1) ? 1 : 0;
assign Check_Bit[1044] = (Bit[1044] == 0) ? 1 : 0;
assign Check_Bit[1045] = (Bit[1045] == 0) ? 1 : 0;
assign Check_Bit[1046] = (Bit[1046] == 1) ? 1 : 0;
assign Check_Bit[1047] = (Bit[1047] == 0) ? 1 : 0;
assign Check_Bit[1048] = (Bit[1048] == 0) ? 1 : 0;
assign Check_Bit[1049] = (Bit[1049] == 0) ? 1 : 0;
assign Check_Bit[1050] = (Bit[1050] == 0) ? 1 : 0;
assign Check_Bit[1051] = (Bit[1051] == 1) ? 1 : 0;
assign Check_Bit[1052] = (Bit[1052] == 1) ? 1 : 0;
assign Check_Bit[1053] = (Bit[1053] == 1) ? 1 : 0;
assign Check_Bit[1054] = (Bit[1054] == 0) ? 1 : 0;
assign Check_Bit[1055] = (Bit[1055] == 0) ? 1 : 0;
assign Check_Bit[1056] = (Bit[1056] == 1) ? 1 : 0;
assign Check_Bit[1057] = (Bit[1057] == 0) ? 1 : 0;
assign Check_Bit[1058] = (Bit[1058] == 1) ? 1 : 0;
assign Check_Bit[1059] = (Bit[1059] == 0) ? 1 : 0;
assign Check_Bit[1060] = (Bit[1060] == 0) ? 1 : 0;
assign Check_Bit[1061] = (Bit[1061] == 0) ? 1 : 0;
assign Check_Bit[1062] = (Bit[1062] == 0) ? 1 : 0;
assign Check_Bit[1063] = (Bit[1063] == 1) ? 1 : 0;
assign Check_Bit[1064] = (Bit[1064] == 0) ? 1 : 0;
assign Check_Bit[1065] = (Bit[1065] == 0) ? 1 : 0;
assign Check_Bit[1066] = (Bit[1066] == 1) ? 1 : 0;
assign Check_Bit[1067] = (Bit[1067] == 0) ? 1 : 0;
assign Check_Bit[1068] = (Bit[1068] == 0) ? 1 : 0;
assign Check_Bit[1069] = (Bit[1069] == 0) ? 1 : 0;
assign Check_Bit[1070] = (Bit[1070] == 1) ? 1 : 0;
assign Check_Bit[1071] = (Bit[1071] == 1) ? 1 : 0;
assign Check_Bit[1072] = (Bit[1072] == 0) ? 1 : 0;
assign Check_Bit[1073] = (Bit[1073] == 0) ? 1 : 0;
assign Check_Bit[1074] = (Bit[1074] == 0) ? 1 : 0;
assign Check_Bit[1075] = (Bit[1075] == 1) ? 1 : 0;
assign Check_Bit[1076] = (Bit[1076] == 0) ? 1 : 0;
assign Check_Bit[1077] = (Bit[1077] == 0) ? 1 : 0;
assign Check_Bit[1078] = (Bit[1078] == 1) ? 1 : 0;
assign Check_Bit[1079] = (Bit[1079] == 0) ? 1 : 0;
assign Check_Bit[1080] = (Bit[1080] == 0) ? 1 : 0;
assign Check_Bit[1081] = (Bit[1081] == 0) ? 1 : 0;
assign Check_Bit[1082] = (Bit[1082] == 0) ? 1 : 0;
assign Check_Bit[1083] = (Bit[1083] == 0) ? 1 : 0;
assign Check_Bit[1084] = (Bit[1084] == 1) ? 1 : 0;
assign Check_Bit[1085] = (Bit[1085] == 0) ? 1 : 0;
assign Check_Bit[1086] = (Bit[1086] == 0) ? 1 : 0;
assign Check_Bit[1087] = (Bit[1087] == 0) ? 1 : 0;
assign Check_Bit[1088] = (Bit[1088] == 1) ? 1 : 0;
assign Check_Bit[1089] = (Bit[1089] == 0) ? 1 : 0;
assign Check_Bit[1090] = (Bit[1090] == 0) ? 1 : 0;
assign Check_Bit[1091] = (Bit[1091] == 1) ? 1 : 0;
assign Check_Bit[1092] = (Bit[1092] == 1) ? 1 : 0;
assign Check_Bit[1093] = (Bit[1093] == 1) ? 1 : 0;
assign Check_Bit[1094] = (Bit[1094] == 1) ? 1 : 0;
assign Check_Bit[1095] = (Bit[1095] == 0) ? 1 : 0;
assign Check_Bit[1096] = (Bit[1096] == 0) ? 1 : 0;
assign Check_Bit[1097] = (Bit[1097] == 0) ? 1 : 0;
assign Check_Bit[1098] = (Bit[1098] == 1) ? 1 : 0;
assign Check_Bit[1099] = (Bit[1099] == 1) ? 1 : 0;
assign Check_Bit[1100] = (Bit[1100] == 1) ? 1 : 0;
assign Check_Bit[1101] = (Bit[1101] == 1) ? 1 : 0;
assign Check_Bit[1102] = (Bit[1102] == 0) ? 1 : 0;
assign Check_Bit[1103] = (Bit[1103] == 1) ? 1 : 0;
assign Check_Bit[1104] = (Bit[1104] == 0) ? 1 : 0;
assign Check_Bit[1105] = (Bit[1105] == 1) ? 1 : 0;
assign Check_Bit[1106] = (Bit[1106] == 1) ? 1 : 0;
assign Check_Bit[1107] = (Bit[1107] == 1) ? 1 : 0;
assign Check_Bit[1108] = (Bit[1108] == 1) ? 1 : 0;
assign Check_Bit[1109] = (Bit[1109] == 0) ? 1 : 0;
assign Check_Bit[1110] = (Bit[1110] == 1) ? 1 : 0;
assign Check_Bit[1111] = (Bit[1111] == 0) ? 1 : 0;
assign Check_Bit[1112] = (Bit[1112] == 1) ? 1 : 0;
assign Check_Bit[1113] = (Bit[1113] == 1) ? 1 : 0;
assign Check_Bit[1114] = (Bit[1114] == 0) ? 1 : 0;
assign Check_Bit[1115] = (Bit[1115] == 1) ? 1 : 0;
assign Check_Bit[1116] = (Bit[1116] == 1) ? 1 : 0;
assign Check_Bit[1117] = (Bit[1117] == 0) ? 1 : 0;
assign Check_Bit[1118] = (Bit[1118] == 0) ? 1 : 0;
assign Check_Bit[1119] = (Bit[1119] == 0) ? 1 : 0;
assign Check_Bit[1120] = (Bit[1120] == 1) ? 1 : 0;
assign Check_Bit[1121] = (Bit[1121] == 1) ? 1 : 0;
assign Check_Bit[1122] = (Bit[1122] == 0) ? 1 : 0;
assign Check_Bit[1123] = (Bit[1123] == 0) ? 1 : 0;
assign Check_Bit[1124] = (Bit[1124] == 1) ? 1 : 0;
assign Check_Bit[1125] = (Bit[1125] == 0) ? 1 : 0;
assign Check_Bit[1126] = (Bit[1126] == 1) ? 1 : 0;
assign Check_Bit[1127] = (Bit[1127] == 1) ? 1 : 0;
assign Check_Bit[1128] = (Bit[1128] == 1) ? 1 : 0;
assign Check_Bit[1129] = (Bit[1129] == 0) ? 1 : 0;
assign Check_Bit[1130] = (Bit[1130] == 0) ? 1 : 0;
assign Check_Bit[1131] = (Bit[1131] == 1) ? 1 : 0;
assign Check_Bit[1132] = (Bit[1132] == 0) ? 1 : 0;
assign Check_Bit[1133] = (Bit[1133] == 1) ? 1 : 0;
assign Check_Bit[1134] = (Bit[1134] == 1) ? 1 : 0;
assign Check_Bit[1135] = (Bit[1135] == 0) ? 1 : 0;
assign Check_Bit[1136] = (Bit[1136] == 1) ? 1 : 0;
assign Check_Bit[1137] = (Bit[1137] == 0) ? 1 : 0;
assign Check_Bit[1138] = (Bit[1138] == 0) ? 1 : 0;
assign Check_Bit[1139] = (Bit[1139] == 1) ? 1 : 0;
assign Check_Bit[1140] = (Bit[1140] == 1) ? 1 : 0;
assign Check_Bit[1141] = (Bit[1141] == 0) ? 1 : 0;
assign Check_Bit[1142] = (Bit[1142] == 0) ? 1 : 0;
assign Check_Bit[1143] = (Bit[1143] == 1) ? 1 : 0;
assign Check_Bit[1144] = (Bit[1144] == 1) ? 1 : 0;
assign Check_Bit[1145] = (Bit[1145] == 0) ? 1 : 0;
assign Check_Bit[1146] = (Bit[1146] == 1) ? 1 : 0;
assign Check_Bit[1147] = (Bit[1147] == 1) ? 1 : 0;
assign Check_Bit[1148] = (Bit[1148] == 0) ? 1 : 0;
assign Check_Bit[1149] = (Bit[1149] == 0) ? 1 : 0;
assign Check_Bit[1150] = (Bit[1150] == 0) ? 1 : 0;
assign Check_Bit[1151] = (Bit[1151] == 1) ? 1 : 0;
assign Check_Bit[1152] = (Bit[1152] == 1) ? 1 : 0;
assign Check_Bit[1153] = (Bit[1153] == 1) ? 1 : 0;
assign Check_Bit[1154] = (Bit[1154] == 1) ? 1 : 0;
assign Check_Bit[1155] = (Bit[1155] == 1) ? 1 : 0;
assign Check_Bit[1156] = (Bit[1156] == 1) ? 1 : 0;
assign Check_Bit[1157] = (Bit[1157] == 1) ? 1 : 0;
assign Check_Bit[1158] = (Bit[1158] == 1) ? 1 : 0;
assign Check_Bit[1159] = (Bit[1159] == 0) ? 1 : 0;
assign Check_Bit[1160] = (Bit[1160] == 1) ? 1 : 0;
assign Check_Bit[1161] = (Bit[1161] == 0) ? 1 : 0;
assign Check_Bit[1162] = (Bit[1162] == 0) ? 1 : 0;
assign Check_Bit[1163] = (Bit[1163] == 1) ? 1 : 0;
assign Check_Bit[1164] = (Bit[1164] == 0) ? 1 : 0;
assign Check_Bit[1165] = (Bit[1165] == 0) ? 1 : 0;
assign Check_Bit[1166] = (Bit[1166] == 0) ? 1 : 0;
assign Check_Bit[1167] = (Bit[1167] == 0) ? 1 : 0;
assign Check_Bit[1168] = (Bit[1168] == 0) ? 1 : 0;
assign Check_Bit[1169] = (Bit[1169] == 1) ? 1 : 0;
assign Check_Bit[1170] = (Bit[1170] == 0) ? 1 : 0;
assign Check_Bit[1171] = (Bit[1171] == 1) ? 1 : 0;
assign Check_Bit[1172] = (Bit[1172] == 0) ? 1 : 0;
assign Check_Bit[1173] = (Bit[1173] == 1) ? 1 : 0;
assign Check_Bit[1174] = (Bit[1174] == 0) ? 1 : 0;
assign Check_Bit[1175] = (Bit[1175] == 0) ? 1 : 0;
assign Check_Bit[1176] = (Bit[1176] == 1) ? 1 : 0;
assign Check_Bit[1177] = (Bit[1177] == 0) ? 1 : 0;
assign Check_Bit[1178] = (Bit[1178] == 0) ? 1 : 0;
assign Check_Bit[1179] = (Bit[1179] == 0) ? 1 : 0;
assign Check_Bit[1180] = (Bit[1180] == 0) ? 1 : 0;
assign Check_Bit[1181] = (Bit[1181] == 1) ? 1 : 0;
assign Check_Bit[1182] = (Bit[1182] == 0) ? 1 : 0;
assign Check_Bit[1183] = (Bit[1183] == 0) ? 1 : 0;
assign Check_Bit[1184] = (Bit[1184] == 1) ? 1 : 0;
assign Check_Bit[1185] = (Bit[1185] == 0) ? 1 : 0;
assign Check_Bit[1186] = (Bit[1186] == 1) ? 1 : 0;
assign Check_Bit[1187] = (Bit[1187] == 1) ? 1 : 0;
assign Check_Bit[1188] = (Bit[1188] == 1) ? 1 : 0;
assign Check_Bit[1189] = (Bit[1189] == 0) ? 1 : 0;
assign Check_Bit[1190] = (Bit[1190] == 1) ? 1 : 0;
assign Check_Bit[1191] = (Bit[1191] == 1) ? 1 : 0;
assign Check_Bit[1192] = (Bit[1192] == 1) ? 1 : 0;
assign Check_Bit[1193] = (Bit[1193] == 0) ? 1 : 0;
assign Check_Bit[1194] = (Bit[1194] == 1) ? 1 : 0;
assign Check_Bit[1195] = (Bit[1195] == 1) ? 1 : 0;
assign Check_Bit[1196] = (Bit[1196] == 1) ? 1 : 0;
assign Check_Bit[1197] = (Bit[1197] == 0) ? 1 : 0;
assign Check_Bit[1198] = (Bit[1198] == 0) ? 1 : 0;
assign Check_Bit[1199] = (Bit[1199] == 0) ? 1 : 0;
assign Check_Bit[1200] = (Bit[1200] == 0) ? 1 : 0;
assign Check_Bit[1201] = (Bit[1201] == 0) ? 1 : 0;
assign Check_Bit[1202] = (Bit[1202] == 1) ? 1 : 0;
assign Check_Bit[1203] = (Bit[1203] == 1) ? 1 : 0;
assign Check_Bit[1204] = (Bit[1204] == 1) ? 1 : 0;
assign Check_Bit[1205] = (Bit[1205] == 0) ? 1 : 0;
assign Check_Bit[1206] = (Bit[1206] == 0) ? 1 : 0;
assign Check_Bit[1207] = (Bit[1207] == 0) ? 1 : 0;
assign Check_Bit[1208] = (Bit[1208] == 1) ? 1 : 0;
assign Check_Bit[1209] = (Bit[1209] == 1) ? 1 : 0;
assign Check_Bit[1210] = (Bit[1210] == 1) ? 1 : 0;
assign Check_Bit[1211] = (Bit[1211] == 0) ? 1 : 0;
assign Check_Bit[1212] = (Bit[1212] == 1) ? 1 : 0;
assign Check_Bit[1213] = (Bit[1213] == 0) ? 1 : 0;
assign Check_Bit[1214] = (Bit[1214] == 1) ? 1 : 0;
assign Check_Bit[1215] = (Bit[1215] == 1) ? 1 : 0;
assign Check_Bit[1216] = (Bit[1216] == 0) ? 1 : 0;
assign Check_Bit[1217] = (Bit[1217] == 1) ? 1 : 0;
assign Check_Bit[1218] = (Bit[1218] == 0) ? 1 : 0;
assign Check_Bit[1219] = (Bit[1219] == 1) ? 1 : 0;
assign Check_Bit[1220] = (Bit[1220] == 1) ? 1 : 0;
assign Check_Bit[1221] = (Bit[1221] == 1) ? 1 : 0;
assign Check_Bit[1222] = (Bit[1222] == 1) ? 1 : 0;
assign Check_Bit[1223] = (Bit[1223] == 0) ? 1 : 0;
assign Check_Bit[1224] = (Bit[1224] == 0) ? 1 : 0;
assign Check_Bit[1225] = (Bit[1225] == 1) ? 1 : 0;
assign Check_Bit[1226] = (Bit[1226] == 1) ? 1 : 0;
assign Check_Bit[1227] = (Bit[1227] == 0) ? 1 : 0;
assign Check_Bit[1228] = (Bit[1228] == 1) ? 1 : 0;
assign Check_Bit[1229] = (Bit[1229] == 0) ? 1 : 0;
assign Check_Bit[1230] = (Bit[1230] == 1) ? 1 : 0;
assign Check_Bit[1231] = (Bit[1231] == 0) ? 1 : 0;
assign Check_Bit[1232] = (Bit[1232] == 1) ? 1 : 0;
assign Check_Bit[1233] = (Bit[1233] == 1) ? 1 : 0;
assign Check_Bit[1234] = (Bit[1234] == 1) ? 1 : 0;
assign Check_Bit[1235] = (Bit[1235] == 1) ? 1 : 0;
assign Check_Bit[1236] = (Bit[1236] == 0) ? 1 : 0;
assign Check_Bit[1237] = (Bit[1237] == 0) ? 1 : 0;
assign Check_Bit[1238] = (Bit[1238] == 1) ? 1 : 0;
assign Check_Bit[1239] = (Bit[1239] == 1) ? 1 : 0;
assign Check_Bit[1240] = (Bit[1240] == 0) ? 1 : 0;
assign Check_Bit[1241] = (Bit[1241] == 0) ? 1 : 0;
assign Check_Bit[1242] = (Bit[1242] == 0) ? 1 : 0;
assign Check_Bit[1243] = (Bit[1243] == 1) ? 1 : 0;
assign Check_Bit[1244] = (Bit[1244] == 1) ? 1 : 0;
assign Check_Bit[1245] = (Bit[1245] == 1) ? 1 : 0;
assign Check_Bit[1246] = (Bit[1246] == 0) ? 1 : 0;
assign Check_Bit[1247] = (Bit[1247] == 0) ? 1 : 0;
assign Check_Bit[1248] = (Bit[1248] == 1) ? 1 : 0;
assign Check_Bit[1249] = (Bit[1249] == 1) ? 1 : 0;
assign Check_Bit[1250] = (Bit[1250] == 1) ? 1 : 0;
assign Check_Bit[1251] = (Bit[1251] == 0) ? 1 : 0;
assign Check_Bit[1252] = (Bit[1252] == 1) ? 1 : 0;
assign Check_Bit[1253] = (Bit[1253] == 1) ? 1 : 0;
assign Check_Bit[1254] = (Bit[1254] == 0) ? 1 : 0;
assign Check_Bit[1255] = (Bit[1255] == 0) ? 1 : 0;
assign Check_Bit[1256] = (Bit[1256] == 1) ? 1 : 0;
assign Check_Bit[1257] = (Bit[1257] == 1) ? 1 : 0;
assign Check_Bit[1258] = (Bit[1258] == 1) ? 1 : 0;
assign Check_Bit[1259] = (Bit[1259] == 1) ? 1 : 0;
assign Check_Bit[1260] = (Bit[1260] == 0) ? 1 : 0;
assign Check_Bit[1261] = (Bit[1261] == 1) ? 1 : 0;
assign Check_Bit[1262] = (Bit[1262] == 1) ? 1 : 0;
assign Check_Bit[1263] = (Bit[1263] == 0) ? 1 : 0;
assign Check_Bit[1264] = (Bit[1264] == 0) ? 1 : 0;
assign Check_Bit[1265] = (Bit[1265] == 1) ? 1 : 0;
assign Check_Bit[1266] = (Bit[1266] == 1) ? 1 : 0;
assign Check_Bit[1267] = (Bit[1267] == 1) ? 1 : 0;
assign Check_Bit[1268] = (Bit[1268] == 0) ? 1 : 0;
assign Check_Bit[1269] = (Bit[1269] == 0) ? 1 : 0;
assign Check_Bit[1270] = (Bit[1270] == 0) ? 1 : 0;
assign Check_Bit[1271] = (Bit[1271] == 0) ? 1 : 0;
assign Check_Bit[1272] = (Bit[1272] == 1) ? 1 : 0;
assign Check_Bit[1273] = (Bit[1273] == 1) ? 1 : 0;
assign Check_Bit[1274] = (Bit[1274] == 1) ? 1 : 0;
assign Check_Bit[1275] = (Bit[1275] == 0) ? 1 : 0;
assign Check_Bit[1276] = (Bit[1276] == 1) ? 1 : 0;
assign Check_Bit[1277] = (Bit[1277] == 0) ? 1 : 0;
assign Check_Bit[1278] = (Bit[1278] == 1) ? 1 : 0;
assign Check_Bit[1279] = (Bit[1279] == 0) ? 1 : 0;
assign Check_Bit[1280] = (Bit[1280] == 1) ? 1 : 0;
assign Check_Bit[1281] = (Bit[1281] == 0) ? 1 : 0;
assign Check_Bit[1282] = (Bit[1282] == 1) ? 1 : 0;
assign Check_Bit[1283] = (Bit[1283] == 1) ? 1 : 0;
assign Check_Bit[1284] = (Bit[1284] == 0) ? 1 : 0;
assign Check_Bit[1285] = (Bit[1285] == 1) ? 1 : 0;
assign Check_Bit[1286] = (Bit[1286] == 1) ? 1 : 0;
assign Check_Bit[1287] = (Bit[1287] == 1) ? 1 : 0;
assign Check_Bit[1288] = (Bit[1288] == 0) ? 1 : 0;
assign Check_Bit[1289] = (Bit[1289] == 1) ? 1 : 0;
assign Check_Bit[1290] = (Bit[1290] == 1) ? 1 : 0;
assign Check_Bit[1291] = (Bit[1291] == 0) ? 1 : 0;
assign Check_Bit[1292] = (Bit[1292] == 0) ? 1 : 0;
assign Check_Bit[1293] = (Bit[1293] == 0) ? 1 : 0;
assign Check_Bit[1294] = (Bit[1294] == 1) ? 1 : 0;
assign Check_Bit[1295] = (Bit[1295] == 1) ? 1 : 0;
assign Check_Bit[1296] = (Bit[1296] == 1) ? 1 : 0;
assign Check_Bit[1297] = (Bit[1297] == 1) ? 1 : 0;
assign Check_Bit[1298] = (Bit[1298] == 0) ? 1 : 0;
assign Check_Bit[1299] = (Bit[1299] == 1) ? 1 : 0;
assign Check_Bit[1300] = (Bit[1300] == 1) ? 1 : 0;
assign Check_Bit[1301] = (Bit[1301] == 0) ? 1 : 0;
assign Check_Bit[1302] = (Bit[1302] == 1) ? 1 : 0;
assign Check_Bit[1303] = (Bit[1303] == 1) ? 1 : 0;
assign Check_Bit[1304] = (Bit[1304] == 1) ? 1 : 0;
assign Check_Bit[1305] = (Bit[1305] == 0) ? 1 : 0;
assign Check_Bit[1306] = (Bit[1306] == 1) ? 1 : 0;
assign Check_Bit[1307] = (Bit[1307] == 0) ? 1 : 0;
assign Check_Bit[1308] = (Bit[1308] == 0) ? 1 : 0;
assign Check_Bit[1309] = (Bit[1309] == 1) ? 1 : 0;
assign Check_Bit[1310] = (Bit[1310] == 0) ? 1 : 0;
assign Check_Bit[1311] = (Bit[1311] == 1) ? 1 : 0;
assign Check_Bit[1312] = (Bit[1312] == 0) ? 1 : 0;
assign Check_Bit[1313] = (Bit[1313] == 0) ? 1 : 0;
assign Check_Bit[1314] = (Bit[1314] == 1) ? 1 : 0;
assign Check_Bit[1315] = (Bit[1315] == 1) ? 1 : 0;
assign Check_Bit[1316] = (Bit[1316] == 0) ? 1 : 0;
assign Check_Bit[1317] = (Bit[1317] == 0) ? 1 : 0;
assign Check_Bit[1318] = (Bit[1318] == 1) ? 1 : 0;
assign Check_Bit[1319] = (Bit[1319] == 1) ? 1 : 0;
assign Check_Bit[1320] = (Bit[1320] == 1) ? 1 : 0;
assign Check_Bit[1321] = (Bit[1321] == 1) ? 1 : 0;
assign Check_Bit[1322] = (Bit[1322] == 0) ? 1 : 0;
assign Check_Bit[1323] = (Bit[1323] == 1) ? 1 : 0;
assign Check_Bit[1324] = (Bit[1324] == 1) ? 1 : 0;
assign Check_Bit[1325] = (Bit[1325] == 1) ? 1 : 0;
assign Check_Bit[1326] = (Bit[1326] == 0) ? 1 : 0;
assign Check_Bit[1327] = (Bit[1327] == 1) ? 1 : 0;
assign Check_Bit[1328] = (Bit[1328] == 1) ? 1 : 0;
assign Check_Bit[1329] = (Bit[1329] == 1) ? 1 : 0;
assign Check_Bit[1330] = (Bit[1330] == 0) ? 1 : 0;
assign Check_Bit[1331] = (Bit[1331] == 1) ? 1 : 0;
assign Check_Bit[1332] = (Bit[1332] == 1) ? 1 : 0;
assign Check_Bit[1333] = (Bit[1333] == 0) ? 1 : 0;
assign Check_Bit[1334] = (Bit[1334] == 1) ? 1 : 0;
assign Check_Bit[1335] = (Bit[1335] == 1) ? 1 : 0;
assign Check_Bit[1336] = (Bit[1336] == 1) ? 1 : 0;
assign Check_Bit[1337] = (Bit[1337] == 0) ? 1 : 0;
assign Check_Bit[1338] = (Bit[1338] == 0) ? 1 : 0;
assign Check_Bit[1339] = (Bit[1339] == 0) ? 1 : 0;
assign Check_Bit[1340] = (Bit[1340] == 1) ? 1 : 0;
assign Check_Bit[1341] = (Bit[1341] == 0) ? 1 : 0;
assign Check_Bit[1342] = (Bit[1342] == 0) ? 1 : 0;
assign Check_Bit[1343] = (Bit[1343] == 0) ? 1 : 0;
assign Check_Bit[1344] = (Bit[1344] == 0) ? 1 : 0;
assign Check_Bit[1345] = (Bit[1345] == 1) ? 1 : 0;
assign Check_Bit[1346] = (Bit[1346] == 1) ? 1 : 0;
assign Check_Bit[1347] = (Bit[1347] == 0) ? 1 : 0;
assign Check_Bit[1348] = (Bit[1348] == 0) ? 1 : 0;
assign Check_Bit[1349] = (Bit[1349] == 0) ? 1 : 0;
assign Check_Bit[1350] = (Bit[1350] == 1) ? 1 : 0;
assign Check_Bit[1351] = (Bit[1351] == 1) ? 1 : 0;
assign Check_Bit[1352] = (Bit[1352] == 1) ? 1 : 0;
assign Check_Bit[1353] = (Bit[1353] == 1) ? 1 : 0;
assign Check_Bit[1354] = (Bit[1354] == 1) ? 1 : 0;
assign Check_Bit[1355] = (Bit[1355] == 0) ? 1 : 0;
assign Check_Bit[1356] = (Bit[1356] == 1) ? 1 : 0;
assign Check_Bit[1357] = (Bit[1357] == 0) ? 1 : 0;
assign Check_Bit[1358] = (Bit[1358] == 0) ? 1 : 0;
assign Check_Bit[1359] = (Bit[1359] == 1) ? 1 : 0;
assign Check_Bit[1360] = (Bit[1360] == 0) ? 1 : 0;
assign Check_Bit[1361] = (Bit[1361] == 1) ? 1 : 0;
assign Check_Bit[1362] = (Bit[1362] == 1) ? 1 : 0;
assign Check_Bit[1363] = (Bit[1363] == 0) ? 1 : 0;
assign Check_Bit[1364] = (Bit[1364] == 0) ? 1 : 0;
assign Check_Bit[1365] = (Bit[1365] == 1) ? 1 : 0;
assign Check_Bit[1366] = (Bit[1366] == 0) ? 1 : 0;
assign Check_Bit[1367] = (Bit[1367] == 0) ? 1 : 0;
assign Check_Bit[1368] = (Bit[1368] == 0) ? 1 : 0;
assign Check_Bit[1369] = (Bit[1369] == 0) ? 1 : 0;
assign Check_Bit[1370] = (Bit[1370] == 1) ? 1 : 0;
assign Check_Bit[1371] = (Bit[1371] == 1) ? 1 : 0;
assign Check_Bit[1372] = (Bit[1372] == 0) ? 1 : 0;
assign Check_Bit[1373] = (Bit[1373] == 1) ? 1 : 0;
assign Check_Bit[1374] = (Bit[1374] == 1) ? 1 : 0;
assign Check_Bit[1375] = (Bit[1375] == 1) ? 1 : 0;
assign Check_Bit[1376] = (Bit[1376] == 0) ? 1 : 0;
assign Check_Bit[1377] = (Bit[1377] == 1) ? 1 : 0;
assign Check_Bit[1378] = (Bit[1378] == 1) ? 1 : 0;
assign Check_Bit[1379] = (Bit[1379] == 0) ? 1 : 0;
assign Check_Bit[1380] = (Bit[1380] == 1) ? 1 : 0;
assign Check_Bit[1381] = (Bit[1381] == 0) ? 1 : 0;
assign Check_Bit[1382] = (Bit[1382] == 0) ? 1 : 0;
assign Check_Bit[1383] = (Bit[1383] == 1) ? 1 : 0;
assign Check_Bit[1384] = (Bit[1384] == 0) ? 1 : 0;
assign Check_Bit[1385] = (Bit[1385] == 1) ? 1 : 0;
assign Check_Bit[1386] = (Bit[1386] == 0) ? 1 : 0;
assign Check_Bit[1387] = (Bit[1387] == 0) ? 1 : 0;
assign Check_Bit[1388] = (Bit[1388] == 1) ? 1 : 0;
assign Check_Bit[1389] = (Bit[1389] == 1) ? 1 : 0;
assign Check_Bit[1390] = (Bit[1390] == 1) ? 1 : 0;
assign Check_Bit[1391] = (Bit[1391] == 0) ? 1 : 0;
assign Check_Bit[1392] = (Bit[1392] == 0) ? 1 : 0;
assign Check_Bit[1393] = (Bit[1393] == 0) ? 1 : 0;
assign Check_Bit[1394] = (Bit[1394] == 1) ? 1 : 0;
assign Check_Bit[1395] = (Bit[1395] == 1) ? 1 : 0;
assign Check_Bit[1396] = (Bit[1396] == 0) ? 1 : 0;
assign Check_Bit[1397] = (Bit[1397] == 1) ? 1 : 0;
assign Check_Bit[1398] = (Bit[1398] == 0) ? 1 : 0;
assign Check_Bit[1399] = (Bit[1399] == 1) ? 1 : 0;
assign Check_Bit[1400] = (Bit[1400] == 1) ? 1 : 0;
assign Check_Bit[1401] = (Bit[1401] == 1) ? 1 : 0;
assign Check_Bit[1402] = (Bit[1402] == 0) ? 1 : 0;
assign Check_Bit[1403] = (Bit[1403] == 0) ? 1 : 0;
assign Check_Bit[1404] = (Bit[1404] == 1) ? 1 : 0;
assign Check_Bit[1405] = (Bit[1405] == 0) ? 1 : 0;
assign Check_Bit[1406] = (Bit[1406] == 0) ? 1 : 0;
assign Check_Bit[1407] = (Bit[1407] == 0) ? 1 : 0;
assign Check_Bit[1408] = (Bit[1408] == 1) ? 1 : 0;
assign Check_Bit[1409] = (Bit[1409] == 1) ? 1 : 0;
assign Check_Bit[1410] = (Bit[1410] == 0) ? 1 : 0;
assign Check_Bit[1411] = (Bit[1411] == 1) ? 1 : 0;
assign Check_Bit[1412] = (Bit[1412] == 1) ? 1 : 0;
assign Check_Bit[1413] = (Bit[1413] == 1) ? 1 : 0;
assign Check_Bit[1414] = (Bit[1414] == 1) ? 1 : 0;
assign Check_Bit[1415] = (Bit[1415] == 1) ? 1 : 0;
assign Check_Bit[1416] = (Bit[1416] == 1) ? 1 : 0;
assign Check_Bit[1417] = (Bit[1417] == 0) ? 1 : 0;
assign Check_Bit[1418] = (Bit[1418] == 0) ? 1 : 0;
assign Check_Bit[1419] = (Bit[1419] == 0) ? 1 : 0;
assign Check_Bit[1420] = (Bit[1420] == 0) ? 1 : 0;
assign Check_Bit[1421] = (Bit[1421] == 0) ? 1 : 0;
assign Check_Bit[1422] = (Bit[1422] == 1) ? 1 : 0;
assign Check_Bit[1423] = (Bit[1423] == 1) ? 1 : 0;
assign Check_Bit[1424] = (Bit[1424] == 0) ? 1 : 0;
assign Check_Bit[1425] = (Bit[1425] == 1) ? 1 : 0;
assign Check_Bit[1426] = (Bit[1426] == 1) ? 1 : 0;
assign Check_Bit[1427] = (Bit[1427] == 1) ? 1 : 0;
assign Check_Bit[1428] = (Bit[1428] == 1) ? 1 : 0;
assign Check_Bit[1429] = (Bit[1429] == 0) ? 1 : 0;
assign Check_Bit[1430] = (Bit[1430] == 0) ? 1 : 0;
assign Check_Bit[1431] = (Bit[1431] == 0) ? 1 : 0;
assign Check_Bit[1432] = (Bit[1432] == 0) ? 1 : 0;
assign Check_Bit[1433] = (Bit[1433] == 1) ? 1 : 0;
assign Check_Bit[1434] = (Bit[1434] == 0) ? 1 : 0;
assign Check_Bit[1435] = (Bit[1435] == 0) ? 1 : 0;
assign Check_Bit[1436] = (Bit[1436] == 0) ? 1 : 0;
assign Check_Bit[1437] = (Bit[1437] == 1) ? 1 : 0;
assign Check_Bit[1438] = (Bit[1438] == 0) ? 1 : 0;
assign Check_Bit[1439] = (Bit[1439] == 0) ? 1 : 0;
wire [63:0] result;
assign result = Check_Bit[0] + Check_Bit[1] + Check_Bit[2] + Check_Bit[3] + Check_Bit[4] + Check_Bit[5] + Check_Bit[6] + Check_Bit[7] + Check_Bit[8] + Check_Bit[9] + Check_Bit[10] + Check_Bit[11] + Check_Bit[12] + Check_Bit[13] + Check_Bit[14] + Check_Bit[15] + Check_Bit[16] + Check_Bit[17] + Check_Bit[18] + Check_Bit[19] + Check_Bit[20] + Check_Bit[21] + Check_Bit[22] + Check_Bit[23] + Check_Bit[24] + Check_Bit[25] + Check_Bit[26] + Check_Bit[27] + Check_Bit[28] + Check_Bit[29] + Check_Bit[30] + Check_Bit[31] + Check_Bit[32] + Check_Bit[33] + Check_Bit[34] + Check_Bit[35] + Check_Bit[36] + Check_Bit[37] + Check_Bit[38] + Check_Bit[39] + Check_Bit[40] + Check_Bit[41] + Check_Bit[42] + Check_Bit[43] + Check_Bit[44] + Check_Bit[45] + Check_Bit[46] + Check_Bit[47] + Check_Bit[48] + Check_Bit[49] + Check_Bit[50] + Check_Bit[51] + Check_Bit[52] + Check_Bit[53] + Check_Bit[54] + Check_Bit[55] + Check_Bit[56] + Check_Bit[57] + Check_Bit[58] + Check_Bit[59] + Check_Bit[60] + Check_Bit[61] + Check_Bit[62] + Check_Bit[63] + Check_Bit[64] + Check_Bit[65] + Check_Bit[66] + Check_Bit[67] + Check_Bit[68] + Check_Bit[69] + Check_Bit[70] + Check_Bit[71] + Check_Bit[72] + Check_Bit[73] + Check_Bit[74] + Check_Bit[75] + Check_Bit[76] + Check_Bit[77] + Check_Bit[78] + Check_Bit[79] + Check_Bit[80] + Check_Bit[81] + Check_Bit[82] + Check_Bit[83] + Check_Bit[84] + Check_Bit[85] + Check_Bit[86] + Check_Bit[87] + Check_Bit[88] + Check_Bit[89] + Check_Bit[90] + Check_Bit[91] + Check_Bit[92] + Check_Bit[93] + Check_Bit[94] + Check_Bit[95] + Check_Bit[96] + Check_Bit[97] + Check_Bit[98] + Check_Bit[99] + Check_Bit[100] + Check_Bit[101] + Check_Bit[102] + Check_Bit[103] + Check_Bit[104] + Check_Bit[105] + Check_Bit[106] + Check_Bit[107] + Check_Bit[108] + Check_Bit[109] + Check_Bit[110] + Check_Bit[111] + Check_Bit[112] + Check_Bit[113] + Check_Bit[114] + Check_Bit[115] + Check_Bit[116] + Check_Bit[117] + Check_Bit[118] + Check_Bit[119] + Check_Bit[120] + Check_Bit[121] + Check_Bit[122] + Check_Bit[123] + Check_Bit[124] + Check_Bit[125] + Check_Bit[126] + Check_Bit[127] + Check_Bit[128] + Check_Bit[129] + Check_Bit[130] + Check_Bit[131] + Check_Bit[132] + Check_Bit[133] + Check_Bit[134] + Check_Bit[135] + Check_Bit[136] + Check_Bit[137] + Check_Bit[138] + Check_Bit[139] + Check_Bit[140] + Check_Bit[141] + Check_Bit[142] + Check_Bit[143] + Check_Bit[144] + Check_Bit[145] + Check_Bit[146] + Check_Bit[147] + Check_Bit[148] + Check_Bit[149] + Check_Bit[150] + Check_Bit[151] + Check_Bit[152] + Check_Bit[153] + Check_Bit[154] + Check_Bit[155] + Check_Bit[156] + Check_Bit[157] + Check_Bit[158] + Check_Bit[159] + Check_Bit[160] + Check_Bit[161] + Check_Bit[162] + Check_Bit[163] + Check_Bit[164] + Check_Bit[165] + Check_Bit[166] + Check_Bit[167] + Check_Bit[168] + Check_Bit[169] + Check_Bit[170] + Check_Bit[171] + Check_Bit[172] + Check_Bit[173] + Check_Bit[174] + Check_Bit[175] + Check_Bit[176] + Check_Bit[177] + Check_Bit[178] + Check_Bit[179] + Check_Bit[180] + Check_Bit[181] + Check_Bit[182] + Check_Bit[183] + Check_Bit[184] + Check_Bit[185] + Check_Bit[186] + Check_Bit[187] + Check_Bit[188] + Check_Bit[189] + Check_Bit[190] + Check_Bit[191] + Check_Bit[192] + Check_Bit[193] + Check_Bit[194] + Check_Bit[195] + Check_Bit[196] + Check_Bit[197] + Check_Bit[198] + Check_Bit[199] + Check_Bit[200] + Check_Bit[201] + Check_Bit[202] + Check_Bit[203] + Check_Bit[204] + Check_Bit[205] + Check_Bit[206] + Check_Bit[207] + Check_Bit[208] + Check_Bit[209] + Check_Bit[210] + Check_Bit[211] + Check_Bit[212] + Check_Bit[213] + Check_Bit[214] + Check_Bit[215] + Check_Bit[216] + Check_Bit[217] + Check_Bit[218] + Check_Bit[219] + Check_Bit[220] + Check_Bit[221] + Check_Bit[222] + Check_Bit[223] + Check_Bit[224] + Check_Bit[225] + Check_Bit[226] + Check_Bit[227] + Check_Bit[228] + Check_Bit[229] + Check_Bit[230] + Check_Bit[231] + Check_Bit[232] + Check_Bit[233] + Check_Bit[234] + Check_Bit[235] + Check_Bit[236] + Check_Bit[237] + Check_Bit[238] + Check_Bit[239] + Check_Bit[240] + Check_Bit[241] + Check_Bit[242] + Check_Bit[243] + Check_Bit[244] + Check_Bit[245] + Check_Bit[246] + Check_Bit[247] + Check_Bit[248] + Check_Bit[249] + Check_Bit[250] + Check_Bit[251] + Check_Bit[252] + Check_Bit[253] + Check_Bit[254] + Check_Bit[255] + Check_Bit[256] + Check_Bit[257] + Check_Bit[258] + Check_Bit[259] + Check_Bit[260] + Check_Bit[261] + Check_Bit[262] + Check_Bit[263] + Check_Bit[264] + Check_Bit[265] + Check_Bit[266] + Check_Bit[267] + Check_Bit[268] + Check_Bit[269] + Check_Bit[270] + Check_Bit[271] + Check_Bit[272] + Check_Bit[273] + Check_Bit[274] + Check_Bit[275] + Check_Bit[276] + Check_Bit[277] + Check_Bit[278] + Check_Bit[279] + Check_Bit[280] + Check_Bit[281] + Check_Bit[282] + Check_Bit[283] + Check_Bit[284] + Check_Bit[285] + Check_Bit[286] + Check_Bit[287] + Check_Bit[288] + Check_Bit[289] + Check_Bit[290] + Check_Bit[291] + Check_Bit[292] + Check_Bit[293] + Check_Bit[294] + Check_Bit[295] + Check_Bit[296] + Check_Bit[297] + Check_Bit[298] + Check_Bit[299] + Check_Bit[300] + Check_Bit[301] + Check_Bit[302] + Check_Bit[303] + Check_Bit[304] + Check_Bit[305] + Check_Bit[306] + Check_Bit[307] + Check_Bit[308] + Check_Bit[309] + Check_Bit[310] + Check_Bit[311] + Check_Bit[312] + Check_Bit[313] + Check_Bit[314] + Check_Bit[315] + Check_Bit[316] + Check_Bit[317] + Check_Bit[318] + Check_Bit[319] + Check_Bit[320] + Check_Bit[321] + Check_Bit[322] + Check_Bit[323] + Check_Bit[324] + Check_Bit[325] + Check_Bit[326] + Check_Bit[327] + Check_Bit[328] + Check_Bit[329] + Check_Bit[330] + Check_Bit[331] + Check_Bit[332] + Check_Bit[333] + Check_Bit[334] + Check_Bit[335] + Check_Bit[336] + Check_Bit[337] + Check_Bit[338] + Check_Bit[339] + Check_Bit[340] + Check_Bit[341] + Check_Bit[342] + Check_Bit[343] + Check_Bit[344] + Check_Bit[345] + Check_Bit[346] + Check_Bit[347] + Check_Bit[348] + Check_Bit[349] + Check_Bit[350] + Check_Bit[351] + Check_Bit[352] + Check_Bit[353] + Check_Bit[354] + Check_Bit[355] + Check_Bit[356] + Check_Bit[357] + Check_Bit[358] + Check_Bit[359] + Check_Bit[360] + Check_Bit[361] + Check_Bit[362] + Check_Bit[363] + Check_Bit[364] + Check_Bit[365] + Check_Bit[366] + Check_Bit[367] + Check_Bit[368] + Check_Bit[369] + Check_Bit[370] + Check_Bit[371] + Check_Bit[372] + Check_Bit[373] + Check_Bit[374] + Check_Bit[375] + Check_Bit[376] + Check_Bit[377] + Check_Bit[378] + Check_Bit[379] + Check_Bit[380] + Check_Bit[381] + Check_Bit[382] + Check_Bit[383] + Check_Bit[384] + Check_Bit[385] + Check_Bit[386] + Check_Bit[387] + Check_Bit[388] + Check_Bit[389] + Check_Bit[390] + Check_Bit[391] + Check_Bit[392] + Check_Bit[393] + Check_Bit[394] + Check_Bit[395] + Check_Bit[396] + Check_Bit[397] + Check_Bit[398] + Check_Bit[399] + Check_Bit[400] + Check_Bit[401] + Check_Bit[402] + Check_Bit[403] + Check_Bit[404] + Check_Bit[405] + Check_Bit[406] + Check_Bit[407] + Check_Bit[408] + Check_Bit[409] + Check_Bit[410] + Check_Bit[411] + Check_Bit[412] + Check_Bit[413] + Check_Bit[414] + Check_Bit[415] + Check_Bit[416] + Check_Bit[417] + Check_Bit[418] + Check_Bit[419] + Check_Bit[420] + Check_Bit[421] + Check_Bit[422] + Check_Bit[423] + Check_Bit[424] + Check_Bit[425] + Check_Bit[426] + Check_Bit[427] + Check_Bit[428] + Check_Bit[429] + Check_Bit[430] + Check_Bit[431] + Check_Bit[432] + Check_Bit[433] + Check_Bit[434] + Check_Bit[435] + Check_Bit[436] + Check_Bit[437] + Check_Bit[438] + Check_Bit[439] + Check_Bit[440] + Check_Bit[441] + Check_Bit[442] + Check_Bit[443] + Check_Bit[444] + Check_Bit[445] + Check_Bit[446] + Check_Bit[447] + Check_Bit[448] + Check_Bit[449] + Check_Bit[450] + Check_Bit[451] + Check_Bit[452] + Check_Bit[453] + Check_Bit[454] + Check_Bit[455] + Check_Bit[456] + Check_Bit[457] + Check_Bit[458] + Check_Bit[459] + Check_Bit[460] + Check_Bit[461] + Check_Bit[462] + Check_Bit[463] + Check_Bit[464] + Check_Bit[465] + Check_Bit[466] + Check_Bit[467] + Check_Bit[468] + Check_Bit[469] + Check_Bit[470] + Check_Bit[471] + Check_Bit[472] + Check_Bit[473] + Check_Bit[474] + Check_Bit[475] + Check_Bit[476] + Check_Bit[477] + Check_Bit[478] + Check_Bit[479] + Check_Bit[480] + Check_Bit[481] + Check_Bit[482] + Check_Bit[483] + Check_Bit[484] + Check_Bit[485] + Check_Bit[486] + Check_Bit[487] + Check_Bit[488] + Check_Bit[489] + Check_Bit[490] + Check_Bit[491] + Check_Bit[492] + Check_Bit[493] + Check_Bit[494] + Check_Bit[495] + Check_Bit[496] + Check_Bit[497] + Check_Bit[498] + Check_Bit[499] + Check_Bit[500] + Check_Bit[501] + Check_Bit[502] + Check_Bit[503] + Check_Bit[504] + Check_Bit[505] + Check_Bit[506] + Check_Bit[507] + Check_Bit[508] + Check_Bit[509] + Check_Bit[510] + Check_Bit[511] + Check_Bit[512] + Check_Bit[513] + Check_Bit[514] + Check_Bit[515] + Check_Bit[516] + Check_Bit[517] + Check_Bit[518] + Check_Bit[519] + Check_Bit[520] + Check_Bit[521] + Check_Bit[522] + Check_Bit[523] + Check_Bit[524] + Check_Bit[525] + Check_Bit[526] + Check_Bit[527] + Check_Bit[528] + Check_Bit[529] + Check_Bit[530] + Check_Bit[531] + Check_Bit[532] + Check_Bit[533] + Check_Bit[534] + Check_Bit[535] + Check_Bit[536] + Check_Bit[537] + Check_Bit[538] + Check_Bit[539] + Check_Bit[540] + Check_Bit[541] + Check_Bit[542] + Check_Bit[543] + Check_Bit[544] + Check_Bit[545] + Check_Bit[546] + Check_Bit[547] + Check_Bit[548] + Check_Bit[549] + Check_Bit[550] + Check_Bit[551] + Check_Bit[552] + Check_Bit[553] + Check_Bit[554] + Check_Bit[555] + Check_Bit[556] + Check_Bit[557] + Check_Bit[558] + Check_Bit[559] + Check_Bit[560] + Check_Bit[561] + Check_Bit[562] + Check_Bit[563] + Check_Bit[564] + Check_Bit[565] + Check_Bit[566] + Check_Bit[567] + Check_Bit[568] + Check_Bit[569] + Check_Bit[570] + Check_Bit[571] + Check_Bit[572] + Check_Bit[573] + Check_Bit[574] + Check_Bit[575] + Check_Bit[576] + Check_Bit[577] + Check_Bit[578] + Check_Bit[579] + Check_Bit[580] + Check_Bit[581] + Check_Bit[582] + Check_Bit[583] + Check_Bit[584] + Check_Bit[585] + Check_Bit[586] + Check_Bit[587] + Check_Bit[588] + Check_Bit[589] + Check_Bit[590] + Check_Bit[591] + Check_Bit[592] + Check_Bit[593] + Check_Bit[594] + Check_Bit[595] + Check_Bit[596] + Check_Bit[597] + Check_Bit[598] + Check_Bit[599] + Check_Bit[600] + Check_Bit[601] + Check_Bit[602] + Check_Bit[603] + Check_Bit[604] + Check_Bit[605] + Check_Bit[606] + Check_Bit[607] + Check_Bit[608] + Check_Bit[609] + Check_Bit[610] + Check_Bit[611] + Check_Bit[612] + Check_Bit[613] + Check_Bit[614] + Check_Bit[615] + Check_Bit[616] + Check_Bit[617] + Check_Bit[618] + Check_Bit[619] + Check_Bit[620] + Check_Bit[621] + Check_Bit[622] + Check_Bit[623] + Check_Bit[624] + Check_Bit[625] + Check_Bit[626] + Check_Bit[627] + Check_Bit[628] + Check_Bit[629] + Check_Bit[630] + Check_Bit[631] + Check_Bit[632] + Check_Bit[633] + Check_Bit[634] + Check_Bit[635] + Check_Bit[636] + Check_Bit[637] + Check_Bit[638] + Check_Bit[639] + Check_Bit[640] + Check_Bit[641] + Check_Bit[642] + Check_Bit[643] + Check_Bit[644] + Check_Bit[645] + Check_Bit[646] + Check_Bit[647] + Check_Bit[648] + Check_Bit[649] + Check_Bit[650] + Check_Bit[651] + Check_Bit[652] + Check_Bit[653] + Check_Bit[654] + Check_Bit[655] + Check_Bit[656] + Check_Bit[657] + Check_Bit[658] + Check_Bit[659] + Check_Bit[660] + Check_Bit[661] + Check_Bit[662] + Check_Bit[663] + Check_Bit[664] + Check_Bit[665] + Check_Bit[666] + Check_Bit[667] + Check_Bit[668] + Check_Bit[669] + Check_Bit[670] + Check_Bit[671] + Check_Bit[672] + Check_Bit[673] + Check_Bit[674] + Check_Bit[675] + Check_Bit[676] + Check_Bit[677] + Check_Bit[678] + Check_Bit[679] + Check_Bit[680] + Check_Bit[681] + Check_Bit[682] + Check_Bit[683] + Check_Bit[684] + Check_Bit[685] + Check_Bit[686] + Check_Bit[687] + Check_Bit[688] + Check_Bit[689] + Check_Bit[690] + Check_Bit[691] + Check_Bit[692] + Check_Bit[693] + Check_Bit[694] + Check_Bit[695] + Check_Bit[696] + Check_Bit[697] + Check_Bit[698] + Check_Bit[699] + Check_Bit[700] + Check_Bit[701] + Check_Bit[702] + Check_Bit[703] + Check_Bit[704] + Check_Bit[705] + Check_Bit[706] + Check_Bit[707] + Check_Bit[708] + Check_Bit[709] + Check_Bit[710] + Check_Bit[711] + Check_Bit[712] + Check_Bit[713] + Check_Bit[714] + Check_Bit[715] + Check_Bit[716] + Check_Bit[717] + Check_Bit[718] + Check_Bit[719] + Check_Bit[720] + Check_Bit[721] + Check_Bit[722] + Check_Bit[723] + Check_Bit[724] + Check_Bit[725] + Check_Bit[726] + Check_Bit[727] + Check_Bit[728] + Check_Bit[729] + Check_Bit[730] + Check_Bit[731] + Check_Bit[732] + Check_Bit[733] + Check_Bit[734] + Check_Bit[735] + Check_Bit[736] + Check_Bit[737] + Check_Bit[738] + Check_Bit[739] + Check_Bit[740] + Check_Bit[741] + Check_Bit[742] + Check_Bit[743] + Check_Bit[744] + Check_Bit[745] + Check_Bit[746] + Check_Bit[747] + Check_Bit[748] + Check_Bit[749] + Check_Bit[750] + Check_Bit[751] + Check_Bit[752] + Check_Bit[753] + Check_Bit[754] + Check_Bit[755] + Check_Bit[756] + Check_Bit[757] + Check_Bit[758] + Check_Bit[759] + Check_Bit[760] + Check_Bit[761] + Check_Bit[762] + Check_Bit[763] + Check_Bit[764] + Check_Bit[765] + Check_Bit[766] + Check_Bit[767] + Check_Bit[768] + Check_Bit[769] + Check_Bit[770] + Check_Bit[771] + Check_Bit[772] + Check_Bit[773] + Check_Bit[774] + Check_Bit[775] + Check_Bit[776] + Check_Bit[777] + Check_Bit[778] + Check_Bit[779] + Check_Bit[780] + Check_Bit[781] + Check_Bit[782] + Check_Bit[783] + Check_Bit[784] + Check_Bit[785] + Check_Bit[786] + Check_Bit[787] + Check_Bit[788] + Check_Bit[789] + Check_Bit[790] + Check_Bit[791] + Check_Bit[792] + Check_Bit[793] + Check_Bit[794] + Check_Bit[795] + Check_Bit[796] + Check_Bit[797] + Check_Bit[798] + Check_Bit[799] + Check_Bit[800] + Check_Bit[801] + Check_Bit[802] + Check_Bit[803] + Check_Bit[804] + Check_Bit[805] + Check_Bit[806] + Check_Bit[807] + Check_Bit[808] + Check_Bit[809] + Check_Bit[810] + Check_Bit[811] + Check_Bit[812] + Check_Bit[813] + Check_Bit[814] + Check_Bit[815] + Check_Bit[816] + Check_Bit[817] + Check_Bit[818] + Check_Bit[819] + Check_Bit[820] + Check_Bit[821] + Check_Bit[822] + Check_Bit[823] + Check_Bit[824] + Check_Bit[825] + Check_Bit[826] + Check_Bit[827] + Check_Bit[828] + Check_Bit[829] + Check_Bit[830] + Check_Bit[831] + Check_Bit[832] + Check_Bit[833] + Check_Bit[834] + Check_Bit[835] + Check_Bit[836] + Check_Bit[837] + Check_Bit[838] + Check_Bit[839] + Check_Bit[840] + Check_Bit[841] + Check_Bit[842] + Check_Bit[843] + Check_Bit[844] + Check_Bit[845] + Check_Bit[846] + Check_Bit[847] + Check_Bit[848] + Check_Bit[849] + Check_Bit[850] + Check_Bit[851] + Check_Bit[852] + Check_Bit[853] + Check_Bit[854] + Check_Bit[855] + Check_Bit[856] + Check_Bit[857] + Check_Bit[858] + Check_Bit[859] + Check_Bit[860] + Check_Bit[861] + Check_Bit[862] + Check_Bit[863] + Check_Bit[864] + Check_Bit[865] + Check_Bit[866] + Check_Bit[867] + Check_Bit[868] + Check_Bit[869] + Check_Bit[870] + Check_Bit[871] + Check_Bit[872] + Check_Bit[873] + Check_Bit[874] + Check_Bit[875] + Check_Bit[876] + Check_Bit[877] + Check_Bit[878] + Check_Bit[879] + Check_Bit[880] + Check_Bit[881] + Check_Bit[882] + Check_Bit[883] + Check_Bit[884] + Check_Bit[885] + Check_Bit[886] + Check_Bit[887] + Check_Bit[888] + Check_Bit[889] + Check_Bit[890] + Check_Bit[891] + Check_Bit[892] + Check_Bit[893] + Check_Bit[894] + Check_Bit[895] + Check_Bit[896] + Check_Bit[897] + Check_Bit[898] + Check_Bit[899] + Check_Bit[900] + Check_Bit[901] + Check_Bit[902] + Check_Bit[903] + Check_Bit[904] + Check_Bit[905] + Check_Bit[906] + Check_Bit[907] + Check_Bit[908] + Check_Bit[909] + Check_Bit[910] + Check_Bit[911] + Check_Bit[912] + Check_Bit[913] + Check_Bit[914] + Check_Bit[915] + Check_Bit[916] + Check_Bit[917] + Check_Bit[918] + Check_Bit[919] + Check_Bit[920] + Check_Bit[921] + Check_Bit[922] + Check_Bit[923] + Check_Bit[924] + Check_Bit[925] + Check_Bit[926] + Check_Bit[927] + Check_Bit[928] + Check_Bit[929] + Check_Bit[930] + Check_Bit[931] + Check_Bit[932] + Check_Bit[933] + Check_Bit[934] + Check_Bit[935] + Check_Bit[936] + Check_Bit[937] + Check_Bit[938] + Check_Bit[939] + Check_Bit[940] + Check_Bit[941] + Check_Bit[942] + Check_Bit[943] + Check_Bit[944] + Check_Bit[945] + Check_Bit[946] + Check_Bit[947] + Check_Bit[948] + Check_Bit[949] + Check_Bit[950] + Check_Bit[951] + Check_Bit[952] + Check_Bit[953] + Check_Bit[954] + Check_Bit[955] + Check_Bit[956] + Check_Bit[957] + Check_Bit[958] + Check_Bit[959] + Check_Bit[960] + Check_Bit[961] + Check_Bit[962] + Check_Bit[963] + Check_Bit[964] + Check_Bit[965] + Check_Bit[966] + Check_Bit[967] + Check_Bit[968] + Check_Bit[969] + Check_Bit[970] + Check_Bit[971] + Check_Bit[972] + Check_Bit[973] + Check_Bit[974] + Check_Bit[975] + Check_Bit[976] + Check_Bit[977] + Check_Bit[978] + Check_Bit[979] + Check_Bit[980] + Check_Bit[981] + Check_Bit[982] + Check_Bit[983] + Check_Bit[984] + Check_Bit[985] + Check_Bit[986] + Check_Bit[987] + Check_Bit[988] + Check_Bit[989] + Check_Bit[990] + Check_Bit[991] + Check_Bit[992] + Check_Bit[993] + Check_Bit[994] + Check_Bit[995] + Check_Bit[996] + Check_Bit[997] + Check_Bit[998] + Check_Bit[999] + Check_Bit[1000] + Check_Bit[1001] + Check_Bit[1002] + Check_Bit[1003] + Check_Bit[1004] + Check_Bit[1005] + Check_Bit[1006] + Check_Bit[1007] + Check_Bit[1008] + Check_Bit[1009] + Check_Bit[1010] + Check_Bit[1011] + Check_Bit[1012] + Check_Bit[1013] + Check_Bit[1014] + Check_Bit[1015] + Check_Bit[1016] + Check_Bit[1017] + Check_Bit[1018] + Check_Bit[1019] + Check_Bit[1020] + Check_Bit[1021] + Check_Bit[1022] + Check_Bit[1023] + Check_Bit[1024] + Check_Bit[1025] + Check_Bit[1026] + Check_Bit[1027] + Check_Bit[1028] + Check_Bit[1029] + Check_Bit[1030] + Check_Bit[1031] + Check_Bit[1032] + Check_Bit[1033] + Check_Bit[1034] + Check_Bit[1035] + Check_Bit[1036] + Check_Bit[1037] + Check_Bit[1038] + Check_Bit[1039] + Check_Bit[1040] + Check_Bit[1041] + Check_Bit[1042] + Check_Bit[1043] + Check_Bit[1044] + Check_Bit[1045] + Check_Bit[1046] + Check_Bit[1047] + Check_Bit[1048] + Check_Bit[1049] + Check_Bit[1050] + Check_Bit[1051] + Check_Bit[1052] + Check_Bit[1053] + Check_Bit[1054] + Check_Bit[1055] + Check_Bit[1056] + Check_Bit[1057] + Check_Bit[1058] + Check_Bit[1059] + Check_Bit[1060] + Check_Bit[1061] + Check_Bit[1062] + Check_Bit[1063] + Check_Bit[1064] + Check_Bit[1065] + Check_Bit[1066] + Check_Bit[1067] + Check_Bit[1068] + Check_Bit[1069] + Check_Bit[1070] + Check_Bit[1071] + Check_Bit[1072] + Check_Bit[1073] + Check_Bit[1074] + Check_Bit[1075] + Check_Bit[1076] + Check_Bit[1077] + Check_Bit[1078] + Check_Bit[1079] + Check_Bit[1080] + Check_Bit[1081] + Check_Bit[1082] + Check_Bit[1083] + Check_Bit[1084] + Check_Bit[1085] + Check_Bit[1086] + Check_Bit[1087] + Check_Bit[1088] + Check_Bit[1089] + Check_Bit[1090] + Check_Bit[1091] + Check_Bit[1092] + Check_Bit[1093] + Check_Bit[1094] + Check_Bit[1095] + Check_Bit[1096] + Check_Bit[1097] + Check_Bit[1098] + Check_Bit[1099] + Check_Bit[1100] + Check_Bit[1101] + Check_Bit[1102] + Check_Bit[1103] + Check_Bit[1104] + Check_Bit[1105] + Check_Bit[1106] + Check_Bit[1107] + Check_Bit[1108] + Check_Bit[1109] + Check_Bit[1110] + Check_Bit[1111] + Check_Bit[1112] + Check_Bit[1113] + Check_Bit[1114] + Check_Bit[1115] + Check_Bit[1116] + Check_Bit[1117] + Check_Bit[1118] + Check_Bit[1119] + Check_Bit[1120] + Check_Bit[1121] + Check_Bit[1122] + Check_Bit[1123] + Check_Bit[1124] + Check_Bit[1125] + Check_Bit[1126] + Check_Bit[1127] + Check_Bit[1128] + Check_Bit[1129] + Check_Bit[1130] + Check_Bit[1131] + Check_Bit[1132] + Check_Bit[1133] + Check_Bit[1134] + Check_Bit[1135] + Check_Bit[1136] + Check_Bit[1137] + Check_Bit[1138] + Check_Bit[1139] + Check_Bit[1140] + Check_Bit[1141] + Check_Bit[1142] + Check_Bit[1143] + Check_Bit[1144] + Check_Bit[1145] + Check_Bit[1146] + Check_Bit[1147] + Check_Bit[1148] + Check_Bit[1149] + Check_Bit[1150] + Check_Bit[1151] + Check_Bit[1152] + Check_Bit[1153] + Check_Bit[1154] + Check_Bit[1155] + Check_Bit[1156] + Check_Bit[1157] + Check_Bit[1158] + Check_Bit[1159] + Check_Bit[1160] + Check_Bit[1161] + Check_Bit[1162] + Check_Bit[1163] + Check_Bit[1164] + Check_Bit[1165] + Check_Bit[1166] + Check_Bit[1167] + Check_Bit[1168] + Check_Bit[1169] + Check_Bit[1170] + Check_Bit[1171] + Check_Bit[1172] + Check_Bit[1173] + Check_Bit[1174] + Check_Bit[1175] + Check_Bit[1176] + Check_Bit[1177] + Check_Bit[1178] + Check_Bit[1179] + Check_Bit[1180] + Check_Bit[1181] + Check_Bit[1182] + Check_Bit[1183] + Check_Bit[1184] + Check_Bit[1185] + Check_Bit[1186] + Check_Bit[1187] + Check_Bit[1188] + Check_Bit[1189] + Check_Bit[1190] + Check_Bit[1191] + Check_Bit[1192] + Check_Bit[1193] + Check_Bit[1194] + Check_Bit[1195] + Check_Bit[1196] + Check_Bit[1197] + Check_Bit[1198] + Check_Bit[1199] + Check_Bit[1200] + Check_Bit[1201] + Check_Bit[1202] + Check_Bit[1203] + Check_Bit[1204] + Check_Bit[1205] + Check_Bit[1206] + Check_Bit[1207] + Check_Bit[1208] + Check_Bit[1209] + Check_Bit[1210] + Check_Bit[1211] + Check_Bit[1212] + Check_Bit[1213] + Check_Bit[1214] + Check_Bit[1215] + Check_Bit[1216] + Check_Bit[1217] + Check_Bit[1218] + Check_Bit[1219] + Check_Bit[1220] + Check_Bit[1221] + Check_Bit[1222] + Check_Bit[1223] + Check_Bit[1224] + Check_Bit[1225] + Check_Bit[1226] + Check_Bit[1227] + Check_Bit[1228] + Check_Bit[1229] + Check_Bit[1230] + Check_Bit[1231] + Check_Bit[1232] + Check_Bit[1233] + Check_Bit[1234] + Check_Bit[1235] + Check_Bit[1236] + Check_Bit[1237] + Check_Bit[1238] + Check_Bit[1239] + Check_Bit[1240] + Check_Bit[1241] + Check_Bit[1242] + Check_Bit[1243] + Check_Bit[1244] + Check_Bit[1245] + Check_Bit[1246] + Check_Bit[1247] + Check_Bit[1248] + Check_Bit[1249] + Check_Bit[1250] + Check_Bit[1251] + Check_Bit[1252] + Check_Bit[1253] + Check_Bit[1254] + Check_Bit[1255] + Check_Bit[1256] + Check_Bit[1257] + Check_Bit[1258] + Check_Bit[1259] + Check_Bit[1260] + Check_Bit[1261] + Check_Bit[1262] + Check_Bit[1263] + Check_Bit[1264] + Check_Bit[1265] + Check_Bit[1266] + Check_Bit[1267] + Check_Bit[1268] + Check_Bit[1269] + Check_Bit[1270] + Check_Bit[1271] + Check_Bit[1272] + Check_Bit[1273] + Check_Bit[1274] + Check_Bit[1275] + Check_Bit[1276] + Check_Bit[1277] + Check_Bit[1278] + Check_Bit[1279] + Check_Bit[1280] + Check_Bit[1281] + Check_Bit[1282] + Check_Bit[1283] + Check_Bit[1284] + Check_Bit[1285] + Check_Bit[1286] + Check_Bit[1287] + Check_Bit[1288] + Check_Bit[1289] + Check_Bit[1290] + Check_Bit[1291] + Check_Bit[1292] + Check_Bit[1293] + Check_Bit[1294] + Check_Bit[1295] + Check_Bit[1296] + Check_Bit[1297] + Check_Bit[1298] + Check_Bit[1299] + Check_Bit[1300] + Check_Bit[1301] + Check_Bit[1302] + Check_Bit[1303] + Check_Bit[1304] + Check_Bit[1305] + Check_Bit[1306] + Check_Bit[1307] + Check_Bit[1308] + Check_Bit[1309] + Check_Bit[1310] + Check_Bit[1311] + Check_Bit[1312] + Check_Bit[1313] + Check_Bit[1314] + Check_Bit[1315] + Check_Bit[1316] + Check_Bit[1317] + Check_Bit[1318] + Check_Bit[1319] + Check_Bit[1320] + Check_Bit[1321] + Check_Bit[1322] + Check_Bit[1323] + Check_Bit[1324] + Check_Bit[1325] + Check_Bit[1326] + Check_Bit[1327] + Check_Bit[1328] + Check_Bit[1329] + Check_Bit[1330] + Check_Bit[1331] + Check_Bit[1332] + Check_Bit[1333] + Check_Bit[1334] + Check_Bit[1335] + Check_Bit[1336] + Check_Bit[1337] + Check_Bit[1338] + Check_Bit[1339] + Check_Bit[1340] + Check_Bit[1341] + Check_Bit[1342] + Check_Bit[1343] + Check_Bit[1344] + Check_Bit[1345] + Check_Bit[1346] + Check_Bit[1347] + Check_Bit[1348] + Check_Bit[1349] + Check_Bit[1350] + Check_Bit[1351] + Check_Bit[1352] + Check_Bit[1353] + Check_Bit[1354] + Check_Bit[1355] + Check_Bit[1356] + Check_Bit[1357] + Check_Bit[1358] + Check_Bit[1359] + Check_Bit[1360] + Check_Bit[1361] + Check_Bit[1362] + Check_Bit[1363] + Check_Bit[1364] + Check_Bit[1365] + Check_Bit[1366] + Check_Bit[1367] + Check_Bit[1368] + Check_Bit[1369] + Check_Bit[1370] + Check_Bit[1371] + Check_Bit[1372] + Check_Bit[1373] + Check_Bit[1374] + Check_Bit[1375] + Check_Bit[1376] + Check_Bit[1377] + Check_Bit[1378] + Check_Bit[1379] + Check_Bit[1380] + Check_Bit[1381] + Check_Bit[1382] + Check_Bit[1383] + Check_Bit[1384] + Check_Bit[1385] + Check_Bit[1386] + Check_Bit[1387] + Check_Bit[1388] + Check_Bit[1389] + Check_Bit[1390] + Check_Bit[1391] + Check_Bit[1392] + Check_Bit[1393] + Check_Bit[1394] + Check_Bit[1395] + Check_Bit[1396] + Check_Bit[1397] + Check_Bit[1398] + Check_Bit[1399] + Check_Bit[1400] + Check_Bit[1401] + Check_Bit[1402] + Check_Bit[1403] + Check_Bit[1404] + Check_Bit[1405] + Check_Bit[1406] + Check_Bit[1407] + Check_Bit[1408] + Check_Bit[1409] + Check_Bit[1410] + Check_Bit[1411] + Check_Bit[1412] + Check_Bit[1413] + Check_Bit[1414] + Check_Bit[1415] + Check_Bit[1416] + Check_Bit[1417] + Check_Bit[1418] + Check_Bit[1419] + Check_Bit[1420] + Check_Bit[1421] + Check_Bit[1422] + Check_Bit[1423] + Check_Bit[1424] + Check_Bit[1425] + Check_Bit[1426] + Check_Bit[1427] + Check_Bit[1428] + Check_Bit[1429] + Check_Bit[1430] + Check_Bit[1431] + Check_Bit[1432] + Check_Bit[1433] + Check_Bit[1434] + Check_Bit[1435] + Check_Bit[1436] + Check_Bit[1437] + Check_Bit[1438] + Check_Bit[1440 - 1];
Decoder Decoder1 (
.clk (clk),
.rst (rst),
.in_valid (in_valid),
.in_index (in_index),
.data_in (L [(in_index+4)*10-1-:10*4]),
.out_valid(out_valid),
//.Bit (Bit),
.out_index (out_index));
endmodule
