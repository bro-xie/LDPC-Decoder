module Decoder #(
	parameter code_length = 1440,
	parameter quan_width = 15
)
(
	input wire clk,
	input wire rst,
	input wire in_valid,
	input wire [15:0] in_index,
	input wire [4 * quan_width - 1: 0] data_in,
	output reg out_valid,
	output reg [15:0] out_index,
	output reg [4 - 1: 0] data_out,
	output wire [code_length - 1:0] Bit
);

reg [code_length * quan_width - 1 : 0] L;
// wire [code_length - 1:0] Bit;
reg [7:0] cnt;
reg [4:0] iter;
reg Check_1, Check_2, Check_3, Check_4, Check_5, Check_6, Check_7, Check_8, Check_9, Check_10, Check_11, Check_12, Check_13, Check_14, Check_15, Check_16, Check_17, Check_18, Check_19, Check_20, Check_21, Check_22, Check_23, Check_24, Check_25, Check_26, Check_27, Check_28, Check_29, Check_30, Check_31, Check_32, Check_33, Check_34, Check_35, Check_36, Check_37, Check_38, Check_39, Check_40, Check_41, Check_42, Check_43, Check_44, Check_45, Check_46, Check_47, Check_48, Check_49, Check_50, Check_51, Check_52, Check_53, Check_54, Check_55, Check_56, Check_57, Check_58, Check_59, Check_60, Check_61, Check_62, Check_63, Check_64, Check_65, Check_66, Check_67, Check_68, Check_69, Check_70, Check_71, Check_72, Check_73, Check_74, Check_75, Check_76, Check_77, Check_78, Check_79, Check_80, Check_81, Check_82, Check_83, Check_84, Check_85, Check_86, Check_87, Check_88, Check_89, Check_90, Check_91, Check_92, Check_93, Check_94, Check_95, Check_96, Check_97, Check_98, Check_99, Check_100, Check_101, Check_102, Check_103, Check_104, Check_105, Check_106, Check_107, Check_108, Check_109, Check_110, Check_111, Check_112, Check_113, Check_114, Check_115, Check_116, Check_117, Check_118, Check_119, Check_120, Check_121, Check_122, Check_123, Check_124, Check_125, Check_126, Check_127, Check_128, Check_129, Check_130, Check_131, Check_132, Check_133, Check_134, Check_135, Check_136, Check_137, Check_138, Check_139, Check_140, Check_141, Check_142, Check_143, Check_144, Check_145, Check_146, Check_147, Check_148, Check_149, Check_150, Check_151, Check_152, Check_153, Check_154, Check_155, Check_156, Check_157, Check_158, Check_159, Check_160, Check_161, Check_162, Check_163, Check_164, Check_165, Check_166, Check_167, Check_168, Check_169, Check_170, Check_171, Check_172, Check_173, Check_174, Check_175, Check_176, Check_177, Check_178, Check_179, Check_180, Check_181, Check_182, Check_183, Check_184, Check_185, Check_186, Check_187, Check_188, Check_189, Check_190, Check_191, Check_192, Check_193, Check_194, Check_195, Check_196, Check_197, Check_198, Check_199, Check_200, Check_201, Check_202, Check_203, Check_204, Check_205, Check_206, Check_207, Check_208, Check_209, Check_210, Check_211, Check_212, Check_213, Check_214, Check_215, Check_216, Check_217, Check_218, Check_219, Check_220, Check_221, Check_222, Check_223, Check_224, Check_225, Check_226, Check_227, Check_228, Check_229, Check_230, Check_231, Check_232, Check_233, Check_234, Check_235, Check_236, Check_237, Check_238, Check_239, Check_240, Check_241, Check_242, Check_243, Check_244, Check_245, Check_246, Check_247, Check_248, Check_249, Check_250, Check_251, Check_252, Check_253, Check_254, Check_255, Check_256, Check_257, Check_258, Check_259, Check_260, Check_261, Check_262, Check_263, Check_264, Check_265, Check_266, Check_267, Check_268, Check_269, Check_270, Check_271, Check_272, Check_273, Check_274, Check_275, Check_276, Check_277, Check_278, Check_279, Check_280, Check_281, Check_282, Check_283, Check_284, Check_285, Check_286, Check_287, Check_288, Check_Sum;
wire [quan_width - 1:0] C2V_1_5, C2V_1_89, C2V_1_109, C2V_1_170, C2V_1_232, C2V_1_275, C2V_1_375, C2V_1_429, C2V_1_526, C2V_1_762, C2V_1_810, C2V_1_858, C2V_1_899, C2V_1_940, C2V_1_974, C2V_1_1013, C2V_1_1087, C2V_1_1146, C2V_1_1153, C2V_2_14, C2V_2_63, C2V_2_119, C2V_2_167, C2V_2_196, C2V_2_265, C2V_2_316, C2V_2_423, C2V_2_512, C2V_2_672, C2V_2_685, C2V_2_853, C2V_2_895, C2V_2_958, C2V_2_989, C2V_2_1021, C2V_2_1088, C2V_2_1119, C2V_2_1153, C2V_2_1154, C2V_3_9, C2V_3_84, C2V_3_101, C2V_3_183, C2V_3_201, C2V_3_268, C2V_3_365, C2V_3_420, C2V_3_531, C2V_3_588, C2V_3_664, C2V_3_768, C2V_3_899, C2V_3_943, C2V_3_968, C2V_3_1028, C2V_3_1058, C2V_3_1151, C2V_3_1154, C2V_3_1155, C2V_4_28, C2V_4_87, C2V_4_126, C2V_4_182, C2V_4_199, C2V_4_253, C2V_4_477, C2V_4_517, C2V_4_553, C2V_4_615, C2V_4_640, C2V_4_686, C2V_4_903, C2V_4_927, C2V_4_963, C2V_4_1041, C2V_4_1068, C2V_4_1132, C2V_4_1155, C2V_4_1156, C2V_5_47, C2V_5_57, C2V_5_140, C2V_5_163, C2V_5_227, C2V_5_245, C2V_5_294, C2V_5_361, C2V_5_440, C2V_5_674, C2V_5_738, C2V_5_792, C2V_5_870, C2V_5_918, C2V_5_961, C2V_5_1013, C2V_5_1062, C2V_5_1110, C2V_5_1156, C2V_5_1157, C2V_6_30, C2V_6_54, C2V_6_142, C2V_6_162, C2V_6_196, C2V_6_275, C2V_6_328, C2V_6_480, C2V_6_529, C2V_6_610, C2V_6_814, C2V_6_842, C2V_6_875, C2V_6_937, C2V_6_972, C2V_6_1039, C2V_6_1103, C2V_6_1105, C2V_6_1157, C2V_6_1158, C2V_7_6, C2V_7_90, C2V_7_110, C2V_7_171, C2V_7_233, C2V_7_276, C2V_7_376, C2V_7_430, C2V_7_527, C2V_7_763, C2V_7_811, C2V_7_859, C2V_7_900, C2V_7_941, C2V_7_975, C2V_7_1014, C2V_7_1088, C2V_7_1147, C2V_7_1158, C2V_7_1159, C2V_8_15, C2V_8_64, C2V_8_120, C2V_8_168, C2V_8_197, C2V_8_266, C2V_8_317, C2V_8_424, C2V_8_513, C2V_8_625, C2V_8_686, C2V_8_854, C2V_8_896, C2V_8_959, C2V_8_990, C2V_8_1022, C2V_8_1089, C2V_8_1120, C2V_8_1159, C2V_8_1160, C2V_9_10, C2V_9_85, C2V_9_102, C2V_9_184, C2V_9_202, C2V_9_269, C2V_9_366, C2V_9_421, C2V_9_532, C2V_9_589, C2V_9_665, C2V_9_721, C2V_9_900, C2V_9_944, C2V_9_969, C2V_9_1029, C2V_9_1059, C2V_9_1152, C2V_9_1160, C2V_9_1161, C2V_10_29, C2V_10_88, C2V_10_127, C2V_10_183, C2V_10_200, C2V_10_254, C2V_10_478, C2V_10_518, C2V_10_554, C2V_10_616, C2V_10_641, C2V_10_687, C2V_10_904, C2V_10_928, C2V_10_964, C2V_10_1042, C2V_10_1069, C2V_10_1133, C2V_10_1161, C2V_10_1162, C2V_11_48, C2V_11_58, C2V_11_141, C2V_11_164, C2V_11_228, C2V_11_246, C2V_11_295, C2V_11_362, C2V_11_441, C2V_11_675, C2V_11_739, C2V_11_793, C2V_11_871, C2V_11_919, C2V_11_962, C2V_11_1014, C2V_11_1063, C2V_11_1111, C2V_11_1162, C2V_11_1163, C2V_12_31, C2V_12_55, C2V_12_143, C2V_12_163, C2V_12_197, C2V_12_276, C2V_12_329, C2V_12_433, C2V_12_530, C2V_12_611, C2V_12_815, C2V_12_843, C2V_12_876, C2V_12_938, C2V_12_973, C2V_12_1040, C2V_12_1104, C2V_12_1106, C2V_12_1163, C2V_12_1164, C2V_13_7, C2V_13_91, C2V_13_111, C2V_13_172, C2V_13_234, C2V_13_277, C2V_13_377, C2V_13_431, C2V_13_528, C2V_13_764, C2V_13_812, C2V_13_860, C2V_13_901, C2V_13_942, C2V_13_976, C2V_13_1015, C2V_13_1089, C2V_13_1148, C2V_13_1164, C2V_13_1165, C2V_14_16, C2V_14_65, C2V_14_121, C2V_14_169, C2V_14_198, C2V_14_267, C2V_14_318, C2V_14_425, C2V_14_514, C2V_14_626, C2V_14_687, C2V_14_855, C2V_14_897, C2V_14_960, C2V_14_991, C2V_14_1023, C2V_14_1090, C2V_14_1121, C2V_14_1165, C2V_14_1166, C2V_15_11, C2V_15_86, C2V_15_103, C2V_15_185, C2V_15_203, C2V_15_270, C2V_15_367, C2V_15_422, C2V_15_533, C2V_15_590, C2V_15_666, C2V_15_722, C2V_15_901, C2V_15_945, C2V_15_970, C2V_15_1030, C2V_15_1060, C2V_15_1105, C2V_15_1166, C2V_15_1167, C2V_16_30, C2V_16_89, C2V_16_128, C2V_16_184, C2V_16_201, C2V_16_255, C2V_16_479, C2V_16_519, C2V_16_555, C2V_16_617, C2V_16_642, C2V_16_688, C2V_16_905, C2V_16_929, C2V_16_965, C2V_16_1043, C2V_16_1070, C2V_16_1134, C2V_16_1167, C2V_16_1168, C2V_17_1, C2V_17_59, C2V_17_142, C2V_17_165, C2V_17_229, C2V_17_247, C2V_17_296, C2V_17_363, C2V_17_442, C2V_17_676, C2V_17_740, C2V_17_794, C2V_17_872, C2V_17_920, C2V_17_963, C2V_17_1015, C2V_17_1064, C2V_17_1112, C2V_17_1168, C2V_17_1169, C2V_18_32, C2V_18_56, C2V_18_144, C2V_18_164, C2V_18_198, C2V_18_277, C2V_18_330, C2V_18_434, C2V_18_531, C2V_18_612, C2V_18_816, C2V_18_844, C2V_18_877, C2V_18_939, C2V_18_974, C2V_18_1041, C2V_18_1057, C2V_18_1107, C2V_18_1169, C2V_18_1170, C2V_19_8, C2V_19_92, C2V_19_112, C2V_19_173, C2V_19_235, C2V_19_278, C2V_19_378, C2V_19_432, C2V_19_481, C2V_19_765, C2V_19_813, C2V_19_861, C2V_19_902, C2V_19_943, C2V_19_977, C2V_19_1016, C2V_19_1090, C2V_19_1149, C2V_19_1170, C2V_19_1171, C2V_20_17, C2V_20_66, C2V_20_122, C2V_20_170, C2V_20_199, C2V_20_268, C2V_20_319, C2V_20_426, C2V_20_515, C2V_20_627, C2V_20_688, C2V_20_856, C2V_20_898, C2V_20_913, C2V_20_992, C2V_20_1024, C2V_20_1091, C2V_20_1122, C2V_20_1171, C2V_20_1172, C2V_21_12, C2V_21_87, C2V_21_104, C2V_21_186, C2V_21_204, C2V_21_271, C2V_21_368, C2V_21_423, C2V_21_534, C2V_21_591, C2V_21_667, C2V_21_723, C2V_21_902, C2V_21_946, C2V_21_971, C2V_21_1031, C2V_21_1061, C2V_21_1106, C2V_21_1172, C2V_21_1173, C2V_22_31, C2V_22_90, C2V_22_129, C2V_22_185, C2V_22_202, C2V_22_256, C2V_22_480, C2V_22_520, C2V_22_556, C2V_22_618, C2V_22_643, C2V_22_689, C2V_22_906, C2V_22_930, C2V_22_966, C2V_22_1044, C2V_22_1071, C2V_22_1135, C2V_22_1173, C2V_22_1174, C2V_23_2, C2V_23_60, C2V_23_143, C2V_23_166, C2V_23_230, C2V_23_248, C2V_23_297, C2V_23_364, C2V_23_443, C2V_23_677, C2V_23_741, C2V_23_795, C2V_23_873, C2V_23_921, C2V_23_964, C2V_23_1016, C2V_23_1065, C2V_23_1113, C2V_23_1174, C2V_23_1175, C2V_24_33, C2V_24_57, C2V_24_97, C2V_24_165, C2V_24_199, C2V_24_278, C2V_24_331, C2V_24_435, C2V_24_532, C2V_24_613, C2V_24_769, C2V_24_845, C2V_24_878, C2V_24_940, C2V_24_975, C2V_24_1042, C2V_24_1058, C2V_24_1108, C2V_24_1175, C2V_24_1176, C2V_25_9, C2V_25_93, C2V_25_113, C2V_25_174, C2V_25_236, C2V_25_279, C2V_25_379, C2V_25_385, C2V_25_482, C2V_25_766, C2V_25_814, C2V_25_862, C2V_25_903, C2V_25_944, C2V_25_978, C2V_25_1017, C2V_25_1091, C2V_25_1150, C2V_25_1176, C2V_25_1177, C2V_26_18, C2V_26_67, C2V_26_123, C2V_26_171, C2V_26_200, C2V_26_269, C2V_26_320, C2V_26_427, C2V_26_516, C2V_26_628, C2V_26_689, C2V_26_857, C2V_26_899, C2V_26_914, C2V_26_993, C2V_26_1025, C2V_26_1092, C2V_26_1123, C2V_26_1177, C2V_26_1178, C2V_27_13, C2V_27_88, C2V_27_105, C2V_27_187, C2V_27_205, C2V_27_272, C2V_27_369, C2V_27_424, C2V_27_535, C2V_27_592, C2V_27_668, C2V_27_724, C2V_27_903, C2V_27_947, C2V_27_972, C2V_27_1032, C2V_27_1062, C2V_27_1107, C2V_27_1178, C2V_27_1179, C2V_28_32, C2V_28_91, C2V_28_130, C2V_28_186, C2V_28_203, C2V_28_257, C2V_28_433, C2V_28_521, C2V_28_557, C2V_28_619, C2V_28_644, C2V_28_690, C2V_28_907, C2V_28_931, C2V_28_967, C2V_28_1045, C2V_28_1072, C2V_28_1136, C2V_28_1179, C2V_28_1180, C2V_29_3, C2V_29_61, C2V_29_144, C2V_29_167, C2V_29_231, C2V_29_249, C2V_29_298, C2V_29_365, C2V_29_444, C2V_29_678, C2V_29_742, C2V_29_796, C2V_29_874, C2V_29_922, C2V_29_965, C2V_29_1017, C2V_29_1066, C2V_29_1114, C2V_29_1180, C2V_29_1181, C2V_30_34, C2V_30_58, C2V_30_98, C2V_30_166, C2V_30_200, C2V_30_279, C2V_30_332, C2V_30_436, C2V_30_533, C2V_30_614, C2V_30_770, C2V_30_846, C2V_30_879, C2V_30_941, C2V_30_976, C2V_30_1043, C2V_30_1059, C2V_30_1109, C2V_30_1181, C2V_30_1182, C2V_31_10, C2V_31_94, C2V_31_114, C2V_31_175, C2V_31_237, C2V_31_280, C2V_31_380, C2V_31_386, C2V_31_483, C2V_31_767, C2V_31_815, C2V_31_863, C2V_31_904, C2V_31_945, C2V_31_979, C2V_31_1018, C2V_31_1092, C2V_31_1151, C2V_31_1182, C2V_31_1183, C2V_32_19, C2V_32_68, C2V_32_124, C2V_32_172, C2V_32_201, C2V_32_270, C2V_32_321, C2V_32_428, C2V_32_517, C2V_32_629, C2V_32_690, C2V_32_858, C2V_32_900, C2V_32_915, C2V_32_994, C2V_32_1026, C2V_32_1093, C2V_32_1124, C2V_32_1183, C2V_32_1184, C2V_33_14, C2V_33_89, C2V_33_106, C2V_33_188, C2V_33_206, C2V_33_273, C2V_33_370, C2V_33_425, C2V_33_536, C2V_33_593, C2V_33_669, C2V_33_725, C2V_33_904, C2V_33_948, C2V_33_973, C2V_33_1033, C2V_33_1063, C2V_33_1108, C2V_33_1184, C2V_33_1185, C2V_34_33, C2V_34_92, C2V_34_131, C2V_34_187, C2V_34_204, C2V_34_258, C2V_34_434, C2V_34_522, C2V_34_558, C2V_34_620, C2V_34_645, C2V_34_691, C2V_34_908, C2V_34_932, C2V_34_968, C2V_34_1046, C2V_34_1073, C2V_34_1137, C2V_34_1185, C2V_34_1186, C2V_35_4, C2V_35_62, C2V_35_97, C2V_35_168, C2V_35_232, C2V_35_250, C2V_35_299, C2V_35_366, C2V_35_445, C2V_35_679, C2V_35_743, C2V_35_797, C2V_35_875, C2V_35_923, C2V_35_966, C2V_35_1018, C2V_35_1067, C2V_35_1115, C2V_35_1186, C2V_35_1187, C2V_36_35, C2V_36_59, C2V_36_99, C2V_36_167, C2V_36_201, C2V_36_280, C2V_36_333, C2V_36_437, C2V_36_534, C2V_36_615, C2V_36_771, C2V_36_847, C2V_36_880, C2V_36_942, C2V_36_977, C2V_36_1044, C2V_36_1060, C2V_36_1110, C2V_36_1187, C2V_36_1188, C2V_37_11, C2V_37_95, C2V_37_115, C2V_37_176, C2V_37_238, C2V_37_281, C2V_37_381, C2V_37_387, C2V_37_484, C2V_37_768, C2V_37_816, C2V_37_864, C2V_37_905, C2V_37_946, C2V_37_980, C2V_37_1019, C2V_37_1093, C2V_37_1152, C2V_37_1188, C2V_37_1189, C2V_38_20, C2V_38_69, C2V_38_125, C2V_38_173, C2V_38_202, C2V_38_271, C2V_38_322, C2V_38_429, C2V_38_518, C2V_38_630, C2V_38_691, C2V_38_859, C2V_38_901, C2V_38_916, C2V_38_995, C2V_38_1027, C2V_38_1094, C2V_38_1125, C2V_38_1189, C2V_38_1190, C2V_39_15, C2V_39_90, C2V_39_107, C2V_39_189, C2V_39_207, C2V_39_274, C2V_39_371, C2V_39_426, C2V_39_537, C2V_39_594, C2V_39_670, C2V_39_726, C2V_39_905, C2V_39_949, C2V_39_974, C2V_39_1034, C2V_39_1064, C2V_39_1109, C2V_39_1190, C2V_39_1191, C2V_40_34, C2V_40_93, C2V_40_132, C2V_40_188, C2V_40_205, C2V_40_259, C2V_40_435, C2V_40_523, C2V_40_559, C2V_40_621, C2V_40_646, C2V_40_692, C2V_40_909, C2V_40_933, C2V_40_969, C2V_40_1047, C2V_40_1074, C2V_40_1138, C2V_40_1191, C2V_40_1192, C2V_41_5, C2V_41_63, C2V_41_98, C2V_41_169, C2V_41_233, C2V_41_251, C2V_41_300, C2V_41_367, C2V_41_446, C2V_41_680, C2V_41_744, C2V_41_798, C2V_41_876, C2V_41_924, C2V_41_967, C2V_41_1019, C2V_41_1068, C2V_41_1116, C2V_41_1192, C2V_41_1193, C2V_42_36, C2V_42_60, C2V_42_100, C2V_42_168, C2V_42_202, C2V_42_281, C2V_42_334, C2V_42_438, C2V_42_535, C2V_42_616, C2V_42_772, C2V_42_848, C2V_42_881, C2V_42_943, C2V_42_978, C2V_42_1045, C2V_42_1061, C2V_42_1111, C2V_42_1193, C2V_42_1194, C2V_43_12, C2V_43_96, C2V_43_116, C2V_43_177, C2V_43_239, C2V_43_282, C2V_43_382, C2V_43_388, C2V_43_485, C2V_43_721, C2V_43_769, C2V_43_817, C2V_43_906, C2V_43_947, C2V_43_981, C2V_43_1020, C2V_43_1094, C2V_43_1105, C2V_43_1194, C2V_43_1195, C2V_44_21, C2V_44_70, C2V_44_126, C2V_44_174, C2V_44_203, C2V_44_272, C2V_44_323, C2V_44_430, C2V_44_519, C2V_44_631, C2V_44_692, C2V_44_860, C2V_44_902, C2V_44_917, C2V_44_996, C2V_44_1028, C2V_44_1095, C2V_44_1126, C2V_44_1195, C2V_44_1196, C2V_45_16, C2V_45_91, C2V_45_108, C2V_45_190, C2V_45_208, C2V_45_275, C2V_45_372, C2V_45_427, C2V_45_538, C2V_45_595, C2V_45_671, C2V_45_727, C2V_45_906, C2V_45_950, C2V_45_975, C2V_45_1035, C2V_45_1065, C2V_45_1110, C2V_45_1196, C2V_45_1197, C2V_46_35, C2V_46_94, C2V_46_133, C2V_46_189, C2V_46_206, C2V_46_260, C2V_46_436, C2V_46_524, C2V_46_560, C2V_46_622, C2V_46_647, C2V_46_693, C2V_46_910, C2V_46_934, C2V_46_970, C2V_46_1048, C2V_46_1075, C2V_46_1139, C2V_46_1197, C2V_46_1198, C2V_47_6, C2V_47_64, C2V_47_99, C2V_47_170, C2V_47_234, C2V_47_252, C2V_47_301, C2V_47_368, C2V_47_447, C2V_47_681, C2V_47_745, C2V_47_799, C2V_47_877, C2V_47_925, C2V_47_968, C2V_47_1020, C2V_47_1069, C2V_47_1117, C2V_47_1198, C2V_47_1199, C2V_48_37, C2V_48_61, C2V_48_101, C2V_48_169, C2V_48_203, C2V_48_282, C2V_48_335, C2V_48_439, C2V_48_536, C2V_48_617, C2V_48_773, C2V_48_849, C2V_48_882, C2V_48_944, C2V_48_979, C2V_48_1046, C2V_48_1062, C2V_48_1112, C2V_48_1199, C2V_48_1200, C2V_49_13, C2V_49_49, C2V_49_117, C2V_49_178, C2V_49_240, C2V_49_283, C2V_49_383, C2V_49_389, C2V_49_486, C2V_49_722, C2V_49_770, C2V_49_818, C2V_49_907, C2V_49_948, C2V_49_982, C2V_49_1021, C2V_49_1095, C2V_49_1106, C2V_49_1200, C2V_49_1201, C2V_50_22, C2V_50_71, C2V_50_127, C2V_50_175, C2V_50_204, C2V_50_273, C2V_50_324, C2V_50_431, C2V_50_520, C2V_50_632, C2V_50_693, C2V_50_861, C2V_50_903, C2V_50_918, C2V_50_997, C2V_50_1029, C2V_50_1096, C2V_50_1127, C2V_50_1201, C2V_50_1202, C2V_51_17, C2V_51_92, C2V_51_109, C2V_51_191, C2V_51_209, C2V_51_276, C2V_51_373, C2V_51_428, C2V_51_539, C2V_51_596, C2V_51_672, C2V_51_728, C2V_51_907, C2V_51_951, C2V_51_976, C2V_51_1036, C2V_51_1066, C2V_51_1111, C2V_51_1202, C2V_51_1203, C2V_52_36, C2V_52_95, C2V_52_134, C2V_52_190, C2V_52_207, C2V_52_261, C2V_52_437, C2V_52_525, C2V_52_561, C2V_52_623, C2V_52_648, C2V_52_694, C2V_52_911, C2V_52_935, C2V_52_971, C2V_52_1049, C2V_52_1076, C2V_52_1140, C2V_52_1203, C2V_52_1204, C2V_53_7, C2V_53_65, C2V_53_100, C2V_53_171, C2V_53_235, C2V_53_253, C2V_53_302, C2V_53_369, C2V_53_448, C2V_53_682, C2V_53_746, C2V_53_800, C2V_53_878, C2V_53_926, C2V_53_969, C2V_53_1021, C2V_53_1070, C2V_53_1118, C2V_53_1204, C2V_53_1205, C2V_54_38, C2V_54_62, C2V_54_102, C2V_54_170, C2V_54_204, C2V_54_283, C2V_54_336, C2V_54_440, C2V_54_537, C2V_54_618, C2V_54_774, C2V_54_850, C2V_54_883, C2V_54_945, C2V_54_980, C2V_54_1047, C2V_54_1063, C2V_54_1113, C2V_54_1205, C2V_54_1206, C2V_55_14, C2V_55_50, C2V_55_118, C2V_55_179, C2V_55_193, C2V_55_284, C2V_55_384, C2V_55_390, C2V_55_487, C2V_55_723, C2V_55_771, C2V_55_819, C2V_55_908, C2V_55_949, C2V_55_983, C2V_55_1022, C2V_55_1096, C2V_55_1107, C2V_55_1206, C2V_55_1207, C2V_56_23, C2V_56_72, C2V_56_128, C2V_56_176, C2V_56_205, C2V_56_274, C2V_56_325, C2V_56_432, C2V_56_521, C2V_56_633, C2V_56_694, C2V_56_862, C2V_56_904, C2V_56_919, C2V_56_998, C2V_56_1030, C2V_56_1097, C2V_56_1128, C2V_56_1207, C2V_56_1208, C2V_57_18, C2V_57_93, C2V_57_110, C2V_57_192, C2V_57_210, C2V_57_277, C2V_57_374, C2V_57_429, C2V_57_540, C2V_57_597, C2V_57_625, C2V_57_729, C2V_57_908, C2V_57_952, C2V_57_977, C2V_57_1037, C2V_57_1067, C2V_57_1112, C2V_57_1208, C2V_57_1209, C2V_58_37, C2V_58_96, C2V_58_135, C2V_58_191, C2V_58_208, C2V_58_262, C2V_58_438, C2V_58_526, C2V_58_562, C2V_58_624, C2V_58_649, C2V_58_695, C2V_58_912, C2V_58_936, C2V_58_972, C2V_58_1050, C2V_58_1077, C2V_58_1141, C2V_58_1209, C2V_58_1210, C2V_59_8, C2V_59_66, C2V_59_101, C2V_59_172, C2V_59_236, C2V_59_254, C2V_59_303, C2V_59_370, C2V_59_449, C2V_59_683, C2V_59_747, C2V_59_801, C2V_59_879, C2V_59_927, C2V_59_970, C2V_59_1022, C2V_59_1071, C2V_59_1119, C2V_59_1210, C2V_59_1211, C2V_60_39, C2V_60_63, C2V_60_103, C2V_60_171, C2V_60_205, C2V_60_284, C2V_60_289, C2V_60_441, C2V_60_538, C2V_60_619, C2V_60_775, C2V_60_851, C2V_60_884, C2V_60_946, C2V_60_981, C2V_60_1048, C2V_60_1064, C2V_60_1114, C2V_60_1211, C2V_60_1212, C2V_61_15, C2V_61_51, C2V_61_119, C2V_61_180, C2V_61_194, C2V_61_285, C2V_61_337, C2V_61_391, C2V_61_488, C2V_61_724, C2V_61_772, C2V_61_820, C2V_61_909, C2V_61_950, C2V_61_984, C2V_61_1023, C2V_61_1097, C2V_61_1108, C2V_61_1212, C2V_61_1213, C2V_62_24, C2V_62_73, C2V_62_129, C2V_62_177, C2V_62_206, C2V_62_275, C2V_62_326, C2V_62_385, C2V_62_522, C2V_62_634, C2V_62_695, C2V_62_863, C2V_62_905, C2V_62_920, C2V_62_999, C2V_62_1031, C2V_62_1098, C2V_62_1129, C2V_62_1213, C2V_62_1214, C2V_63_19, C2V_63_94, C2V_63_111, C2V_63_145, C2V_63_211, C2V_63_278, C2V_63_375, C2V_63_430, C2V_63_541, C2V_63_598, C2V_63_626, C2V_63_730, C2V_63_909, C2V_63_953, C2V_63_978, C2V_63_1038, C2V_63_1068, C2V_63_1113, C2V_63_1214, C2V_63_1215, C2V_64_38, C2V_64_49, C2V_64_136, C2V_64_192, C2V_64_209, C2V_64_263, C2V_64_439, C2V_64_527, C2V_64_563, C2V_64_577, C2V_64_650, C2V_64_696, C2V_64_865, C2V_64_937, C2V_64_973, C2V_64_1051, C2V_64_1078, C2V_64_1142, C2V_64_1215, C2V_64_1216, C2V_65_9, C2V_65_67, C2V_65_102, C2V_65_173, C2V_65_237, C2V_65_255, C2V_65_304, C2V_65_371, C2V_65_450, C2V_65_684, C2V_65_748, C2V_65_802, C2V_65_880, C2V_65_928, C2V_65_971, C2V_65_1023, C2V_65_1072, C2V_65_1120, C2V_65_1216, C2V_65_1217, C2V_66_40, C2V_66_64, C2V_66_104, C2V_66_172, C2V_66_206, C2V_66_285, C2V_66_290, C2V_66_442, C2V_66_539, C2V_66_620, C2V_66_776, C2V_66_852, C2V_66_885, C2V_66_947, C2V_66_982, C2V_66_1049, C2V_66_1065, C2V_66_1115, C2V_66_1217, C2V_66_1218, C2V_67_16, C2V_67_52, C2V_67_120, C2V_67_181, C2V_67_195, C2V_67_286, C2V_67_338, C2V_67_392, C2V_67_489, C2V_67_725, C2V_67_773, C2V_67_821, C2V_67_910, C2V_67_951, C2V_67_985, C2V_67_1024, C2V_67_1098, C2V_67_1109, C2V_67_1218, C2V_67_1219, C2V_68_25, C2V_68_74, C2V_68_130, C2V_68_178, C2V_68_207, C2V_68_276, C2V_68_327, C2V_68_386, C2V_68_523, C2V_68_635, C2V_68_696, C2V_68_864, C2V_68_906, C2V_68_921, C2V_68_1000, C2V_68_1032, C2V_68_1099, C2V_68_1130, C2V_68_1219, C2V_68_1220, C2V_69_20, C2V_69_95, C2V_69_112, C2V_69_146, C2V_69_212, C2V_69_279, C2V_69_376, C2V_69_431, C2V_69_542, C2V_69_599, C2V_69_627, C2V_69_731, C2V_69_910, C2V_69_954, C2V_69_979, C2V_69_1039, C2V_69_1069, C2V_69_1114, C2V_69_1220, C2V_69_1221, C2V_70_39, C2V_70_50, C2V_70_137, C2V_70_145, C2V_70_210, C2V_70_264, C2V_70_440, C2V_70_528, C2V_70_564, C2V_70_578, C2V_70_651, C2V_70_697, C2V_70_866, C2V_70_938, C2V_70_974, C2V_70_1052, C2V_70_1079, C2V_70_1143, C2V_70_1221, C2V_70_1222, C2V_71_10, C2V_71_68, C2V_71_103, C2V_71_174, C2V_71_238, C2V_71_256, C2V_71_305, C2V_71_372, C2V_71_451, C2V_71_685, C2V_71_749, C2V_71_803, C2V_71_881, C2V_71_929, C2V_71_972, C2V_71_1024, C2V_71_1073, C2V_71_1121, C2V_71_1222, C2V_71_1223, C2V_72_41, C2V_72_65, C2V_72_105, C2V_72_173, C2V_72_207, C2V_72_286, C2V_72_291, C2V_72_443, C2V_72_540, C2V_72_621, C2V_72_777, C2V_72_853, C2V_72_886, C2V_72_948, C2V_72_983, C2V_72_1050, C2V_72_1066, C2V_72_1116, C2V_72_1223, C2V_72_1224, C2V_73_17, C2V_73_53, C2V_73_121, C2V_73_182, C2V_73_196, C2V_73_287, C2V_73_339, C2V_73_393, C2V_73_490, C2V_73_726, C2V_73_774, C2V_73_822, C2V_73_911, C2V_73_952, C2V_73_986, C2V_73_1025, C2V_73_1099, C2V_73_1110, C2V_73_1224, C2V_73_1225, C2V_74_26, C2V_74_75, C2V_74_131, C2V_74_179, C2V_74_208, C2V_74_277, C2V_74_328, C2V_74_387, C2V_74_524, C2V_74_636, C2V_74_697, C2V_74_817, C2V_74_907, C2V_74_922, C2V_74_1001, C2V_74_1033, C2V_74_1100, C2V_74_1131, C2V_74_1225, C2V_74_1226, C2V_75_21, C2V_75_96, C2V_75_113, C2V_75_147, C2V_75_213, C2V_75_280, C2V_75_377, C2V_75_432, C2V_75_543, C2V_75_600, C2V_75_628, C2V_75_732, C2V_75_911, C2V_75_955, C2V_75_980, C2V_75_1040, C2V_75_1070, C2V_75_1115, C2V_75_1226, C2V_75_1227, C2V_76_40, C2V_76_51, C2V_76_138, C2V_76_146, C2V_76_211, C2V_76_265, C2V_76_441, C2V_76_481, C2V_76_565, C2V_76_579, C2V_76_652, C2V_76_698, C2V_76_867, C2V_76_939, C2V_76_975, C2V_76_1053, C2V_76_1080, C2V_76_1144, C2V_76_1227, C2V_76_1228, C2V_77_11, C2V_77_69, C2V_77_104, C2V_77_175, C2V_77_239, C2V_77_257, C2V_77_306, C2V_77_373, C2V_77_452, C2V_77_686, C2V_77_750, C2V_77_804, C2V_77_882, C2V_77_930, C2V_77_973, C2V_77_1025, C2V_77_1074, C2V_77_1122, C2V_77_1228, C2V_77_1229, C2V_78_42, C2V_78_66, C2V_78_106, C2V_78_174, C2V_78_208, C2V_78_287, C2V_78_292, C2V_78_444, C2V_78_541, C2V_78_622, C2V_78_778, C2V_78_854, C2V_78_887, C2V_78_949, C2V_78_984, C2V_78_1051, C2V_78_1067, C2V_78_1117, C2V_78_1229, C2V_78_1230, C2V_79_18, C2V_79_54, C2V_79_122, C2V_79_183, C2V_79_197, C2V_79_288, C2V_79_340, C2V_79_394, C2V_79_491, C2V_79_727, C2V_79_775, C2V_79_823, C2V_79_912, C2V_79_953, C2V_79_987, C2V_79_1026, C2V_79_1100, C2V_79_1111, C2V_79_1230, C2V_79_1231, C2V_80_27, C2V_80_76, C2V_80_132, C2V_80_180, C2V_80_209, C2V_80_278, C2V_80_329, C2V_80_388, C2V_80_525, C2V_80_637, C2V_80_698, C2V_80_818, C2V_80_908, C2V_80_923, C2V_80_1002, C2V_80_1034, C2V_80_1101, C2V_80_1132, C2V_80_1231, C2V_80_1232, C2V_81_22, C2V_81_49, C2V_81_114, C2V_81_148, C2V_81_214, C2V_81_281, C2V_81_378, C2V_81_385, C2V_81_544, C2V_81_601, C2V_81_629, C2V_81_733, C2V_81_912, C2V_81_956, C2V_81_981, C2V_81_1041, C2V_81_1071, C2V_81_1116, C2V_81_1232, C2V_81_1233, C2V_82_41, C2V_82_52, C2V_82_139, C2V_82_147, C2V_82_212, C2V_82_266, C2V_82_442, C2V_82_482, C2V_82_566, C2V_82_580, C2V_82_653, C2V_82_699, C2V_82_868, C2V_82_940, C2V_82_976, C2V_82_1054, C2V_82_1081, C2V_82_1145, C2V_82_1233, C2V_82_1234, C2V_83_12, C2V_83_70, C2V_83_105, C2V_83_176, C2V_83_240, C2V_83_258, C2V_83_307, C2V_83_374, C2V_83_453, C2V_83_687, C2V_83_751, C2V_83_805, C2V_83_883, C2V_83_931, C2V_83_974, C2V_83_1026, C2V_83_1075, C2V_83_1123, C2V_83_1234, C2V_83_1235, C2V_84_43, C2V_84_67, C2V_84_107, C2V_84_175, C2V_84_209, C2V_84_288, C2V_84_293, C2V_84_445, C2V_84_542, C2V_84_623, C2V_84_779, C2V_84_855, C2V_84_888, C2V_84_950, C2V_84_985, C2V_84_1052, C2V_84_1068, C2V_84_1118, C2V_84_1235, C2V_84_1236, C2V_85_19, C2V_85_55, C2V_85_123, C2V_85_184, C2V_85_198, C2V_85_241, C2V_85_341, C2V_85_395, C2V_85_492, C2V_85_728, C2V_85_776, C2V_85_824, C2V_85_865, C2V_85_954, C2V_85_988, C2V_85_1027, C2V_85_1101, C2V_85_1112, C2V_85_1236, C2V_85_1237, C2V_86_28, C2V_86_77, C2V_86_133, C2V_86_181, C2V_86_210, C2V_86_279, C2V_86_330, C2V_86_389, C2V_86_526, C2V_86_638, C2V_86_699, C2V_86_819, C2V_86_909, C2V_86_924, C2V_86_1003, C2V_86_1035, C2V_86_1102, C2V_86_1133, C2V_86_1237, C2V_86_1238, C2V_87_23, C2V_87_50, C2V_87_115, C2V_87_149, C2V_87_215, C2V_87_282, C2V_87_379, C2V_87_386, C2V_87_545, C2V_87_602, C2V_87_630, C2V_87_734, C2V_87_865, C2V_87_957, C2V_87_982, C2V_87_1042, C2V_87_1072, C2V_87_1117, C2V_87_1238, C2V_87_1239, C2V_88_42, C2V_88_53, C2V_88_140, C2V_88_148, C2V_88_213, C2V_88_267, C2V_88_443, C2V_88_483, C2V_88_567, C2V_88_581, C2V_88_654, C2V_88_700, C2V_88_869, C2V_88_941, C2V_88_977, C2V_88_1055, C2V_88_1082, C2V_88_1146, C2V_88_1239, C2V_88_1240, C2V_89_13, C2V_89_71, C2V_89_106, C2V_89_177, C2V_89_193, C2V_89_259, C2V_89_308, C2V_89_375, C2V_89_454, C2V_89_688, C2V_89_752, C2V_89_806, C2V_89_884, C2V_89_932, C2V_89_975, C2V_89_1027, C2V_89_1076, C2V_89_1124, C2V_89_1240, C2V_89_1241, C2V_90_44, C2V_90_68, C2V_90_108, C2V_90_176, C2V_90_210, C2V_90_241, C2V_90_294, C2V_90_446, C2V_90_543, C2V_90_624, C2V_90_780, C2V_90_856, C2V_90_889, C2V_90_951, C2V_90_986, C2V_90_1053, C2V_90_1069, C2V_90_1119, C2V_90_1241, C2V_90_1242, C2V_91_20, C2V_91_56, C2V_91_124, C2V_91_185, C2V_91_199, C2V_91_242, C2V_91_342, C2V_91_396, C2V_91_493, C2V_91_729, C2V_91_777, C2V_91_825, C2V_91_866, C2V_91_955, C2V_91_989, C2V_91_1028, C2V_91_1102, C2V_91_1113, C2V_91_1242, C2V_91_1243, C2V_92_29, C2V_92_78, C2V_92_134, C2V_92_182, C2V_92_211, C2V_92_280, C2V_92_331, C2V_92_390, C2V_92_527, C2V_92_639, C2V_92_700, C2V_92_820, C2V_92_910, C2V_92_925, C2V_92_1004, C2V_92_1036, C2V_92_1103, C2V_92_1134, C2V_92_1243, C2V_92_1244, C2V_93_24, C2V_93_51, C2V_93_116, C2V_93_150, C2V_93_216, C2V_93_283, C2V_93_380, C2V_93_387, C2V_93_546, C2V_93_603, C2V_93_631, C2V_93_735, C2V_93_866, C2V_93_958, C2V_93_983, C2V_93_1043, C2V_93_1073, C2V_93_1118, C2V_93_1244, C2V_93_1245, C2V_94_43, C2V_94_54, C2V_94_141, C2V_94_149, C2V_94_214, C2V_94_268, C2V_94_444, C2V_94_484, C2V_94_568, C2V_94_582, C2V_94_655, C2V_94_701, C2V_94_870, C2V_94_942, C2V_94_978, C2V_94_1056, C2V_94_1083, C2V_94_1147, C2V_94_1245, C2V_94_1246, C2V_95_14, C2V_95_72, C2V_95_107, C2V_95_178, C2V_95_194, C2V_95_260, C2V_95_309, C2V_95_376, C2V_95_455, C2V_95_689, C2V_95_753, C2V_95_807, C2V_95_885, C2V_95_933, C2V_95_976, C2V_95_1028, C2V_95_1077, C2V_95_1125, C2V_95_1246, C2V_95_1247, C2V_96_45, C2V_96_69, C2V_96_109, C2V_96_177, C2V_96_211, C2V_96_242, C2V_96_295, C2V_96_447, C2V_96_544, C2V_96_577, C2V_96_781, C2V_96_857, C2V_96_890, C2V_96_952, C2V_96_987, C2V_96_1054, C2V_96_1070, C2V_96_1120, C2V_96_1247, C2V_96_1248, C2V_97_21, C2V_97_57, C2V_97_125, C2V_97_186, C2V_97_200, C2V_97_243, C2V_97_343, C2V_97_397, C2V_97_494, C2V_97_730, C2V_97_778, C2V_97_826, C2V_97_867, C2V_97_956, C2V_97_990, C2V_97_1029, C2V_97_1103, C2V_97_1114, C2V_97_1248, C2V_97_1249, C2V_98_30, C2V_98_79, C2V_98_135, C2V_98_183, C2V_98_212, C2V_98_281, C2V_98_332, C2V_98_391, C2V_98_528, C2V_98_640, C2V_98_701, C2V_98_821, C2V_98_911, C2V_98_926, C2V_98_1005, C2V_98_1037, C2V_98_1104, C2V_98_1135, C2V_98_1249, C2V_98_1250, C2V_99_25, C2V_99_52, C2V_99_117, C2V_99_151, C2V_99_217, C2V_99_284, C2V_99_381, C2V_99_388, C2V_99_547, C2V_99_604, C2V_99_632, C2V_99_736, C2V_99_867, C2V_99_959, C2V_99_984, C2V_99_1044, C2V_99_1074, C2V_99_1119, C2V_99_1250, C2V_99_1251, C2V_100_44, C2V_100_55, C2V_100_142, C2V_100_150, C2V_100_215, C2V_100_269, C2V_100_445, C2V_100_485, C2V_100_569, C2V_100_583, C2V_100_656, C2V_100_702, C2V_100_871, C2V_100_943, C2V_100_979, C2V_100_1009, C2V_100_1084, C2V_100_1148, C2V_100_1251, C2V_100_1252, C2V_101_15, C2V_101_73, C2V_101_108, C2V_101_179, C2V_101_195, C2V_101_261, C2V_101_310, C2V_101_377, C2V_101_456, C2V_101_690, C2V_101_754, C2V_101_808, C2V_101_886, C2V_101_934, C2V_101_977, C2V_101_1029, C2V_101_1078, C2V_101_1126, C2V_101_1252, C2V_101_1253, C2V_102_46, C2V_102_70, C2V_102_110, C2V_102_178, C2V_102_212, C2V_102_243, C2V_102_296, C2V_102_448, C2V_102_545, C2V_102_578, C2V_102_782, C2V_102_858, C2V_102_891, C2V_102_953, C2V_102_988, C2V_102_1055, C2V_102_1071, C2V_102_1121, C2V_102_1253, C2V_102_1254, C2V_103_22, C2V_103_58, C2V_103_126, C2V_103_187, C2V_103_201, C2V_103_244, C2V_103_344, C2V_103_398, C2V_103_495, C2V_103_731, C2V_103_779, C2V_103_827, C2V_103_868, C2V_103_957, C2V_103_991, C2V_103_1030, C2V_103_1104, C2V_103_1115, C2V_103_1254, C2V_103_1255, C2V_104_31, C2V_104_80, C2V_104_136, C2V_104_184, C2V_104_213, C2V_104_282, C2V_104_333, C2V_104_392, C2V_104_481, C2V_104_641, C2V_104_702, C2V_104_822, C2V_104_912, C2V_104_927, C2V_104_1006, C2V_104_1038, C2V_104_1057, C2V_104_1136, C2V_104_1255, C2V_104_1256, C2V_105_26, C2V_105_53, C2V_105_118, C2V_105_152, C2V_105_218, C2V_105_285, C2V_105_382, C2V_105_389, C2V_105_548, C2V_105_605, C2V_105_633, C2V_105_737, C2V_105_868, C2V_105_960, C2V_105_985, C2V_105_1045, C2V_105_1075, C2V_105_1120, C2V_105_1256, C2V_105_1257, C2V_106_45, C2V_106_56, C2V_106_143, C2V_106_151, C2V_106_216, C2V_106_270, C2V_106_446, C2V_106_486, C2V_106_570, C2V_106_584, C2V_106_657, C2V_106_703, C2V_106_872, C2V_106_944, C2V_106_980, C2V_106_1010, C2V_106_1085, C2V_106_1149, C2V_106_1257, C2V_106_1258, C2V_107_16, C2V_107_74, C2V_107_109, C2V_107_180, C2V_107_196, C2V_107_262, C2V_107_311, C2V_107_378, C2V_107_457, C2V_107_691, C2V_107_755, C2V_107_809, C2V_107_887, C2V_107_935, C2V_107_978, C2V_107_1030, C2V_107_1079, C2V_107_1127, C2V_107_1258, C2V_107_1259, C2V_108_47, C2V_108_71, C2V_108_111, C2V_108_179, C2V_108_213, C2V_108_244, C2V_108_297, C2V_108_449, C2V_108_546, C2V_108_579, C2V_108_783, C2V_108_859, C2V_108_892, C2V_108_954, C2V_108_989, C2V_108_1056, C2V_108_1072, C2V_108_1122, C2V_108_1259, C2V_108_1260, C2V_109_23, C2V_109_59, C2V_109_127, C2V_109_188, C2V_109_202, C2V_109_245, C2V_109_345, C2V_109_399, C2V_109_496, C2V_109_732, C2V_109_780, C2V_109_828, C2V_109_869, C2V_109_958, C2V_109_992, C2V_109_1031, C2V_109_1057, C2V_109_1116, C2V_109_1260, C2V_109_1261, C2V_110_32, C2V_110_81, C2V_110_137, C2V_110_185, C2V_110_214, C2V_110_283, C2V_110_334, C2V_110_393, C2V_110_482, C2V_110_642, C2V_110_703, C2V_110_823, C2V_110_865, C2V_110_928, C2V_110_1007, C2V_110_1039, C2V_110_1058, C2V_110_1137, C2V_110_1261, C2V_110_1262, C2V_111_27, C2V_111_54, C2V_111_119, C2V_111_153, C2V_111_219, C2V_111_286, C2V_111_383, C2V_111_390, C2V_111_549, C2V_111_606, C2V_111_634, C2V_111_738, C2V_111_869, C2V_111_913, C2V_111_986, C2V_111_1046, C2V_111_1076, C2V_111_1121, C2V_111_1262, C2V_111_1263, C2V_112_46, C2V_112_57, C2V_112_144, C2V_112_152, C2V_112_217, C2V_112_271, C2V_112_447, C2V_112_487, C2V_112_571, C2V_112_585, C2V_112_658, C2V_112_704, C2V_112_873, C2V_112_945, C2V_112_981, C2V_112_1011, C2V_112_1086, C2V_112_1150, C2V_112_1263, C2V_112_1264, C2V_113_17, C2V_113_75, C2V_113_110, C2V_113_181, C2V_113_197, C2V_113_263, C2V_113_312, C2V_113_379, C2V_113_458, C2V_113_692, C2V_113_756, C2V_113_810, C2V_113_888, C2V_113_936, C2V_113_979, C2V_113_1031, C2V_113_1080, C2V_113_1128, C2V_113_1264, C2V_113_1265, C2V_114_48, C2V_114_72, C2V_114_112, C2V_114_180, C2V_114_214, C2V_114_245, C2V_114_298, C2V_114_450, C2V_114_547, C2V_114_580, C2V_114_784, C2V_114_860, C2V_114_893, C2V_114_955, C2V_114_990, C2V_114_1009, C2V_114_1073, C2V_114_1123, C2V_114_1265, C2V_114_1266, C2V_115_24, C2V_115_60, C2V_115_128, C2V_115_189, C2V_115_203, C2V_115_246, C2V_115_346, C2V_115_400, C2V_115_497, C2V_115_733, C2V_115_781, C2V_115_829, C2V_115_870, C2V_115_959, C2V_115_993, C2V_115_1032, C2V_115_1058, C2V_115_1117, C2V_115_1266, C2V_115_1267, C2V_116_33, C2V_116_82, C2V_116_138, C2V_116_186, C2V_116_215, C2V_116_284, C2V_116_335, C2V_116_394, C2V_116_483, C2V_116_643, C2V_116_704, C2V_116_824, C2V_116_866, C2V_116_929, C2V_116_1008, C2V_116_1040, C2V_116_1059, C2V_116_1138, C2V_116_1267, C2V_116_1268, C2V_117_28, C2V_117_55, C2V_117_120, C2V_117_154, C2V_117_220, C2V_117_287, C2V_117_384, C2V_117_391, C2V_117_550, C2V_117_607, C2V_117_635, C2V_117_739, C2V_117_870, C2V_117_914, C2V_117_987, C2V_117_1047, C2V_117_1077, C2V_117_1122, C2V_117_1268, C2V_117_1269, C2V_118_47, C2V_118_58, C2V_118_97, C2V_118_153, C2V_118_218, C2V_118_272, C2V_118_448, C2V_118_488, C2V_118_572, C2V_118_586, C2V_118_659, C2V_118_705, C2V_118_874, C2V_118_946, C2V_118_982, C2V_118_1012, C2V_118_1087, C2V_118_1151, C2V_118_1269, C2V_118_1270, C2V_119_18, C2V_119_76, C2V_119_111, C2V_119_182, C2V_119_198, C2V_119_264, C2V_119_313, C2V_119_380, C2V_119_459, C2V_119_693, C2V_119_757, C2V_119_811, C2V_119_889, C2V_119_937, C2V_119_980, C2V_119_1032, C2V_119_1081, C2V_119_1129, C2V_119_1270, C2V_119_1271, C2V_120_1, C2V_120_73, C2V_120_113, C2V_120_181, C2V_120_215, C2V_120_246, C2V_120_299, C2V_120_451, C2V_120_548, C2V_120_581, C2V_120_785, C2V_120_861, C2V_120_894, C2V_120_956, C2V_120_991, C2V_120_1010, C2V_120_1074, C2V_120_1124, C2V_120_1271, C2V_120_1272, C2V_121_25, C2V_121_61, C2V_121_129, C2V_121_190, C2V_121_204, C2V_121_247, C2V_121_347, C2V_121_401, C2V_121_498, C2V_121_734, C2V_121_782, C2V_121_830, C2V_121_871, C2V_121_960, C2V_121_994, C2V_121_1033, C2V_121_1059, C2V_121_1118, C2V_121_1272, C2V_121_1273, C2V_122_34, C2V_122_83, C2V_122_139, C2V_122_187, C2V_122_216, C2V_122_285, C2V_122_336, C2V_122_395, C2V_122_484, C2V_122_644, C2V_122_705, C2V_122_825, C2V_122_867, C2V_122_930, C2V_122_961, C2V_122_1041, C2V_122_1060, C2V_122_1139, C2V_122_1273, C2V_122_1274, C2V_123_29, C2V_123_56, C2V_123_121, C2V_123_155, C2V_123_221, C2V_123_288, C2V_123_337, C2V_123_392, C2V_123_551, C2V_123_608, C2V_123_636, C2V_123_740, C2V_123_871, C2V_123_915, C2V_123_988, C2V_123_1048, C2V_123_1078, C2V_123_1123, C2V_123_1274, C2V_123_1275, C2V_124_48, C2V_124_59, C2V_124_98, C2V_124_154, C2V_124_219, C2V_124_273, C2V_124_449, C2V_124_489, C2V_124_573, C2V_124_587, C2V_124_660, C2V_124_706, C2V_124_875, C2V_124_947, C2V_124_983, C2V_124_1013, C2V_124_1088, C2V_124_1152, C2V_124_1275, C2V_124_1276, C2V_125_19, C2V_125_77, C2V_125_112, C2V_125_183, C2V_125_199, C2V_125_265, C2V_125_314, C2V_125_381, C2V_125_460, C2V_125_694, C2V_125_758, C2V_125_812, C2V_125_890, C2V_125_938, C2V_125_981, C2V_125_1033, C2V_125_1082, C2V_125_1130, C2V_125_1276, C2V_125_1277, C2V_126_2, C2V_126_74, C2V_126_114, C2V_126_182, C2V_126_216, C2V_126_247, C2V_126_300, C2V_126_452, C2V_126_549, C2V_126_582, C2V_126_786, C2V_126_862, C2V_126_895, C2V_126_957, C2V_126_992, C2V_126_1011, C2V_126_1075, C2V_126_1125, C2V_126_1277, C2V_126_1278, C2V_127_26, C2V_127_62, C2V_127_130, C2V_127_191, C2V_127_205, C2V_127_248, C2V_127_348, C2V_127_402, C2V_127_499, C2V_127_735, C2V_127_783, C2V_127_831, C2V_127_872, C2V_127_913, C2V_127_995, C2V_127_1034, C2V_127_1060, C2V_127_1119, C2V_127_1278, C2V_127_1279, C2V_128_35, C2V_128_84, C2V_128_140, C2V_128_188, C2V_128_217, C2V_128_286, C2V_128_289, C2V_128_396, C2V_128_485, C2V_128_645, C2V_128_706, C2V_128_826, C2V_128_868, C2V_128_931, C2V_128_962, C2V_128_1042, C2V_128_1061, C2V_128_1140, C2V_128_1279, C2V_128_1280, C2V_129_30, C2V_129_57, C2V_129_122, C2V_129_156, C2V_129_222, C2V_129_241, C2V_129_338, C2V_129_393, C2V_129_552, C2V_129_609, C2V_129_637, C2V_129_741, C2V_129_872, C2V_129_916, C2V_129_989, C2V_129_1049, C2V_129_1079, C2V_129_1124, C2V_129_1280, C2V_129_1281, C2V_130_1, C2V_130_60, C2V_130_99, C2V_130_155, C2V_130_220, C2V_130_274, C2V_130_450, C2V_130_490, C2V_130_574, C2V_130_588, C2V_130_661, C2V_130_707, C2V_130_876, C2V_130_948, C2V_130_984, C2V_130_1014, C2V_130_1089, C2V_130_1105, C2V_130_1281, C2V_130_1282, C2V_131_20, C2V_131_78, C2V_131_113, C2V_131_184, C2V_131_200, C2V_131_266, C2V_131_315, C2V_131_382, C2V_131_461, C2V_131_695, C2V_131_759, C2V_131_813, C2V_131_891, C2V_131_939, C2V_131_982, C2V_131_1034, C2V_131_1083, C2V_131_1131, C2V_131_1282, C2V_131_1283, C2V_132_3, C2V_132_75, C2V_132_115, C2V_132_183, C2V_132_217, C2V_132_248, C2V_132_301, C2V_132_453, C2V_132_550, C2V_132_583, C2V_132_787, C2V_132_863, C2V_132_896, C2V_132_958, C2V_132_993, C2V_132_1012, C2V_132_1076, C2V_132_1126, C2V_132_1283, C2V_132_1284, C2V_133_27, C2V_133_63, C2V_133_131, C2V_133_192, C2V_133_206, C2V_133_249, C2V_133_349, C2V_133_403, C2V_133_500, C2V_133_736, C2V_133_784, C2V_133_832, C2V_133_873, C2V_133_914, C2V_133_996, C2V_133_1035, C2V_133_1061, C2V_133_1120, C2V_133_1284, C2V_133_1285, C2V_134_36, C2V_134_85, C2V_134_141, C2V_134_189, C2V_134_218, C2V_134_287, C2V_134_290, C2V_134_397, C2V_134_486, C2V_134_646, C2V_134_707, C2V_134_827, C2V_134_869, C2V_134_932, C2V_134_963, C2V_134_1043, C2V_134_1062, C2V_134_1141, C2V_134_1285, C2V_134_1286, C2V_135_31, C2V_135_58, C2V_135_123, C2V_135_157, C2V_135_223, C2V_135_242, C2V_135_339, C2V_135_394, C2V_135_553, C2V_135_610, C2V_135_638, C2V_135_742, C2V_135_873, C2V_135_917, C2V_135_990, C2V_135_1050, C2V_135_1080, C2V_135_1125, C2V_135_1286, C2V_135_1287, C2V_136_2, C2V_136_61, C2V_136_100, C2V_136_156, C2V_136_221, C2V_136_275, C2V_136_451, C2V_136_491, C2V_136_575, C2V_136_589, C2V_136_662, C2V_136_708, C2V_136_877, C2V_136_949, C2V_136_985, C2V_136_1015, C2V_136_1090, C2V_136_1106, C2V_136_1287, C2V_136_1288, C2V_137_21, C2V_137_79, C2V_137_114, C2V_137_185, C2V_137_201, C2V_137_267, C2V_137_316, C2V_137_383, C2V_137_462, C2V_137_696, C2V_137_760, C2V_137_814, C2V_137_892, C2V_137_940, C2V_137_983, C2V_137_1035, C2V_137_1084, C2V_137_1132, C2V_137_1288, C2V_137_1289, C2V_138_4, C2V_138_76, C2V_138_116, C2V_138_184, C2V_138_218, C2V_138_249, C2V_138_302, C2V_138_454, C2V_138_551, C2V_138_584, C2V_138_788, C2V_138_864, C2V_138_897, C2V_138_959, C2V_138_994, C2V_138_1013, C2V_138_1077, C2V_138_1127, C2V_138_1289, C2V_138_1290, C2V_139_28, C2V_139_64, C2V_139_132, C2V_139_145, C2V_139_207, C2V_139_250, C2V_139_350, C2V_139_404, C2V_139_501, C2V_139_737, C2V_139_785, C2V_139_833, C2V_139_874, C2V_139_915, C2V_139_997, C2V_139_1036, C2V_139_1062, C2V_139_1121, C2V_139_1290, C2V_139_1291, C2V_140_37, C2V_140_86, C2V_140_142, C2V_140_190, C2V_140_219, C2V_140_288, C2V_140_291, C2V_140_398, C2V_140_487, C2V_140_647, C2V_140_708, C2V_140_828, C2V_140_870, C2V_140_933, C2V_140_964, C2V_140_1044, C2V_140_1063, C2V_140_1142, C2V_140_1291, C2V_140_1292, C2V_141_32, C2V_141_59, C2V_141_124, C2V_141_158, C2V_141_224, C2V_141_243, C2V_141_340, C2V_141_395, C2V_141_554, C2V_141_611, C2V_141_639, C2V_141_743, C2V_141_874, C2V_141_918, C2V_141_991, C2V_141_1051, C2V_141_1081, C2V_141_1126, C2V_141_1292, C2V_141_1293, C2V_142_3, C2V_142_62, C2V_142_101, C2V_142_157, C2V_142_222, C2V_142_276, C2V_142_452, C2V_142_492, C2V_142_576, C2V_142_590, C2V_142_663, C2V_142_709, C2V_142_878, C2V_142_950, C2V_142_986, C2V_142_1016, C2V_142_1091, C2V_142_1107, C2V_142_1293, C2V_142_1294, C2V_143_22, C2V_143_80, C2V_143_115, C2V_143_186, C2V_143_202, C2V_143_268, C2V_143_317, C2V_143_384, C2V_143_463, C2V_143_697, C2V_143_761, C2V_143_815, C2V_143_893, C2V_143_941, C2V_143_984, C2V_143_1036, C2V_143_1085, C2V_143_1133, C2V_143_1294, C2V_143_1295, C2V_144_5, C2V_144_77, C2V_144_117, C2V_144_185, C2V_144_219, C2V_144_250, C2V_144_303, C2V_144_455, C2V_144_552, C2V_144_585, C2V_144_789, C2V_144_817, C2V_144_898, C2V_144_960, C2V_144_995, C2V_144_1014, C2V_144_1078, C2V_144_1128, C2V_144_1295, C2V_144_1296, C2V_145_29, C2V_145_65, C2V_145_133, C2V_145_146, C2V_145_208, C2V_145_251, C2V_145_351, C2V_145_405, C2V_145_502, C2V_145_738, C2V_145_786, C2V_145_834, C2V_145_875, C2V_145_916, C2V_145_998, C2V_145_1037, C2V_145_1063, C2V_145_1122, C2V_145_1296, C2V_145_1297, C2V_146_38, C2V_146_87, C2V_146_143, C2V_146_191, C2V_146_220, C2V_146_241, C2V_146_292, C2V_146_399, C2V_146_488, C2V_146_648, C2V_146_709, C2V_146_829, C2V_146_871, C2V_146_934, C2V_146_965, C2V_146_1045, C2V_146_1064, C2V_146_1143, C2V_146_1297, C2V_146_1298, C2V_147_33, C2V_147_60, C2V_147_125, C2V_147_159, C2V_147_225, C2V_147_244, C2V_147_341, C2V_147_396, C2V_147_555, C2V_147_612, C2V_147_640, C2V_147_744, C2V_147_875, C2V_147_919, C2V_147_992, C2V_147_1052, C2V_147_1082, C2V_147_1127, C2V_147_1298, C2V_147_1299, C2V_148_4, C2V_148_63, C2V_148_102, C2V_148_158, C2V_148_223, C2V_148_277, C2V_148_453, C2V_148_493, C2V_148_529, C2V_148_591, C2V_148_664, C2V_148_710, C2V_148_879, C2V_148_951, C2V_148_987, C2V_148_1017, C2V_148_1092, C2V_148_1108, C2V_148_1299, C2V_148_1300, C2V_149_23, C2V_149_81, C2V_149_116, C2V_149_187, C2V_149_203, C2V_149_269, C2V_149_318, C2V_149_337, C2V_149_464, C2V_149_698, C2V_149_762, C2V_149_816, C2V_149_894, C2V_149_942, C2V_149_985, C2V_149_1037, C2V_149_1086, C2V_149_1134, C2V_149_1300, C2V_149_1301, C2V_150_6, C2V_150_78, C2V_150_118, C2V_150_186, C2V_150_220, C2V_150_251, C2V_150_304, C2V_150_456, C2V_150_553, C2V_150_586, C2V_150_790, C2V_150_818, C2V_150_899, C2V_150_913, C2V_150_996, C2V_150_1015, C2V_150_1079, C2V_150_1129, C2V_150_1301, C2V_150_1302, C2V_151_30, C2V_151_66, C2V_151_134, C2V_151_147, C2V_151_209, C2V_151_252, C2V_151_352, C2V_151_406, C2V_151_503, C2V_151_739, C2V_151_787, C2V_151_835, C2V_151_876, C2V_151_917, C2V_151_999, C2V_151_1038, C2V_151_1064, C2V_151_1123, C2V_151_1302, C2V_151_1303, C2V_152_39, C2V_152_88, C2V_152_144, C2V_152_192, C2V_152_221, C2V_152_242, C2V_152_293, C2V_152_400, C2V_152_489, C2V_152_649, C2V_152_710, C2V_152_830, C2V_152_872, C2V_152_935, C2V_152_966, C2V_152_1046, C2V_152_1065, C2V_152_1144, C2V_152_1303, C2V_152_1304, C2V_153_34, C2V_153_61, C2V_153_126, C2V_153_160, C2V_153_226, C2V_153_245, C2V_153_342, C2V_153_397, C2V_153_556, C2V_153_613, C2V_153_641, C2V_153_745, C2V_153_876, C2V_153_920, C2V_153_993, C2V_153_1053, C2V_153_1083, C2V_153_1128, C2V_153_1304, C2V_153_1305, C2V_154_5, C2V_154_64, C2V_154_103, C2V_154_159, C2V_154_224, C2V_154_278, C2V_154_454, C2V_154_494, C2V_154_530, C2V_154_592, C2V_154_665, C2V_154_711, C2V_154_880, C2V_154_952, C2V_154_988, C2V_154_1018, C2V_154_1093, C2V_154_1109, C2V_154_1305, C2V_154_1306, C2V_155_24, C2V_155_82, C2V_155_117, C2V_155_188, C2V_155_204, C2V_155_270, C2V_155_319, C2V_155_338, C2V_155_465, C2V_155_699, C2V_155_763, C2V_155_769, C2V_155_895, C2V_155_943, C2V_155_986, C2V_155_1038, C2V_155_1087, C2V_155_1135, C2V_155_1306, C2V_155_1307, C2V_156_7, C2V_156_79, C2V_156_119, C2V_156_187, C2V_156_221, C2V_156_252, C2V_156_305, C2V_156_457, C2V_156_554, C2V_156_587, C2V_156_791, C2V_156_819, C2V_156_900, C2V_156_914, C2V_156_997, C2V_156_1016, C2V_156_1080, C2V_156_1130, C2V_156_1307, C2V_156_1308, C2V_157_31, C2V_157_67, C2V_157_135, C2V_157_148, C2V_157_210, C2V_157_253, C2V_157_353, C2V_157_407, C2V_157_504, C2V_157_740, C2V_157_788, C2V_157_836, C2V_157_877, C2V_157_918, C2V_157_1000, C2V_157_1039, C2V_157_1065, C2V_157_1124, C2V_157_1308, C2V_157_1309, C2V_158_40, C2V_158_89, C2V_158_97, C2V_158_145, C2V_158_222, C2V_158_243, C2V_158_294, C2V_158_401, C2V_158_490, C2V_158_650, C2V_158_711, C2V_158_831, C2V_158_873, C2V_158_936, C2V_158_967, C2V_158_1047, C2V_158_1066, C2V_158_1145, C2V_158_1309, C2V_158_1310, C2V_159_35, C2V_159_62, C2V_159_127, C2V_159_161, C2V_159_227, C2V_159_246, C2V_159_343, C2V_159_398, C2V_159_557, C2V_159_614, C2V_159_642, C2V_159_746, C2V_159_877, C2V_159_921, C2V_159_994, C2V_159_1054, C2V_159_1084, C2V_159_1129, C2V_159_1310, C2V_159_1311, C2V_160_6, C2V_160_65, C2V_160_104, C2V_160_160, C2V_160_225, C2V_160_279, C2V_160_455, C2V_160_495, C2V_160_531, C2V_160_593, C2V_160_666, C2V_160_712, C2V_160_881, C2V_160_953, C2V_160_989, C2V_160_1019, C2V_160_1094, C2V_160_1110, C2V_160_1311, C2V_160_1312, C2V_161_25, C2V_161_83, C2V_161_118, C2V_161_189, C2V_161_205, C2V_161_271, C2V_161_320, C2V_161_339, C2V_161_466, C2V_161_700, C2V_161_764, C2V_161_770, C2V_161_896, C2V_161_944, C2V_161_987, C2V_161_1039, C2V_161_1088, C2V_161_1136, C2V_161_1312, C2V_161_1313, C2V_162_8, C2V_162_80, C2V_162_120, C2V_162_188, C2V_162_222, C2V_162_253, C2V_162_306, C2V_162_458, C2V_162_555, C2V_162_588, C2V_162_792, C2V_162_820, C2V_162_901, C2V_162_915, C2V_162_998, C2V_162_1017, C2V_162_1081, C2V_162_1131, C2V_162_1313, C2V_162_1314, C2V_163_32, C2V_163_68, C2V_163_136, C2V_163_149, C2V_163_211, C2V_163_254, C2V_163_354, C2V_163_408, C2V_163_505, C2V_163_741, C2V_163_789, C2V_163_837, C2V_163_878, C2V_163_919, C2V_163_1001, C2V_163_1040, C2V_163_1066, C2V_163_1125, C2V_163_1314, C2V_163_1315, C2V_164_41, C2V_164_90, C2V_164_98, C2V_164_146, C2V_164_223, C2V_164_244, C2V_164_295, C2V_164_402, C2V_164_491, C2V_164_651, C2V_164_712, C2V_164_832, C2V_164_874, C2V_164_937, C2V_164_968, C2V_164_1048, C2V_164_1067, C2V_164_1146, C2V_164_1315, C2V_164_1316, C2V_165_36, C2V_165_63, C2V_165_128, C2V_165_162, C2V_165_228, C2V_165_247, C2V_165_344, C2V_165_399, C2V_165_558, C2V_165_615, C2V_165_643, C2V_165_747, C2V_165_878, C2V_165_922, C2V_165_995, C2V_165_1055, C2V_165_1085, C2V_165_1130, C2V_165_1316, C2V_165_1317, C2V_166_7, C2V_166_66, C2V_166_105, C2V_166_161, C2V_166_226, C2V_166_280, C2V_166_456, C2V_166_496, C2V_166_532, C2V_166_594, C2V_166_667, C2V_166_713, C2V_166_882, C2V_166_954, C2V_166_990, C2V_166_1020, C2V_166_1095, C2V_166_1111, C2V_166_1317, C2V_166_1318, C2V_167_26, C2V_167_84, C2V_167_119, C2V_167_190, C2V_167_206, C2V_167_272, C2V_167_321, C2V_167_340, C2V_167_467, C2V_167_701, C2V_167_765, C2V_167_771, C2V_167_897, C2V_167_945, C2V_167_988, C2V_167_1040, C2V_167_1089, C2V_167_1137, C2V_167_1318, C2V_167_1319, C2V_168_9, C2V_168_81, C2V_168_121, C2V_168_189, C2V_168_223, C2V_168_254, C2V_168_307, C2V_168_459, C2V_168_556, C2V_168_589, C2V_168_793, C2V_168_821, C2V_168_902, C2V_168_916, C2V_168_999, C2V_168_1018, C2V_168_1082, C2V_168_1132, C2V_168_1319, C2V_168_1320, C2V_169_33, C2V_169_69, C2V_169_137, C2V_169_150, C2V_169_212, C2V_169_255, C2V_169_355, C2V_169_409, C2V_169_506, C2V_169_742, C2V_169_790, C2V_169_838, C2V_169_879, C2V_169_920, C2V_169_1002, C2V_169_1041, C2V_169_1067, C2V_169_1126, C2V_169_1320, C2V_169_1321, C2V_170_42, C2V_170_91, C2V_170_99, C2V_170_147, C2V_170_224, C2V_170_245, C2V_170_296, C2V_170_403, C2V_170_492, C2V_170_652, C2V_170_713, C2V_170_833, C2V_170_875, C2V_170_938, C2V_170_969, C2V_170_1049, C2V_170_1068, C2V_170_1147, C2V_170_1321, C2V_170_1322, C2V_171_37, C2V_171_64, C2V_171_129, C2V_171_163, C2V_171_229, C2V_171_248, C2V_171_345, C2V_171_400, C2V_171_559, C2V_171_616, C2V_171_644, C2V_171_748, C2V_171_879, C2V_171_923, C2V_171_996, C2V_171_1056, C2V_171_1086, C2V_171_1131, C2V_171_1322, C2V_171_1323, C2V_172_8, C2V_172_67, C2V_172_106, C2V_172_162, C2V_172_227, C2V_172_281, C2V_172_457, C2V_172_497, C2V_172_533, C2V_172_595, C2V_172_668, C2V_172_714, C2V_172_883, C2V_172_955, C2V_172_991, C2V_172_1021, C2V_172_1096, C2V_172_1112, C2V_172_1323, C2V_172_1324, C2V_173_27, C2V_173_85, C2V_173_120, C2V_173_191, C2V_173_207, C2V_173_273, C2V_173_322, C2V_173_341, C2V_173_468, C2V_173_702, C2V_173_766, C2V_173_772, C2V_173_898, C2V_173_946, C2V_173_989, C2V_173_1041, C2V_173_1090, C2V_173_1138, C2V_173_1324, C2V_173_1325, C2V_174_10, C2V_174_82, C2V_174_122, C2V_174_190, C2V_174_224, C2V_174_255, C2V_174_308, C2V_174_460, C2V_174_557, C2V_174_590, C2V_174_794, C2V_174_822, C2V_174_903, C2V_174_917, C2V_174_1000, C2V_174_1019, C2V_174_1083, C2V_174_1133, C2V_174_1325, C2V_174_1326, C2V_175_34, C2V_175_70, C2V_175_138, C2V_175_151, C2V_175_213, C2V_175_256, C2V_175_356, C2V_175_410, C2V_175_507, C2V_175_743, C2V_175_791, C2V_175_839, C2V_175_880, C2V_175_921, C2V_175_1003, C2V_175_1042, C2V_175_1068, C2V_175_1127, C2V_175_1326, C2V_175_1327, C2V_176_43, C2V_176_92, C2V_176_100, C2V_176_148, C2V_176_225, C2V_176_246, C2V_176_297, C2V_176_404, C2V_176_493, C2V_176_653, C2V_176_714, C2V_176_834, C2V_176_876, C2V_176_939, C2V_176_970, C2V_176_1050, C2V_176_1069, C2V_176_1148, C2V_176_1327, C2V_176_1328, C2V_177_38, C2V_177_65, C2V_177_130, C2V_177_164, C2V_177_230, C2V_177_249, C2V_177_346, C2V_177_401, C2V_177_560, C2V_177_617, C2V_177_645, C2V_177_749, C2V_177_880, C2V_177_924, C2V_177_997, C2V_177_1009, C2V_177_1087, C2V_177_1132, C2V_177_1328, C2V_177_1329, C2V_178_9, C2V_178_68, C2V_178_107, C2V_178_163, C2V_178_228, C2V_178_282, C2V_178_458, C2V_178_498, C2V_178_534, C2V_178_596, C2V_178_669, C2V_178_715, C2V_178_884, C2V_178_956, C2V_178_992, C2V_178_1022, C2V_178_1097, C2V_178_1113, C2V_178_1329, C2V_178_1330, C2V_179_28, C2V_179_86, C2V_179_121, C2V_179_192, C2V_179_208, C2V_179_274, C2V_179_323, C2V_179_342, C2V_179_469, C2V_179_703, C2V_179_767, C2V_179_773, C2V_179_899, C2V_179_947, C2V_179_990, C2V_179_1042, C2V_179_1091, C2V_179_1139, C2V_179_1330, C2V_179_1331, C2V_180_11, C2V_180_83, C2V_180_123, C2V_180_191, C2V_180_225, C2V_180_256, C2V_180_309, C2V_180_461, C2V_180_558, C2V_180_591, C2V_180_795, C2V_180_823, C2V_180_904, C2V_180_918, C2V_180_1001, C2V_180_1020, C2V_180_1084, C2V_180_1134, C2V_180_1331, C2V_180_1332, C2V_181_35, C2V_181_71, C2V_181_139, C2V_181_152, C2V_181_214, C2V_181_257, C2V_181_357, C2V_181_411, C2V_181_508, C2V_181_744, C2V_181_792, C2V_181_840, C2V_181_881, C2V_181_922, C2V_181_1004, C2V_181_1043, C2V_181_1069, C2V_181_1128, C2V_181_1332, C2V_181_1333, C2V_182_44, C2V_182_93, C2V_182_101, C2V_182_149, C2V_182_226, C2V_182_247, C2V_182_298, C2V_182_405, C2V_182_494, C2V_182_654, C2V_182_715, C2V_182_835, C2V_182_877, C2V_182_940, C2V_182_971, C2V_182_1051, C2V_182_1070, C2V_182_1149, C2V_182_1333, C2V_182_1334, C2V_183_39, C2V_183_66, C2V_183_131, C2V_183_165, C2V_183_231, C2V_183_250, C2V_183_347, C2V_183_402, C2V_183_561, C2V_183_618, C2V_183_646, C2V_183_750, C2V_183_881, C2V_183_925, C2V_183_998, C2V_183_1010, C2V_183_1088, C2V_183_1133, C2V_183_1334, C2V_183_1335, C2V_184_10, C2V_184_69, C2V_184_108, C2V_184_164, C2V_184_229, C2V_184_283, C2V_184_459, C2V_184_499, C2V_184_535, C2V_184_597, C2V_184_670, C2V_184_716, C2V_184_885, C2V_184_957, C2V_184_993, C2V_184_1023, C2V_184_1098, C2V_184_1114, C2V_184_1335, C2V_184_1336, C2V_185_29, C2V_185_87, C2V_185_122, C2V_185_145, C2V_185_209, C2V_185_275, C2V_185_324, C2V_185_343, C2V_185_470, C2V_185_704, C2V_185_768, C2V_185_774, C2V_185_900, C2V_185_948, C2V_185_991, C2V_185_1043, C2V_185_1092, C2V_185_1140, C2V_185_1336, C2V_185_1337, C2V_186_12, C2V_186_84, C2V_186_124, C2V_186_192, C2V_186_226, C2V_186_257, C2V_186_310, C2V_186_462, C2V_186_559, C2V_186_592, C2V_186_796, C2V_186_824, C2V_186_905, C2V_186_919, C2V_186_1002, C2V_186_1021, C2V_186_1085, C2V_186_1135, C2V_186_1337, C2V_186_1338, C2V_187_36, C2V_187_72, C2V_187_140, C2V_187_153, C2V_187_215, C2V_187_258, C2V_187_358, C2V_187_412, C2V_187_509, C2V_187_745, C2V_187_793, C2V_187_841, C2V_187_882, C2V_187_923, C2V_187_1005, C2V_187_1044, C2V_187_1070, C2V_187_1129, C2V_187_1338, C2V_187_1339, C2V_188_45, C2V_188_94, C2V_188_102, C2V_188_150, C2V_188_227, C2V_188_248, C2V_188_299, C2V_188_406, C2V_188_495, C2V_188_655, C2V_188_716, C2V_188_836, C2V_188_878, C2V_188_941, C2V_188_972, C2V_188_1052, C2V_188_1071, C2V_188_1150, C2V_188_1339, C2V_188_1340, C2V_189_40, C2V_189_67, C2V_189_132, C2V_189_166, C2V_189_232, C2V_189_251, C2V_189_348, C2V_189_403, C2V_189_562, C2V_189_619, C2V_189_647, C2V_189_751, C2V_189_882, C2V_189_926, C2V_189_999, C2V_189_1011, C2V_189_1089, C2V_189_1134, C2V_189_1340, C2V_189_1341, C2V_190_11, C2V_190_70, C2V_190_109, C2V_190_165, C2V_190_230, C2V_190_284, C2V_190_460, C2V_190_500, C2V_190_536, C2V_190_598, C2V_190_671, C2V_190_717, C2V_190_886, C2V_190_958, C2V_190_994, C2V_190_1024, C2V_190_1099, C2V_190_1115, C2V_190_1341, C2V_190_1342, C2V_191_30, C2V_191_88, C2V_191_123, C2V_191_146, C2V_191_210, C2V_191_276, C2V_191_325, C2V_191_344, C2V_191_471, C2V_191_705, C2V_191_721, C2V_191_775, C2V_191_901, C2V_191_949, C2V_191_992, C2V_191_1044, C2V_191_1093, C2V_191_1141, C2V_191_1342, C2V_191_1343, C2V_192_13, C2V_192_85, C2V_192_125, C2V_192_145, C2V_192_227, C2V_192_258, C2V_192_311, C2V_192_463, C2V_192_560, C2V_192_593, C2V_192_797, C2V_192_825, C2V_192_906, C2V_192_920, C2V_192_1003, C2V_192_1022, C2V_192_1086, C2V_192_1136, C2V_192_1343, C2V_192_1344, C2V_193_37, C2V_193_73, C2V_193_141, C2V_193_154, C2V_193_216, C2V_193_259, C2V_193_359, C2V_193_413, C2V_193_510, C2V_193_746, C2V_193_794, C2V_193_842, C2V_193_883, C2V_193_924, C2V_193_1006, C2V_193_1045, C2V_193_1071, C2V_193_1130, C2V_193_1344, C2V_193_1345, C2V_194_46, C2V_194_95, C2V_194_103, C2V_194_151, C2V_194_228, C2V_194_249, C2V_194_300, C2V_194_407, C2V_194_496, C2V_194_656, C2V_194_717, C2V_194_837, C2V_194_879, C2V_194_942, C2V_194_973, C2V_194_1053, C2V_194_1072, C2V_194_1151, C2V_194_1345, C2V_194_1346, C2V_195_41, C2V_195_68, C2V_195_133, C2V_195_167, C2V_195_233, C2V_195_252, C2V_195_349, C2V_195_404, C2V_195_563, C2V_195_620, C2V_195_648, C2V_195_752, C2V_195_883, C2V_195_927, C2V_195_1000, C2V_195_1012, C2V_195_1090, C2V_195_1135, C2V_195_1346, C2V_195_1347, C2V_196_12, C2V_196_71, C2V_196_110, C2V_196_166, C2V_196_231, C2V_196_285, C2V_196_461, C2V_196_501, C2V_196_537, C2V_196_599, C2V_196_672, C2V_196_718, C2V_196_887, C2V_196_959, C2V_196_995, C2V_196_1025, C2V_196_1100, C2V_196_1116, C2V_196_1347, C2V_196_1348, C2V_197_31, C2V_197_89, C2V_197_124, C2V_197_147, C2V_197_211, C2V_197_277, C2V_197_326, C2V_197_345, C2V_197_472, C2V_197_706, C2V_197_722, C2V_197_776, C2V_197_902, C2V_197_950, C2V_197_993, C2V_197_1045, C2V_197_1094, C2V_197_1142, C2V_197_1348, C2V_197_1349, C2V_198_14, C2V_198_86, C2V_198_126, C2V_198_146, C2V_198_228, C2V_198_259, C2V_198_312, C2V_198_464, C2V_198_561, C2V_198_594, C2V_198_798, C2V_198_826, C2V_198_907, C2V_198_921, C2V_198_1004, C2V_198_1023, C2V_198_1087, C2V_198_1137, C2V_198_1349, C2V_198_1350, C2V_199_38, C2V_199_74, C2V_199_142, C2V_199_155, C2V_199_217, C2V_199_260, C2V_199_360, C2V_199_414, C2V_199_511, C2V_199_747, C2V_199_795, C2V_199_843, C2V_199_884, C2V_199_925, C2V_199_1007, C2V_199_1046, C2V_199_1072, C2V_199_1131, C2V_199_1350, C2V_199_1351, C2V_200_47, C2V_200_96, C2V_200_104, C2V_200_152, C2V_200_229, C2V_200_250, C2V_200_301, C2V_200_408, C2V_200_497, C2V_200_657, C2V_200_718, C2V_200_838, C2V_200_880, C2V_200_943, C2V_200_974, C2V_200_1054, C2V_200_1073, C2V_200_1152, C2V_200_1351, C2V_200_1352, C2V_201_42, C2V_201_69, C2V_201_134, C2V_201_168, C2V_201_234, C2V_201_253, C2V_201_350, C2V_201_405, C2V_201_564, C2V_201_621, C2V_201_649, C2V_201_753, C2V_201_884, C2V_201_928, C2V_201_1001, C2V_201_1013, C2V_201_1091, C2V_201_1136, C2V_201_1352, C2V_201_1353, C2V_202_13, C2V_202_72, C2V_202_111, C2V_202_167, C2V_202_232, C2V_202_286, C2V_202_462, C2V_202_502, C2V_202_538, C2V_202_600, C2V_202_625, C2V_202_719, C2V_202_888, C2V_202_960, C2V_202_996, C2V_202_1026, C2V_202_1101, C2V_202_1117, C2V_202_1353, C2V_202_1354, C2V_203_32, C2V_203_90, C2V_203_125, C2V_203_148, C2V_203_212, C2V_203_278, C2V_203_327, C2V_203_346, C2V_203_473, C2V_203_707, C2V_203_723, C2V_203_777, C2V_203_903, C2V_203_951, C2V_203_994, C2V_203_1046, C2V_203_1095, C2V_203_1143, C2V_203_1354, C2V_203_1355, C2V_204_15, C2V_204_87, C2V_204_127, C2V_204_147, C2V_204_229, C2V_204_260, C2V_204_313, C2V_204_465, C2V_204_562, C2V_204_595, C2V_204_799, C2V_204_827, C2V_204_908, C2V_204_922, C2V_204_1005, C2V_204_1024, C2V_204_1088, C2V_204_1138, C2V_204_1355, C2V_204_1356, C2V_205_39, C2V_205_75, C2V_205_143, C2V_205_156, C2V_205_218, C2V_205_261, C2V_205_361, C2V_205_415, C2V_205_512, C2V_205_748, C2V_205_796, C2V_205_844, C2V_205_885, C2V_205_926, C2V_205_1008, C2V_205_1047, C2V_205_1073, C2V_205_1132, C2V_205_1356, C2V_205_1357, C2V_206_48, C2V_206_49, C2V_206_105, C2V_206_153, C2V_206_230, C2V_206_251, C2V_206_302, C2V_206_409, C2V_206_498, C2V_206_658, C2V_206_719, C2V_206_839, C2V_206_881, C2V_206_944, C2V_206_975, C2V_206_1055, C2V_206_1074, C2V_206_1105, C2V_206_1357, C2V_206_1358, C2V_207_43, C2V_207_70, C2V_207_135, C2V_207_169, C2V_207_235, C2V_207_254, C2V_207_351, C2V_207_406, C2V_207_565, C2V_207_622, C2V_207_650, C2V_207_754, C2V_207_885, C2V_207_929, C2V_207_1002, C2V_207_1014, C2V_207_1092, C2V_207_1137, C2V_207_1358, C2V_207_1359, C2V_208_14, C2V_208_73, C2V_208_112, C2V_208_168, C2V_208_233, C2V_208_287, C2V_208_463, C2V_208_503, C2V_208_539, C2V_208_601, C2V_208_626, C2V_208_720, C2V_208_889, C2V_208_913, C2V_208_997, C2V_208_1027, C2V_208_1102, C2V_208_1118, C2V_208_1359, C2V_208_1360, C2V_209_33, C2V_209_91, C2V_209_126, C2V_209_149, C2V_209_213, C2V_209_279, C2V_209_328, C2V_209_347, C2V_209_474, C2V_209_708, C2V_209_724, C2V_209_778, C2V_209_904, C2V_209_952, C2V_209_995, C2V_209_1047, C2V_209_1096, C2V_209_1144, C2V_209_1360, C2V_209_1361, C2V_210_16, C2V_210_88, C2V_210_128, C2V_210_148, C2V_210_230, C2V_210_261, C2V_210_314, C2V_210_466, C2V_210_563, C2V_210_596, C2V_210_800, C2V_210_828, C2V_210_909, C2V_210_923, C2V_210_1006, C2V_210_1025, C2V_210_1089, C2V_210_1139, C2V_210_1361, C2V_210_1362, C2V_211_40, C2V_211_76, C2V_211_144, C2V_211_157, C2V_211_219, C2V_211_262, C2V_211_362, C2V_211_416, C2V_211_513, C2V_211_749, C2V_211_797, C2V_211_845, C2V_211_886, C2V_211_927, C2V_211_961, C2V_211_1048, C2V_211_1074, C2V_211_1133, C2V_211_1362, C2V_211_1363, C2V_212_1, C2V_212_50, C2V_212_106, C2V_212_154, C2V_212_231, C2V_212_252, C2V_212_303, C2V_212_410, C2V_212_499, C2V_212_659, C2V_212_720, C2V_212_840, C2V_212_882, C2V_212_945, C2V_212_976, C2V_212_1056, C2V_212_1075, C2V_212_1106, C2V_212_1363, C2V_212_1364, C2V_213_44, C2V_213_71, C2V_213_136, C2V_213_170, C2V_213_236, C2V_213_255, C2V_213_352, C2V_213_407, C2V_213_566, C2V_213_623, C2V_213_651, C2V_213_755, C2V_213_886, C2V_213_930, C2V_213_1003, C2V_213_1015, C2V_213_1093, C2V_213_1138, C2V_213_1364, C2V_213_1365, C2V_214_15, C2V_214_74, C2V_214_113, C2V_214_169, C2V_214_234, C2V_214_288, C2V_214_464, C2V_214_504, C2V_214_540, C2V_214_602, C2V_214_627, C2V_214_673, C2V_214_890, C2V_214_914, C2V_214_998, C2V_214_1028, C2V_214_1103, C2V_214_1119, C2V_214_1365, C2V_214_1366, C2V_215_34, C2V_215_92, C2V_215_127, C2V_215_150, C2V_215_214, C2V_215_280, C2V_215_329, C2V_215_348, C2V_215_475, C2V_215_709, C2V_215_725, C2V_215_779, C2V_215_905, C2V_215_953, C2V_215_996, C2V_215_1048, C2V_215_1097, C2V_215_1145, C2V_215_1366, C2V_215_1367, C2V_216_17, C2V_216_89, C2V_216_129, C2V_216_149, C2V_216_231, C2V_216_262, C2V_216_315, C2V_216_467, C2V_216_564, C2V_216_597, C2V_216_801, C2V_216_829, C2V_216_910, C2V_216_924, C2V_216_1007, C2V_216_1026, C2V_216_1090, C2V_216_1140, C2V_216_1367, C2V_216_1368, C2V_217_41, C2V_217_77, C2V_217_97, C2V_217_158, C2V_217_220, C2V_217_263, C2V_217_363, C2V_217_417, C2V_217_514, C2V_217_750, C2V_217_798, C2V_217_846, C2V_217_887, C2V_217_928, C2V_217_962, C2V_217_1049, C2V_217_1075, C2V_217_1134, C2V_217_1368, C2V_217_1369, C2V_218_2, C2V_218_51, C2V_218_107, C2V_218_155, C2V_218_232, C2V_218_253, C2V_218_304, C2V_218_411, C2V_218_500, C2V_218_660, C2V_218_673, C2V_218_841, C2V_218_883, C2V_218_946, C2V_218_977, C2V_218_1009, C2V_218_1076, C2V_218_1107, C2V_218_1369, C2V_218_1370, C2V_219_45, C2V_219_72, C2V_219_137, C2V_219_171, C2V_219_237, C2V_219_256, C2V_219_353, C2V_219_408, C2V_219_567, C2V_219_624, C2V_219_652, C2V_219_756, C2V_219_887, C2V_219_931, C2V_219_1004, C2V_219_1016, C2V_219_1094, C2V_219_1139, C2V_219_1370, C2V_219_1371, C2V_220_16, C2V_220_75, C2V_220_114, C2V_220_170, C2V_220_235, C2V_220_241, C2V_220_465, C2V_220_505, C2V_220_541, C2V_220_603, C2V_220_628, C2V_220_674, C2V_220_891, C2V_220_915, C2V_220_999, C2V_220_1029, C2V_220_1104, C2V_220_1120, C2V_220_1371, C2V_220_1372, C2V_221_35, C2V_221_93, C2V_221_128, C2V_221_151, C2V_221_215, C2V_221_281, C2V_221_330, C2V_221_349, C2V_221_476, C2V_221_710, C2V_221_726, C2V_221_780, C2V_221_906, C2V_221_954, C2V_221_997, C2V_221_1049, C2V_221_1098, C2V_221_1146, C2V_221_1372, C2V_221_1373, C2V_222_18, C2V_222_90, C2V_222_130, C2V_222_150, C2V_222_232, C2V_222_263, C2V_222_316, C2V_222_468, C2V_222_565, C2V_222_598, C2V_222_802, C2V_222_830, C2V_222_911, C2V_222_925, C2V_222_1008, C2V_222_1027, C2V_222_1091, C2V_222_1141, C2V_222_1373, C2V_222_1374, C2V_223_42, C2V_223_78, C2V_223_98, C2V_223_159, C2V_223_221, C2V_223_264, C2V_223_364, C2V_223_418, C2V_223_515, C2V_223_751, C2V_223_799, C2V_223_847, C2V_223_888, C2V_223_929, C2V_223_963, C2V_223_1050, C2V_223_1076, C2V_223_1135, C2V_223_1374, C2V_223_1375, C2V_224_3, C2V_224_52, C2V_224_108, C2V_224_156, C2V_224_233, C2V_224_254, C2V_224_305, C2V_224_412, C2V_224_501, C2V_224_661, C2V_224_674, C2V_224_842, C2V_224_884, C2V_224_947, C2V_224_978, C2V_224_1010, C2V_224_1077, C2V_224_1108, C2V_224_1375, C2V_224_1376, C2V_225_46, C2V_225_73, C2V_225_138, C2V_225_172, C2V_225_238, C2V_225_257, C2V_225_354, C2V_225_409, C2V_225_568, C2V_225_577, C2V_225_653, C2V_225_757, C2V_225_888, C2V_225_932, C2V_225_1005, C2V_225_1017, C2V_225_1095, C2V_225_1140, C2V_225_1376, C2V_225_1377, C2V_226_17, C2V_226_76, C2V_226_115, C2V_226_171, C2V_226_236, C2V_226_242, C2V_226_466, C2V_226_506, C2V_226_542, C2V_226_604, C2V_226_629, C2V_226_675, C2V_226_892, C2V_226_916, C2V_226_1000, C2V_226_1030, C2V_226_1057, C2V_226_1121, C2V_226_1377, C2V_226_1378, C2V_227_36, C2V_227_94, C2V_227_129, C2V_227_152, C2V_227_216, C2V_227_282, C2V_227_331, C2V_227_350, C2V_227_477, C2V_227_711, C2V_227_727, C2V_227_781, C2V_227_907, C2V_227_955, C2V_227_998, C2V_227_1050, C2V_227_1099, C2V_227_1147, C2V_227_1378, C2V_227_1379, C2V_228_19, C2V_228_91, C2V_228_131, C2V_228_151, C2V_228_233, C2V_228_264, C2V_228_317, C2V_228_469, C2V_228_566, C2V_228_599, C2V_228_803, C2V_228_831, C2V_228_912, C2V_228_926, C2V_228_961, C2V_228_1028, C2V_228_1092, C2V_228_1142, C2V_228_1379, C2V_228_1380, C2V_229_43, C2V_229_79, C2V_229_99, C2V_229_160, C2V_229_222, C2V_229_265, C2V_229_365, C2V_229_419, C2V_229_516, C2V_229_752, C2V_229_800, C2V_229_848, C2V_229_889, C2V_229_930, C2V_229_964, C2V_229_1051, C2V_229_1077, C2V_229_1136, C2V_229_1380, C2V_229_1381, C2V_230_4, C2V_230_53, C2V_230_109, C2V_230_157, C2V_230_234, C2V_230_255, C2V_230_306, C2V_230_413, C2V_230_502, C2V_230_662, C2V_230_675, C2V_230_843, C2V_230_885, C2V_230_948, C2V_230_979, C2V_230_1011, C2V_230_1078, C2V_230_1109, C2V_230_1381, C2V_230_1382, C2V_231_47, C2V_231_74, C2V_231_139, C2V_231_173, C2V_231_239, C2V_231_258, C2V_231_355, C2V_231_410, C2V_231_569, C2V_231_578, C2V_231_654, C2V_231_758, C2V_231_889, C2V_231_933, C2V_231_1006, C2V_231_1018, C2V_231_1096, C2V_231_1141, C2V_231_1382, C2V_231_1383, C2V_232_18, C2V_232_77, C2V_232_116, C2V_232_172, C2V_232_237, C2V_232_243, C2V_232_467, C2V_232_507, C2V_232_543, C2V_232_605, C2V_232_630, C2V_232_676, C2V_232_893, C2V_232_917, C2V_232_1001, C2V_232_1031, C2V_232_1058, C2V_232_1122, C2V_232_1383, C2V_232_1384, C2V_233_37, C2V_233_95, C2V_233_130, C2V_233_153, C2V_233_217, C2V_233_283, C2V_233_332, C2V_233_351, C2V_233_478, C2V_233_712, C2V_233_728, C2V_233_782, C2V_233_908, C2V_233_956, C2V_233_999, C2V_233_1051, C2V_233_1100, C2V_233_1148, C2V_233_1384, C2V_233_1385, C2V_234_20, C2V_234_92, C2V_234_132, C2V_234_152, C2V_234_234, C2V_234_265, C2V_234_318, C2V_234_470, C2V_234_567, C2V_234_600, C2V_234_804, C2V_234_832, C2V_234_865, C2V_234_927, C2V_234_962, C2V_234_1029, C2V_234_1093, C2V_234_1143, C2V_234_1385, C2V_234_1386, C2V_235_44, C2V_235_80, C2V_235_100, C2V_235_161, C2V_235_223, C2V_235_266, C2V_235_366, C2V_235_420, C2V_235_517, C2V_235_753, C2V_235_801, C2V_235_849, C2V_235_890, C2V_235_931, C2V_235_965, C2V_235_1052, C2V_235_1078, C2V_235_1137, C2V_235_1386, C2V_235_1387, C2V_236_5, C2V_236_54, C2V_236_110, C2V_236_158, C2V_236_235, C2V_236_256, C2V_236_307, C2V_236_414, C2V_236_503, C2V_236_663, C2V_236_676, C2V_236_844, C2V_236_886, C2V_236_949, C2V_236_980, C2V_236_1012, C2V_236_1079, C2V_236_1110, C2V_236_1387, C2V_236_1388, C2V_237_48, C2V_237_75, C2V_237_140, C2V_237_174, C2V_237_240, C2V_237_259, C2V_237_356, C2V_237_411, C2V_237_570, C2V_237_579, C2V_237_655, C2V_237_759, C2V_237_890, C2V_237_934, C2V_237_1007, C2V_237_1019, C2V_237_1097, C2V_237_1142, C2V_237_1388, C2V_237_1389, C2V_238_19, C2V_238_78, C2V_238_117, C2V_238_173, C2V_238_238, C2V_238_244, C2V_238_468, C2V_238_508, C2V_238_544, C2V_238_606, C2V_238_631, C2V_238_677, C2V_238_894, C2V_238_918, C2V_238_1002, C2V_238_1032, C2V_238_1059, C2V_238_1123, C2V_238_1389, C2V_238_1390, C2V_239_38, C2V_239_96, C2V_239_131, C2V_239_154, C2V_239_218, C2V_239_284, C2V_239_333, C2V_239_352, C2V_239_479, C2V_239_713, C2V_239_729, C2V_239_783, C2V_239_909, C2V_239_957, C2V_239_1000, C2V_239_1052, C2V_239_1101, C2V_239_1149, C2V_239_1390, C2V_239_1391, C2V_240_21, C2V_240_93, C2V_240_133, C2V_240_153, C2V_240_235, C2V_240_266, C2V_240_319, C2V_240_471, C2V_240_568, C2V_240_601, C2V_240_805, C2V_240_833, C2V_240_866, C2V_240_928, C2V_240_963, C2V_240_1030, C2V_240_1094, C2V_240_1144, C2V_240_1391, C2V_240_1392, C2V_241_45, C2V_241_81, C2V_241_101, C2V_241_162, C2V_241_224, C2V_241_267, C2V_241_367, C2V_241_421, C2V_241_518, C2V_241_754, C2V_241_802, C2V_241_850, C2V_241_891, C2V_241_932, C2V_241_966, C2V_241_1053, C2V_241_1079, C2V_241_1138, C2V_241_1392, C2V_241_1393, C2V_242_6, C2V_242_55, C2V_242_111, C2V_242_159, C2V_242_236, C2V_242_257, C2V_242_308, C2V_242_415, C2V_242_504, C2V_242_664, C2V_242_677, C2V_242_845, C2V_242_887, C2V_242_950, C2V_242_981, C2V_242_1013, C2V_242_1080, C2V_242_1111, C2V_242_1393, C2V_242_1394, C2V_243_1, C2V_243_76, C2V_243_141, C2V_243_175, C2V_243_193, C2V_243_260, C2V_243_357, C2V_243_412, C2V_243_571, C2V_243_580, C2V_243_656, C2V_243_760, C2V_243_891, C2V_243_935, C2V_243_1008, C2V_243_1020, C2V_243_1098, C2V_243_1143, C2V_243_1394, C2V_243_1395, C2V_244_20, C2V_244_79, C2V_244_118, C2V_244_174, C2V_244_239, C2V_244_245, C2V_244_469, C2V_244_509, C2V_244_545, C2V_244_607, C2V_244_632, C2V_244_678, C2V_244_895, C2V_244_919, C2V_244_1003, C2V_244_1033, C2V_244_1060, C2V_244_1124, C2V_244_1395, C2V_244_1396, C2V_245_39, C2V_245_49, C2V_245_132, C2V_245_155, C2V_245_219, C2V_245_285, C2V_245_334, C2V_245_353, C2V_245_480, C2V_245_714, C2V_245_730, C2V_245_784, C2V_245_910, C2V_245_958, C2V_245_1001, C2V_245_1053, C2V_245_1102, C2V_245_1150, C2V_245_1396, C2V_245_1397, C2V_246_22, C2V_246_94, C2V_246_134, C2V_246_154, C2V_246_236, C2V_246_267, C2V_246_320, C2V_246_472, C2V_246_569, C2V_246_602, C2V_246_806, C2V_246_834, C2V_246_867, C2V_246_929, C2V_246_964, C2V_246_1031, C2V_246_1095, C2V_246_1145, C2V_246_1397, C2V_246_1398, C2V_247_46, C2V_247_82, C2V_247_102, C2V_247_163, C2V_247_225, C2V_247_268, C2V_247_368, C2V_247_422, C2V_247_519, C2V_247_755, C2V_247_803, C2V_247_851, C2V_247_892, C2V_247_933, C2V_247_967, C2V_247_1054, C2V_247_1080, C2V_247_1139, C2V_247_1398, C2V_247_1399, C2V_248_7, C2V_248_56, C2V_248_112, C2V_248_160, C2V_248_237, C2V_248_258, C2V_248_309, C2V_248_416, C2V_248_505, C2V_248_665, C2V_248_678, C2V_248_846, C2V_248_888, C2V_248_951, C2V_248_982, C2V_248_1014, C2V_248_1081, C2V_248_1112, C2V_248_1399, C2V_248_1400, C2V_249_2, C2V_249_77, C2V_249_142, C2V_249_176, C2V_249_194, C2V_249_261, C2V_249_358, C2V_249_413, C2V_249_572, C2V_249_581, C2V_249_657, C2V_249_761, C2V_249_892, C2V_249_936, C2V_249_961, C2V_249_1021, C2V_249_1099, C2V_249_1144, C2V_249_1400, C2V_249_1401, C2V_250_21, C2V_250_80, C2V_250_119, C2V_250_175, C2V_250_240, C2V_250_246, C2V_250_470, C2V_250_510, C2V_250_546, C2V_250_608, C2V_250_633, C2V_250_679, C2V_250_896, C2V_250_920, C2V_250_1004, C2V_250_1034, C2V_250_1061, C2V_250_1125, C2V_250_1401, C2V_250_1402, C2V_251_40, C2V_251_50, C2V_251_133, C2V_251_156, C2V_251_220, C2V_251_286, C2V_251_335, C2V_251_354, C2V_251_433, C2V_251_715, C2V_251_731, C2V_251_785, C2V_251_911, C2V_251_959, C2V_251_1002, C2V_251_1054, C2V_251_1103, C2V_251_1151, C2V_251_1402, C2V_251_1403, C2V_252_23, C2V_252_95, C2V_252_135, C2V_252_155, C2V_252_237, C2V_252_268, C2V_252_321, C2V_252_473, C2V_252_570, C2V_252_603, C2V_252_807, C2V_252_835, C2V_252_868, C2V_252_930, C2V_252_965, C2V_252_1032, C2V_252_1096, C2V_252_1146, C2V_252_1403, C2V_252_1404, C2V_253_47, C2V_253_83, C2V_253_103, C2V_253_164, C2V_253_226, C2V_253_269, C2V_253_369, C2V_253_423, C2V_253_520, C2V_253_756, C2V_253_804, C2V_253_852, C2V_253_893, C2V_253_934, C2V_253_968, C2V_253_1055, C2V_253_1081, C2V_253_1140, C2V_253_1404, C2V_253_1405, C2V_254_8, C2V_254_57, C2V_254_113, C2V_254_161, C2V_254_238, C2V_254_259, C2V_254_310, C2V_254_417, C2V_254_506, C2V_254_666, C2V_254_679, C2V_254_847, C2V_254_889, C2V_254_952, C2V_254_983, C2V_254_1015, C2V_254_1082, C2V_254_1113, C2V_254_1405, C2V_254_1406, C2V_255_3, C2V_255_78, C2V_255_143, C2V_255_177, C2V_255_195, C2V_255_262, C2V_255_359, C2V_255_414, C2V_255_573, C2V_255_582, C2V_255_658, C2V_255_762, C2V_255_893, C2V_255_937, C2V_255_962, C2V_255_1022, C2V_255_1100, C2V_255_1145, C2V_255_1406, C2V_255_1407, C2V_256_22, C2V_256_81, C2V_256_120, C2V_256_176, C2V_256_193, C2V_256_247, C2V_256_471, C2V_256_511, C2V_256_547, C2V_256_609, C2V_256_634, C2V_256_680, C2V_256_897, C2V_256_921, C2V_256_1005, C2V_256_1035, C2V_256_1062, C2V_256_1126, C2V_256_1407, C2V_256_1408, C2V_257_41, C2V_257_51, C2V_257_134, C2V_257_157, C2V_257_221, C2V_257_287, C2V_257_336, C2V_257_355, C2V_257_434, C2V_257_716, C2V_257_732, C2V_257_786, C2V_257_912, C2V_257_960, C2V_257_1003, C2V_257_1055, C2V_257_1104, C2V_257_1152, C2V_257_1408, C2V_257_1409, C2V_258_24, C2V_258_96, C2V_258_136, C2V_258_156, C2V_258_238, C2V_258_269, C2V_258_322, C2V_258_474, C2V_258_571, C2V_258_604, C2V_258_808, C2V_258_836, C2V_258_869, C2V_258_931, C2V_258_966, C2V_258_1033, C2V_258_1097, C2V_258_1147, C2V_258_1409, C2V_258_1410, C2V_259_48, C2V_259_84, C2V_259_104, C2V_259_165, C2V_259_227, C2V_259_270, C2V_259_370, C2V_259_424, C2V_259_521, C2V_259_757, C2V_259_805, C2V_259_853, C2V_259_894, C2V_259_935, C2V_259_969, C2V_259_1056, C2V_259_1082, C2V_259_1141, C2V_259_1410, C2V_259_1411, C2V_260_9, C2V_260_58, C2V_260_114, C2V_260_162, C2V_260_239, C2V_260_260, C2V_260_311, C2V_260_418, C2V_260_507, C2V_260_667, C2V_260_680, C2V_260_848, C2V_260_890, C2V_260_953, C2V_260_984, C2V_260_1016, C2V_260_1083, C2V_260_1114, C2V_260_1411, C2V_260_1412, C2V_261_4, C2V_261_79, C2V_261_144, C2V_261_178, C2V_261_196, C2V_261_263, C2V_261_360, C2V_261_415, C2V_261_574, C2V_261_583, C2V_261_659, C2V_261_763, C2V_261_894, C2V_261_938, C2V_261_963, C2V_261_1023, C2V_261_1101, C2V_261_1146, C2V_261_1412, C2V_261_1413, C2V_262_23, C2V_262_82, C2V_262_121, C2V_262_177, C2V_262_194, C2V_262_248, C2V_262_472, C2V_262_512, C2V_262_548, C2V_262_610, C2V_262_635, C2V_262_681, C2V_262_898, C2V_262_922, C2V_262_1006, C2V_262_1036, C2V_262_1063, C2V_262_1127, C2V_262_1413, C2V_262_1414, C2V_263_42, C2V_263_52, C2V_263_135, C2V_263_158, C2V_263_222, C2V_263_288, C2V_263_289, C2V_263_356, C2V_263_435, C2V_263_717, C2V_263_733, C2V_263_787, C2V_263_865, C2V_263_913, C2V_263_1004, C2V_263_1056, C2V_263_1057, C2V_263_1105, C2V_263_1414, C2V_263_1415, C2V_264_25, C2V_264_49, C2V_264_137, C2V_264_157, C2V_264_239, C2V_264_270, C2V_264_323, C2V_264_475, C2V_264_572, C2V_264_605, C2V_264_809, C2V_264_837, C2V_264_870, C2V_264_932, C2V_264_967, C2V_264_1034, C2V_264_1098, C2V_264_1148, C2V_264_1415, C2V_264_1416, C2V_265_1, C2V_265_85, C2V_265_105, C2V_265_166, C2V_265_228, C2V_265_271, C2V_265_371, C2V_265_425, C2V_265_522, C2V_265_758, C2V_265_806, C2V_265_854, C2V_265_895, C2V_265_936, C2V_265_970, C2V_265_1009, C2V_265_1083, C2V_265_1142, C2V_265_1416, C2V_265_1417, C2V_266_10, C2V_266_59, C2V_266_115, C2V_266_163, C2V_266_240, C2V_266_261, C2V_266_312, C2V_266_419, C2V_266_508, C2V_266_668, C2V_266_681, C2V_266_849, C2V_266_891, C2V_266_954, C2V_266_985, C2V_266_1017, C2V_266_1084, C2V_266_1115, C2V_266_1417, C2V_266_1418, C2V_267_5, C2V_267_80, C2V_267_97, C2V_267_179, C2V_267_197, C2V_267_264, C2V_267_361, C2V_267_416, C2V_267_575, C2V_267_584, C2V_267_660, C2V_267_764, C2V_267_895, C2V_267_939, C2V_267_964, C2V_267_1024, C2V_267_1102, C2V_267_1147, C2V_267_1418, C2V_267_1419, C2V_268_24, C2V_268_83, C2V_268_122, C2V_268_178, C2V_268_195, C2V_268_249, C2V_268_473, C2V_268_513, C2V_268_549, C2V_268_611, C2V_268_636, C2V_268_682, C2V_268_899, C2V_268_923, C2V_268_1007, C2V_268_1037, C2V_268_1064, C2V_268_1128, C2V_268_1419, C2V_268_1420, C2V_269_43, C2V_269_53, C2V_269_136, C2V_269_159, C2V_269_223, C2V_269_241, C2V_269_290, C2V_269_357, C2V_269_436, C2V_269_718, C2V_269_734, C2V_269_788, C2V_269_866, C2V_269_914, C2V_269_1005, C2V_269_1009, C2V_269_1058, C2V_269_1106, C2V_269_1420, C2V_269_1421, C2V_270_26, C2V_270_50, C2V_270_138, C2V_270_158, C2V_270_240, C2V_270_271, C2V_270_324, C2V_270_476, C2V_270_573, C2V_270_606, C2V_270_810, C2V_270_838, C2V_270_871, C2V_270_933, C2V_270_968, C2V_270_1035, C2V_270_1099, C2V_270_1149, C2V_270_1421, C2V_270_1422, C2V_271_2, C2V_271_86, C2V_271_106, C2V_271_167, C2V_271_229, C2V_271_272, C2V_271_372, C2V_271_426, C2V_271_523, C2V_271_759, C2V_271_807, C2V_271_855, C2V_271_896, C2V_271_937, C2V_271_971, C2V_271_1010, C2V_271_1084, C2V_271_1143, C2V_271_1422, C2V_271_1423, C2V_272_11, C2V_272_60, C2V_272_116, C2V_272_164, C2V_272_193, C2V_272_262, C2V_272_313, C2V_272_420, C2V_272_509, C2V_272_669, C2V_272_682, C2V_272_850, C2V_272_892, C2V_272_955, C2V_272_986, C2V_272_1018, C2V_272_1085, C2V_272_1116, C2V_272_1423, C2V_272_1424, C2V_273_6, C2V_273_81, C2V_273_98, C2V_273_180, C2V_273_198, C2V_273_265, C2V_273_362, C2V_273_417, C2V_273_576, C2V_273_585, C2V_273_661, C2V_273_765, C2V_273_896, C2V_273_940, C2V_273_965, C2V_273_1025, C2V_273_1103, C2V_273_1148, C2V_273_1424, C2V_273_1425, C2V_274_25, C2V_274_84, C2V_274_123, C2V_274_179, C2V_274_196, C2V_274_250, C2V_274_474, C2V_274_514, C2V_274_550, C2V_274_612, C2V_274_637, C2V_274_683, C2V_274_900, C2V_274_924, C2V_274_1008, C2V_274_1038, C2V_274_1065, C2V_274_1129, C2V_274_1425, C2V_274_1426, C2V_275_44, C2V_275_54, C2V_275_137, C2V_275_160, C2V_275_224, C2V_275_242, C2V_275_291, C2V_275_358, C2V_275_437, C2V_275_719, C2V_275_735, C2V_275_789, C2V_275_867, C2V_275_915, C2V_275_1006, C2V_275_1010, C2V_275_1059, C2V_275_1107, C2V_275_1426, C2V_275_1427, C2V_276_27, C2V_276_51, C2V_276_139, C2V_276_159, C2V_276_193, C2V_276_272, C2V_276_325, C2V_276_477, C2V_276_574, C2V_276_607, C2V_276_811, C2V_276_839, C2V_276_872, C2V_276_934, C2V_276_969, C2V_276_1036, C2V_276_1100, C2V_276_1150, C2V_276_1427, C2V_276_1428, C2V_277_3, C2V_277_87, C2V_277_107, C2V_277_168, C2V_277_230, C2V_277_273, C2V_277_373, C2V_277_427, C2V_277_524, C2V_277_760, C2V_277_808, C2V_277_856, C2V_277_897, C2V_277_938, C2V_277_972, C2V_277_1011, C2V_277_1085, C2V_277_1144, C2V_277_1428, C2V_277_1429, C2V_278_12, C2V_278_61, C2V_278_117, C2V_278_165, C2V_278_194, C2V_278_263, C2V_278_314, C2V_278_421, C2V_278_510, C2V_278_670, C2V_278_683, C2V_278_851, C2V_278_893, C2V_278_956, C2V_278_987, C2V_278_1019, C2V_278_1086, C2V_278_1117, C2V_278_1429, C2V_278_1430, C2V_279_7, C2V_279_82, C2V_279_99, C2V_279_181, C2V_279_199, C2V_279_266, C2V_279_363, C2V_279_418, C2V_279_529, C2V_279_586, C2V_279_662, C2V_279_766, C2V_279_897, C2V_279_941, C2V_279_966, C2V_279_1026, C2V_279_1104, C2V_279_1149, C2V_279_1430, C2V_279_1431, C2V_280_26, C2V_280_85, C2V_280_124, C2V_280_180, C2V_280_197, C2V_280_251, C2V_280_475, C2V_280_515, C2V_280_551, C2V_280_613, C2V_280_638, C2V_280_684, C2V_280_901, C2V_280_925, C2V_280_961, C2V_280_1039, C2V_280_1066, C2V_280_1130, C2V_280_1431, C2V_280_1432, C2V_281_45, C2V_281_55, C2V_281_138, C2V_281_161, C2V_281_225, C2V_281_243, C2V_281_292, C2V_281_359, C2V_281_438, C2V_281_720, C2V_281_736, C2V_281_790, C2V_281_868, C2V_281_916, C2V_281_1007, C2V_281_1011, C2V_281_1060, C2V_281_1108, C2V_281_1432, C2V_281_1433, C2V_282_28, C2V_282_52, C2V_282_140, C2V_282_160, C2V_282_194, C2V_282_273, C2V_282_326, C2V_282_478, C2V_282_575, C2V_282_608, C2V_282_812, C2V_282_840, C2V_282_873, C2V_282_935, C2V_282_970, C2V_282_1037, C2V_282_1101, C2V_282_1151, C2V_282_1433, C2V_282_1434, C2V_283_4, C2V_283_88, C2V_283_108, C2V_283_169, C2V_283_231, C2V_283_274, C2V_283_374, C2V_283_428, C2V_283_525, C2V_283_761, C2V_283_809, C2V_283_857, C2V_283_898, C2V_283_939, C2V_283_973, C2V_283_1012, C2V_283_1086, C2V_283_1145, C2V_283_1434, C2V_283_1435, C2V_284_13, C2V_284_62, C2V_284_118, C2V_284_166, C2V_284_195, C2V_284_264, C2V_284_315, C2V_284_422, C2V_284_511, C2V_284_671, C2V_284_684, C2V_284_852, C2V_284_894, C2V_284_957, C2V_284_988, C2V_284_1020, C2V_284_1087, C2V_284_1118, C2V_284_1435, C2V_284_1436, C2V_285_8, C2V_285_83, C2V_285_100, C2V_285_182, C2V_285_200, C2V_285_267, C2V_285_364, C2V_285_419, C2V_285_530, C2V_285_587, C2V_285_663, C2V_285_767, C2V_285_898, C2V_285_942, C2V_285_967, C2V_285_1027, C2V_285_1057, C2V_285_1150, C2V_285_1436, C2V_285_1437, C2V_286_27, C2V_286_86, C2V_286_125, C2V_286_181, C2V_286_198, C2V_286_252, C2V_286_476, C2V_286_516, C2V_286_552, C2V_286_614, C2V_286_639, C2V_286_685, C2V_286_902, C2V_286_926, C2V_286_962, C2V_286_1040, C2V_286_1067, C2V_286_1131, C2V_286_1437, C2V_286_1438, C2V_287_46, C2V_287_56, C2V_287_139, C2V_287_162, C2V_287_226, C2V_287_244, C2V_287_293, C2V_287_360, C2V_287_439, C2V_287_673, C2V_287_737, C2V_287_791, C2V_287_869, C2V_287_917, C2V_287_1008, C2V_287_1012, C2V_287_1061, C2V_287_1109, C2V_287_1438, C2V_287_1439, C2V_288_29, C2V_288_53, C2V_288_141, C2V_288_161, C2V_288_195, C2V_288_274, C2V_288_327, C2V_288_479, C2V_288_576, C2V_288_609, C2V_288_813, C2V_288_841, C2V_288_874, C2V_288_936, C2V_288_971, C2V_288_1038, C2V_288_1102, C2V_288_1152, C2V_288_1439, C2V_288_1440, C2V_0_0;
wire [quan_width - 1:0] V2C_5_1, V2C_89_1, V2C_109_1, V2C_170_1, V2C_232_1, V2C_275_1, V2C_375_1, V2C_429_1, V2C_526_1, V2C_762_1, V2C_810_1, V2C_858_1, V2C_899_1, V2C_940_1, V2C_974_1, V2C_1013_1, V2C_1087_1, V2C_1146_1, V2C_1153_1, V2C_14_2, V2C_63_2, V2C_119_2, V2C_167_2, V2C_196_2, V2C_265_2, V2C_316_2, V2C_423_2, V2C_512_2, V2C_672_2, V2C_685_2, V2C_853_2, V2C_895_2, V2C_958_2, V2C_989_2, V2C_1021_2, V2C_1088_2, V2C_1119_2, V2C_1153_2, V2C_1154_2, V2C_9_3, V2C_84_3, V2C_101_3, V2C_183_3, V2C_201_3, V2C_268_3, V2C_365_3, V2C_420_3, V2C_531_3, V2C_588_3, V2C_664_3, V2C_768_3, V2C_899_3, V2C_943_3, V2C_968_3, V2C_1028_3, V2C_1058_3, V2C_1151_3, V2C_1154_3, V2C_1155_3, V2C_28_4, V2C_87_4, V2C_126_4, V2C_182_4, V2C_199_4, V2C_253_4, V2C_477_4, V2C_517_4, V2C_553_4, V2C_615_4, V2C_640_4, V2C_686_4, V2C_903_4, V2C_927_4, V2C_963_4, V2C_1041_4, V2C_1068_4, V2C_1132_4, V2C_1155_4, V2C_1156_4, V2C_47_5, V2C_57_5, V2C_140_5, V2C_163_5, V2C_227_5, V2C_245_5, V2C_294_5, V2C_361_5, V2C_440_5, V2C_674_5, V2C_738_5, V2C_792_5, V2C_870_5, V2C_918_5, V2C_961_5, V2C_1013_5, V2C_1062_5, V2C_1110_5, V2C_1156_5, V2C_1157_5, V2C_30_6, V2C_54_6, V2C_142_6, V2C_162_6, V2C_196_6, V2C_275_6, V2C_328_6, V2C_480_6, V2C_529_6, V2C_610_6, V2C_814_6, V2C_842_6, V2C_875_6, V2C_937_6, V2C_972_6, V2C_1039_6, V2C_1103_6, V2C_1105_6, V2C_1157_6, V2C_1158_6, V2C_6_7, V2C_90_7, V2C_110_7, V2C_171_7, V2C_233_7, V2C_276_7, V2C_376_7, V2C_430_7, V2C_527_7, V2C_763_7, V2C_811_7, V2C_859_7, V2C_900_7, V2C_941_7, V2C_975_7, V2C_1014_7, V2C_1088_7, V2C_1147_7, V2C_1158_7, V2C_1159_7, V2C_15_8, V2C_64_8, V2C_120_8, V2C_168_8, V2C_197_8, V2C_266_8, V2C_317_8, V2C_424_8, V2C_513_8, V2C_625_8, V2C_686_8, V2C_854_8, V2C_896_8, V2C_959_8, V2C_990_8, V2C_1022_8, V2C_1089_8, V2C_1120_8, V2C_1159_8, V2C_1160_8, V2C_10_9, V2C_85_9, V2C_102_9, V2C_184_9, V2C_202_9, V2C_269_9, V2C_366_9, V2C_421_9, V2C_532_9, V2C_589_9, V2C_665_9, V2C_721_9, V2C_900_9, V2C_944_9, V2C_969_9, V2C_1029_9, V2C_1059_9, V2C_1152_9, V2C_1160_9, V2C_1161_9, V2C_29_10, V2C_88_10, V2C_127_10, V2C_183_10, V2C_200_10, V2C_254_10, V2C_478_10, V2C_518_10, V2C_554_10, V2C_616_10, V2C_641_10, V2C_687_10, V2C_904_10, V2C_928_10, V2C_964_10, V2C_1042_10, V2C_1069_10, V2C_1133_10, V2C_1161_10, V2C_1162_10, V2C_48_11, V2C_58_11, V2C_141_11, V2C_164_11, V2C_228_11, V2C_246_11, V2C_295_11, V2C_362_11, V2C_441_11, V2C_675_11, V2C_739_11, V2C_793_11, V2C_871_11, V2C_919_11, V2C_962_11, V2C_1014_11, V2C_1063_11, V2C_1111_11, V2C_1162_11, V2C_1163_11, V2C_31_12, V2C_55_12, V2C_143_12, V2C_163_12, V2C_197_12, V2C_276_12, V2C_329_12, V2C_433_12, V2C_530_12, V2C_611_12, V2C_815_12, V2C_843_12, V2C_876_12, V2C_938_12, V2C_973_12, V2C_1040_12, V2C_1104_12, V2C_1106_12, V2C_1163_12, V2C_1164_12, V2C_7_13, V2C_91_13, V2C_111_13, V2C_172_13, V2C_234_13, V2C_277_13, V2C_377_13, V2C_431_13, V2C_528_13, V2C_764_13, V2C_812_13, V2C_860_13, V2C_901_13, V2C_942_13, V2C_976_13, V2C_1015_13, V2C_1089_13, V2C_1148_13, V2C_1164_13, V2C_1165_13, V2C_16_14, V2C_65_14, V2C_121_14, V2C_169_14, V2C_198_14, V2C_267_14, V2C_318_14, V2C_425_14, V2C_514_14, V2C_626_14, V2C_687_14, V2C_855_14, V2C_897_14, V2C_960_14, V2C_991_14, V2C_1023_14, V2C_1090_14, V2C_1121_14, V2C_1165_14, V2C_1166_14, V2C_11_15, V2C_86_15, V2C_103_15, V2C_185_15, V2C_203_15, V2C_270_15, V2C_367_15, V2C_422_15, V2C_533_15, V2C_590_15, V2C_666_15, V2C_722_15, V2C_901_15, V2C_945_15, V2C_970_15, V2C_1030_15, V2C_1060_15, V2C_1105_15, V2C_1166_15, V2C_1167_15, V2C_30_16, V2C_89_16, V2C_128_16, V2C_184_16, V2C_201_16, V2C_255_16, V2C_479_16, V2C_519_16, V2C_555_16, V2C_617_16, V2C_642_16, V2C_688_16, V2C_905_16, V2C_929_16, V2C_965_16, V2C_1043_16, V2C_1070_16, V2C_1134_16, V2C_1167_16, V2C_1168_16, V2C_1_17, V2C_59_17, V2C_142_17, V2C_165_17, V2C_229_17, V2C_247_17, V2C_296_17, V2C_363_17, V2C_442_17, V2C_676_17, V2C_740_17, V2C_794_17, V2C_872_17, V2C_920_17, V2C_963_17, V2C_1015_17, V2C_1064_17, V2C_1112_17, V2C_1168_17, V2C_1169_17, V2C_32_18, V2C_56_18, V2C_144_18, V2C_164_18, V2C_198_18, V2C_277_18, V2C_330_18, V2C_434_18, V2C_531_18, V2C_612_18, V2C_816_18, V2C_844_18, V2C_877_18, V2C_939_18, V2C_974_18, V2C_1041_18, V2C_1057_18, V2C_1107_18, V2C_1169_18, V2C_1170_18, V2C_8_19, V2C_92_19, V2C_112_19, V2C_173_19, V2C_235_19, V2C_278_19, V2C_378_19, V2C_432_19, V2C_481_19, V2C_765_19, V2C_813_19, V2C_861_19, V2C_902_19, V2C_943_19, V2C_977_19, V2C_1016_19, V2C_1090_19, V2C_1149_19, V2C_1170_19, V2C_1171_19, V2C_17_20, V2C_66_20, V2C_122_20, V2C_170_20, V2C_199_20, V2C_268_20, V2C_319_20, V2C_426_20, V2C_515_20, V2C_627_20, V2C_688_20, V2C_856_20, V2C_898_20, V2C_913_20, V2C_992_20, V2C_1024_20, V2C_1091_20, V2C_1122_20, V2C_1171_20, V2C_1172_20, V2C_12_21, V2C_87_21, V2C_104_21, V2C_186_21, V2C_204_21, V2C_271_21, V2C_368_21, V2C_423_21, V2C_534_21, V2C_591_21, V2C_667_21, V2C_723_21, V2C_902_21, V2C_946_21, V2C_971_21, V2C_1031_21, V2C_1061_21, V2C_1106_21, V2C_1172_21, V2C_1173_21, V2C_31_22, V2C_90_22, V2C_129_22, V2C_185_22, V2C_202_22, V2C_256_22, V2C_480_22, V2C_520_22, V2C_556_22, V2C_618_22, V2C_643_22, V2C_689_22, V2C_906_22, V2C_930_22, V2C_966_22, V2C_1044_22, V2C_1071_22, V2C_1135_22, V2C_1173_22, V2C_1174_22, V2C_2_23, V2C_60_23, V2C_143_23, V2C_166_23, V2C_230_23, V2C_248_23, V2C_297_23, V2C_364_23, V2C_443_23, V2C_677_23, V2C_741_23, V2C_795_23, V2C_873_23, V2C_921_23, V2C_964_23, V2C_1016_23, V2C_1065_23, V2C_1113_23, V2C_1174_23, V2C_1175_23, V2C_33_24, V2C_57_24, V2C_97_24, V2C_165_24, V2C_199_24, V2C_278_24, V2C_331_24, V2C_435_24, V2C_532_24, V2C_613_24, V2C_769_24, V2C_845_24, V2C_878_24, V2C_940_24, V2C_975_24, V2C_1042_24, V2C_1058_24, V2C_1108_24, V2C_1175_24, V2C_1176_24, V2C_9_25, V2C_93_25, V2C_113_25, V2C_174_25, V2C_236_25, V2C_279_25, V2C_379_25, V2C_385_25, V2C_482_25, V2C_766_25, V2C_814_25, V2C_862_25, V2C_903_25, V2C_944_25, V2C_978_25, V2C_1017_25, V2C_1091_25, V2C_1150_25, V2C_1176_25, V2C_1177_25, V2C_18_26, V2C_67_26, V2C_123_26, V2C_171_26, V2C_200_26, V2C_269_26, V2C_320_26, V2C_427_26, V2C_516_26, V2C_628_26, V2C_689_26, V2C_857_26, V2C_899_26, V2C_914_26, V2C_993_26, V2C_1025_26, V2C_1092_26, V2C_1123_26, V2C_1177_26, V2C_1178_26, V2C_13_27, V2C_88_27, V2C_105_27, V2C_187_27, V2C_205_27, V2C_272_27, V2C_369_27, V2C_424_27, V2C_535_27, V2C_592_27, V2C_668_27, V2C_724_27, V2C_903_27, V2C_947_27, V2C_972_27, V2C_1032_27, V2C_1062_27, V2C_1107_27, V2C_1178_27, V2C_1179_27, V2C_32_28, V2C_91_28, V2C_130_28, V2C_186_28, V2C_203_28, V2C_257_28, V2C_433_28, V2C_521_28, V2C_557_28, V2C_619_28, V2C_644_28, V2C_690_28, V2C_907_28, V2C_931_28, V2C_967_28, V2C_1045_28, V2C_1072_28, V2C_1136_28, V2C_1179_28, V2C_1180_28, V2C_3_29, V2C_61_29, V2C_144_29, V2C_167_29, V2C_231_29, V2C_249_29, V2C_298_29, V2C_365_29, V2C_444_29, V2C_678_29, V2C_742_29, V2C_796_29, V2C_874_29, V2C_922_29, V2C_965_29, V2C_1017_29, V2C_1066_29, V2C_1114_29, V2C_1180_29, V2C_1181_29, V2C_34_30, V2C_58_30, V2C_98_30, V2C_166_30, V2C_200_30, V2C_279_30, V2C_332_30, V2C_436_30, V2C_533_30, V2C_614_30, V2C_770_30, V2C_846_30, V2C_879_30, V2C_941_30, V2C_976_30, V2C_1043_30, V2C_1059_30, V2C_1109_30, V2C_1181_30, V2C_1182_30, V2C_10_31, V2C_94_31, V2C_114_31, V2C_175_31, V2C_237_31, V2C_280_31, V2C_380_31, V2C_386_31, V2C_483_31, V2C_767_31, V2C_815_31, V2C_863_31, V2C_904_31, V2C_945_31, V2C_979_31, V2C_1018_31, V2C_1092_31, V2C_1151_31, V2C_1182_31, V2C_1183_31, V2C_19_32, V2C_68_32, V2C_124_32, V2C_172_32, V2C_201_32, V2C_270_32, V2C_321_32, V2C_428_32, V2C_517_32, V2C_629_32, V2C_690_32, V2C_858_32, V2C_900_32, V2C_915_32, V2C_994_32, V2C_1026_32, V2C_1093_32, V2C_1124_32, V2C_1183_32, V2C_1184_32, V2C_14_33, V2C_89_33, V2C_106_33, V2C_188_33, V2C_206_33, V2C_273_33, V2C_370_33, V2C_425_33, V2C_536_33, V2C_593_33, V2C_669_33, V2C_725_33, V2C_904_33, V2C_948_33, V2C_973_33, V2C_1033_33, V2C_1063_33, V2C_1108_33, V2C_1184_33, V2C_1185_33, V2C_33_34, V2C_92_34, V2C_131_34, V2C_187_34, V2C_204_34, V2C_258_34, V2C_434_34, V2C_522_34, V2C_558_34, V2C_620_34, V2C_645_34, V2C_691_34, V2C_908_34, V2C_932_34, V2C_968_34, V2C_1046_34, V2C_1073_34, V2C_1137_34, V2C_1185_34, V2C_1186_34, V2C_4_35, V2C_62_35, V2C_97_35, V2C_168_35, V2C_232_35, V2C_250_35, V2C_299_35, V2C_366_35, V2C_445_35, V2C_679_35, V2C_743_35, V2C_797_35, V2C_875_35, V2C_923_35, V2C_966_35, V2C_1018_35, V2C_1067_35, V2C_1115_35, V2C_1186_35, V2C_1187_35, V2C_35_36, V2C_59_36, V2C_99_36, V2C_167_36, V2C_201_36, V2C_280_36, V2C_333_36, V2C_437_36, V2C_534_36, V2C_615_36, V2C_771_36, V2C_847_36, V2C_880_36, V2C_942_36, V2C_977_36, V2C_1044_36, V2C_1060_36, V2C_1110_36, V2C_1187_36, V2C_1188_36, V2C_11_37, V2C_95_37, V2C_115_37, V2C_176_37, V2C_238_37, V2C_281_37, V2C_381_37, V2C_387_37, V2C_484_37, V2C_768_37, V2C_816_37, V2C_864_37, V2C_905_37, V2C_946_37, V2C_980_37, V2C_1019_37, V2C_1093_37, V2C_1152_37, V2C_1188_37, V2C_1189_37, V2C_20_38, V2C_69_38, V2C_125_38, V2C_173_38, V2C_202_38, V2C_271_38, V2C_322_38, V2C_429_38, V2C_518_38, V2C_630_38, V2C_691_38, V2C_859_38, V2C_901_38, V2C_916_38, V2C_995_38, V2C_1027_38, V2C_1094_38, V2C_1125_38, V2C_1189_38, V2C_1190_38, V2C_15_39, V2C_90_39, V2C_107_39, V2C_189_39, V2C_207_39, V2C_274_39, V2C_371_39, V2C_426_39, V2C_537_39, V2C_594_39, V2C_670_39, V2C_726_39, V2C_905_39, V2C_949_39, V2C_974_39, V2C_1034_39, V2C_1064_39, V2C_1109_39, V2C_1190_39, V2C_1191_39, V2C_34_40, V2C_93_40, V2C_132_40, V2C_188_40, V2C_205_40, V2C_259_40, V2C_435_40, V2C_523_40, V2C_559_40, V2C_621_40, V2C_646_40, V2C_692_40, V2C_909_40, V2C_933_40, V2C_969_40, V2C_1047_40, V2C_1074_40, V2C_1138_40, V2C_1191_40, V2C_1192_40, V2C_5_41, V2C_63_41, V2C_98_41, V2C_169_41, V2C_233_41, V2C_251_41, V2C_300_41, V2C_367_41, V2C_446_41, V2C_680_41, V2C_744_41, V2C_798_41, V2C_876_41, V2C_924_41, V2C_967_41, V2C_1019_41, V2C_1068_41, V2C_1116_41, V2C_1192_41, V2C_1193_41, V2C_36_42, V2C_60_42, V2C_100_42, V2C_168_42, V2C_202_42, V2C_281_42, V2C_334_42, V2C_438_42, V2C_535_42, V2C_616_42, V2C_772_42, V2C_848_42, V2C_881_42, V2C_943_42, V2C_978_42, V2C_1045_42, V2C_1061_42, V2C_1111_42, V2C_1193_42, V2C_1194_42, V2C_12_43, V2C_96_43, V2C_116_43, V2C_177_43, V2C_239_43, V2C_282_43, V2C_382_43, V2C_388_43, V2C_485_43, V2C_721_43, V2C_769_43, V2C_817_43, V2C_906_43, V2C_947_43, V2C_981_43, V2C_1020_43, V2C_1094_43, V2C_1105_43, V2C_1194_43, V2C_1195_43, V2C_21_44, V2C_70_44, V2C_126_44, V2C_174_44, V2C_203_44, V2C_272_44, V2C_323_44, V2C_430_44, V2C_519_44, V2C_631_44, V2C_692_44, V2C_860_44, V2C_902_44, V2C_917_44, V2C_996_44, V2C_1028_44, V2C_1095_44, V2C_1126_44, V2C_1195_44, V2C_1196_44, V2C_16_45, V2C_91_45, V2C_108_45, V2C_190_45, V2C_208_45, V2C_275_45, V2C_372_45, V2C_427_45, V2C_538_45, V2C_595_45, V2C_671_45, V2C_727_45, V2C_906_45, V2C_950_45, V2C_975_45, V2C_1035_45, V2C_1065_45, V2C_1110_45, V2C_1196_45, V2C_1197_45, V2C_35_46, V2C_94_46, V2C_133_46, V2C_189_46, V2C_206_46, V2C_260_46, V2C_436_46, V2C_524_46, V2C_560_46, V2C_622_46, V2C_647_46, V2C_693_46, V2C_910_46, V2C_934_46, V2C_970_46, V2C_1048_46, V2C_1075_46, V2C_1139_46, V2C_1197_46, V2C_1198_46, V2C_6_47, V2C_64_47, V2C_99_47, V2C_170_47, V2C_234_47, V2C_252_47, V2C_301_47, V2C_368_47, V2C_447_47, V2C_681_47, V2C_745_47, V2C_799_47, V2C_877_47, V2C_925_47, V2C_968_47, V2C_1020_47, V2C_1069_47, V2C_1117_47, V2C_1198_47, V2C_1199_47, V2C_37_48, V2C_61_48, V2C_101_48, V2C_169_48, V2C_203_48, V2C_282_48, V2C_335_48, V2C_439_48, V2C_536_48, V2C_617_48, V2C_773_48, V2C_849_48, V2C_882_48, V2C_944_48, V2C_979_48, V2C_1046_48, V2C_1062_48, V2C_1112_48, V2C_1199_48, V2C_1200_48, V2C_13_49, V2C_49_49, V2C_117_49, V2C_178_49, V2C_240_49, V2C_283_49, V2C_383_49, V2C_389_49, V2C_486_49, V2C_722_49, V2C_770_49, V2C_818_49, V2C_907_49, V2C_948_49, V2C_982_49, V2C_1021_49, V2C_1095_49, V2C_1106_49, V2C_1200_49, V2C_1201_49, V2C_22_50, V2C_71_50, V2C_127_50, V2C_175_50, V2C_204_50, V2C_273_50, V2C_324_50, V2C_431_50, V2C_520_50, V2C_632_50, V2C_693_50, V2C_861_50, V2C_903_50, V2C_918_50, V2C_997_50, V2C_1029_50, V2C_1096_50, V2C_1127_50, V2C_1201_50, V2C_1202_50, V2C_17_51, V2C_92_51, V2C_109_51, V2C_191_51, V2C_209_51, V2C_276_51, V2C_373_51, V2C_428_51, V2C_539_51, V2C_596_51, V2C_672_51, V2C_728_51, V2C_907_51, V2C_951_51, V2C_976_51, V2C_1036_51, V2C_1066_51, V2C_1111_51, V2C_1202_51, V2C_1203_51, V2C_36_52, V2C_95_52, V2C_134_52, V2C_190_52, V2C_207_52, V2C_261_52, V2C_437_52, V2C_525_52, V2C_561_52, V2C_623_52, V2C_648_52, V2C_694_52, V2C_911_52, V2C_935_52, V2C_971_52, V2C_1049_52, V2C_1076_52, V2C_1140_52, V2C_1203_52, V2C_1204_52, V2C_7_53, V2C_65_53, V2C_100_53, V2C_171_53, V2C_235_53, V2C_253_53, V2C_302_53, V2C_369_53, V2C_448_53, V2C_682_53, V2C_746_53, V2C_800_53, V2C_878_53, V2C_926_53, V2C_969_53, V2C_1021_53, V2C_1070_53, V2C_1118_53, V2C_1204_53, V2C_1205_53, V2C_38_54, V2C_62_54, V2C_102_54, V2C_170_54, V2C_204_54, V2C_283_54, V2C_336_54, V2C_440_54, V2C_537_54, V2C_618_54, V2C_774_54, V2C_850_54, V2C_883_54, V2C_945_54, V2C_980_54, V2C_1047_54, V2C_1063_54, V2C_1113_54, V2C_1205_54, V2C_1206_54, V2C_14_55, V2C_50_55, V2C_118_55, V2C_179_55, V2C_193_55, V2C_284_55, V2C_384_55, V2C_390_55, V2C_487_55, V2C_723_55, V2C_771_55, V2C_819_55, V2C_908_55, V2C_949_55, V2C_983_55, V2C_1022_55, V2C_1096_55, V2C_1107_55, V2C_1206_55, V2C_1207_55, V2C_23_56, V2C_72_56, V2C_128_56, V2C_176_56, V2C_205_56, V2C_274_56, V2C_325_56, V2C_432_56, V2C_521_56, V2C_633_56, V2C_694_56, V2C_862_56, V2C_904_56, V2C_919_56, V2C_998_56, V2C_1030_56, V2C_1097_56, V2C_1128_56, V2C_1207_56, V2C_1208_56, V2C_18_57, V2C_93_57, V2C_110_57, V2C_192_57, V2C_210_57, V2C_277_57, V2C_374_57, V2C_429_57, V2C_540_57, V2C_597_57, V2C_625_57, V2C_729_57, V2C_908_57, V2C_952_57, V2C_977_57, V2C_1037_57, V2C_1067_57, V2C_1112_57, V2C_1208_57, V2C_1209_57, V2C_37_58, V2C_96_58, V2C_135_58, V2C_191_58, V2C_208_58, V2C_262_58, V2C_438_58, V2C_526_58, V2C_562_58, V2C_624_58, V2C_649_58, V2C_695_58, V2C_912_58, V2C_936_58, V2C_972_58, V2C_1050_58, V2C_1077_58, V2C_1141_58, V2C_1209_58, V2C_1210_58, V2C_8_59, V2C_66_59, V2C_101_59, V2C_172_59, V2C_236_59, V2C_254_59, V2C_303_59, V2C_370_59, V2C_449_59, V2C_683_59, V2C_747_59, V2C_801_59, V2C_879_59, V2C_927_59, V2C_970_59, V2C_1022_59, V2C_1071_59, V2C_1119_59, V2C_1210_59, V2C_1211_59, V2C_39_60, V2C_63_60, V2C_103_60, V2C_171_60, V2C_205_60, V2C_284_60, V2C_289_60, V2C_441_60, V2C_538_60, V2C_619_60, V2C_775_60, V2C_851_60, V2C_884_60, V2C_946_60, V2C_981_60, V2C_1048_60, V2C_1064_60, V2C_1114_60, V2C_1211_60, V2C_1212_60, V2C_15_61, V2C_51_61, V2C_119_61, V2C_180_61, V2C_194_61, V2C_285_61, V2C_337_61, V2C_391_61, V2C_488_61, V2C_724_61, V2C_772_61, V2C_820_61, V2C_909_61, V2C_950_61, V2C_984_61, V2C_1023_61, V2C_1097_61, V2C_1108_61, V2C_1212_61, V2C_1213_61, V2C_24_62, V2C_73_62, V2C_129_62, V2C_177_62, V2C_206_62, V2C_275_62, V2C_326_62, V2C_385_62, V2C_522_62, V2C_634_62, V2C_695_62, V2C_863_62, V2C_905_62, V2C_920_62, V2C_999_62, V2C_1031_62, V2C_1098_62, V2C_1129_62, V2C_1213_62, V2C_1214_62, V2C_19_63, V2C_94_63, V2C_111_63, V2C_145_63, V2C_211_63, V2C_278_63, V2C_375_63, V2C_430_63, V2C_541_63, V2C_598_63, V2C_626_63, V2C_730_63, V2C_909_63, V2C_953_63, V2C_978_63, V2C_1038_63, V2C_1068_63, V2C_1113_63, V2C_1214_63, V2C_1215_63, V2C_38_64, V2C_49_64, V2C_136_64, V2C_192_64, V2C_209_64, V2C_263_64, V2C_439_64, V2C_527_64, V2C_563_64, V2C_577_64, V2C_650_64, V2C_696_64, V2C_865_64, V2C_937_64, V2C_973_64, V2C_1051_64, V2C_1078_64, V2C_1142_64, V2C_1215_64, V2C_1216_64, V2C_9_65, V2C_67_65, V2C_102_65, V2C_173_65, V2C_237_65, V2C_255_65, V2C_304_65, V2C_371_65, V2C_450_65, V2C_684_65, V2C_748_65, V2C_802_65, V2C_880_65, V2C_928_65, V2C_971_65, V2C_1023_65, V2C_1072_65, V2C_1120_65, V2C_1216_65, V2C_1217_65, V2C_40_66, V2C_64_66, V2C_104_66, V2C_172_66, V2C_206_66, V2C_285_66, V2C_290_66, V2C_442_66, V2C_539_66, V2C_620_66, V2C_776_66, V2C_852_66, V2C_885_66, V2C_947_66, V2C_982_66, V2C_1049_66, V2C_1065_66, V2C_1115_66, V2C_1217_66, V2C_1218_66, V2C_16_67, V2C_52_67, V2C_120_67, V2C_181_67, V2C_195_67, V2C_286_67, V2C_338_67, V2C_392_67, V2C_489_67, V2C_725_67, V2C_773_67, V2C_821_67, V2C_910_67, V2C_951_67, V2C_985_67, V2C_1024_67, V2C_1098_67, V2C_1109_67, V2C_1218_67, V2C_1219_67, V2C_25_68, V2C_74_68, V2C_130_68, V2C_178_68, V2C_207_68, V2C_276_68, V2C_327_68, V2C_386_68, V2C_523_68, V2C_635_68, V2C_696_68, V2C_864_68, V2C_906_68, V2C_921_68, V2C_1000_68, V2C_1032_68, V2C_1099_68, V2C_1130_68, V2C_1219_68, V2C_1220_68, V2C_20_69, V2C_95_69, V2C_112_69, V2C_146_69, V2C_212_69, V2C_279_69, V2C_376_69, V2C_431_69, V2C_542_69, V2C_599_69, V2C_627_69, V2C_731_69, V2C_910_69, V2C_954_69, V2C_979_69, V2C_1039_69, V2C_1069_69, V2C_1114_69, V2C_1220_69, V2C_1221_69, V2C_39_70, V2C_50_70, V2C_137_70, V2C_145_70, V2C_210_70, V2C_264_70, V2C_440_70, V2C_528_70, V2C_564_70, V2C_578_70, V2C_651_70, V2C_697_70, V2C_866_70, V2C_938_70, V2C_974_70, V2C_1052_70, V2C_1079_70, V2C_1143_70, V2C_1221_70, V2C_1222_70, V2C_10_71, V2C_68_71, V2C_103_71, V2C_174_71, V2C_238_71, V2C_256_71, V2C_305_71, V2C_372_71, V2C_451_71, V2C_685_71, V2C_749_71, V2C_803_71, V2C_881_71, V2C_929_71, V2C_972_71, V2C_1024_71, V2C_1073_71, V2C_1121_71, V2C_1222_71, V2C_1223_71, V2C_41_72, V2C_65_72, V2C_105_72, V2C_173_72, V2C_207_72, V2C_286_72, V2C_291_72, V2C_443_72, V2C_540_72, V2C_621_72, V2C_777_72, V2C_853_72, V2C_886_72, V2C_948_72, V2C_983_72, V2C_1050_72, V2C_1066_72, V2C_1116_72, V2C_1223_72, V2C_1224_72, V2C_17_73, V2C_53_73, V2C_121_73, V2C_182_73, V2C_196_73, V2C_287_73, V2C_339_73, V2C_393_73, V2C_490_73, V2C_726_73, V2C_774_73, V2C_822_73, V2C_911_73, V2C_952_73, V2C_986_73, V2C_1025_73, V2C_1099_73, V2C_1110_73, V2C_1224_73, V2C_1225_73, V2C_26_74, V2C_75_74, V2C_131_74, V2C_179_74, V2C_208_74, V2C_277_74, V2C_328_74, V2C_387_74, V2C_524_74, V2C_636_74, V2C_697_74, V2C_817_74, V2C_907_74, V2C_922_74, V2C_1001_74, V2C_1033_74, V2C_1100_74, V2C_1131_74, V2C_1225_74, V2C_1226_74, V2C_21_75, V2C_96_75, V2C_113_75, V2C_147_75, V2C_213_75, V2C_280_75, V2C_377_75, V2C_432_75, V2C_543_75, V2C_600_75, V2C_628_75, V2C_732_75, V2C_911_75, V2C_955_75, V2C_980_75, V2C_1040_75, V2C_1070_75, V2C_1115_75, V2C_1226_75, V2C_1227_75, V2C_40_76, V2C_51_76, V2C_138_76, V2C_146_76, V2C_211_76, V2C_265_76, V2C_441_76, V2C_481_76, V2C_565_76, V2C_579_76, V2C_652_76, V2C_698_76, V2C_867_76, V2C_939_76, V2C_975_76, V2C_1053_76, V2C_1080_76, V2C_1144_76, V2C_1227_76, V2C_1228_76, V2C_11_77, V2C_69_77, V2C_104_77, V2C_175_77, V2C_239_77, V2C_257_77, V2C_306_77, V2C_373_77, V2C_452_77, V2C_686_77, V2C_750_77, V2C_804_77, V2C_882_77, V2C_930_77, V2C_973_77, V2C_1025_77, V2C_1074_77, V2C_1122_77, V2C_1228_77, V2C_1229_77, V2C_42_78, V2C_66_78, V2C_106_78, V2C_174_78, V2C_208_78, V2C_287_78, V2C_292_78, V2C_444_78, V2C_541_78, V2C_622_78, V2C_778_78, V2C_854_78, V2C_887_78, V2C_949_78, V2C_984_78, V2C_1051_78, V2C_1067_78, V2C_1117_78, V2C_1229_78, V2C_1230_78, V2C_18_79, V2C_54_79, V2C_122_79, V2C_183_79, V2C_197_79, V2C_288_79, V2C_340_79, V2C_394_79, V2C_491_79, V2C_727_79, V2C_775_79, V2C_823_79, V2C_912_79, V2C_953_79, V2C_987_79, V2C_1026_79, V2C_1100_79, V2C_1111_79, V2C_1230_79, V2C_1231_79, V2C_27_80, V2C_76_80, V2C_132_80, V2C_180_80, V2C_209_80, V2C_278_80, V2C_329_80, V2C_388_80, V2C_525_80, V2C_637_80, V2C_698_80, V2C_818_80, V2C_908_80, V2C_923_80, V2C_1002_80, V2C_1034_80, V2C_1101_80, V2C_1132_80, V2C_1231_80, V2C_1232_80, V2C_22_81, V2C_49_81, V2C_114_81, V2C_148_81, V2C_214_81, V2C_281_81, V2C_378_81, V2C_385_81, V2C_544_81, V2C_601_81, V2C_629_81, V2C_733_81, V2C_912_81, V2C_956_81, V2C_981_81, V2C_1041_81, V2C_1071_81, V2C_1116_81, V2C_1232_81, V2C_1233_81, V2C_41_82, V2C_52_82, V2C_139_82, V2C_147_82, V2C_212_82, V2C_266_82, V2C_442_82, V2C_482_82, V2C_566_82, V2C_580_82, V2C_653_82, V2C_699_82, V2C_868_82, V2C_940_82, V2C_976_82, V2C_1054_82, V2C_1081_82, V2C_1145_82, V2C_1233_82, V2C_1234_82, V2C_12_83, V2C_70_83, V2C_105_83, V2C_176_83, V2C_240_83, V2C_258_83, V2C_307_83, V2C_374_83, V2C_453_83, V2C_687_83, V2C_751_83, V2C_805_83, V2C_883_83, V2C_931_83, V2C_974_83, V2C_1026_83, V2C_1075_83, V2C_1123_83, V2C_1234_83, V2C_1235_83, V2C_43_84, V2C_67_84, V2C_107_84, V2C_175_84, V2C_209_84, V2C_288_84, V2C_293_84, V2C_445_84, V2C_542_84, V2C_623_84, V2C_779_84, V2C_855_84, V2C_888_84, V2C_950_84, V2C_985_84, V2C_1052_84, V2C_1068_84, V2C_1118_84, V2C_1235_84, V2C_1236_84, V2C_19_85, V2C_55_85, V2C_123_85, V2C_184_85, V2C_198_85, V2C_241_85, V2C_341_85, V2C_395_85, V2C_492_85, V2C_728_85, V2C_776_85, V2C_824_85, V2C_865_85, V2C_954_85, V2C_988_85, V2C_1027_85, V2C_1101_85, V2C_1112_85, V2C_1236_85, V2C_1237_85, V2C_28_86, V2C_77_86, V2C_133_86, V2C_181_86, V2C_210_86, V2C_279_86, V2C_330_86, V2C_389_86, V2C_526_86, V2C_638_86, V2C_699_86, V2C_819_86, V2C_909_86, V2C_924_86, V2C_1003_86, V2C_1035_86, V2C_1102_86, V2C_1133_86, V2C_1237_86, V2C_1238_86, V2C_23_87, V2C_50_87, V2C_115_87, V2C_149_87, V2C_215_87, V2C_282_87, V2C_379_87, V2C_386_87, V2C_545_87, V2C_602_87, V2C_630_87, V2C_734_87, V2C_865_87, V2C_957_87, V2C_982_87, V2C_1042_87, V2C_1072_87, V2C_1117_87, V2C_1238_87, V2C_1239_87, V2C_42_88, V2C_53_88, V2C_140_88, V2C_148_88, V2C_213_88, V2C_267_88, V2C_443_88, V2C_483_88, V2C_567_88, V2C_581_88, V2C_654_88, V2C_700_88, V2C_869_88, V2C_941_88, V2C_977_88, V2C_1055_88, V2C_1082_88, V2C_1146_88, V2C_1239_88, V2C_1240_88, V2C_13_89, V2C_71_89, V2C_106_89, V2C_177_89, V2C_193_89, V2C_259_89, V2C_308_89, V2C_375_89, V2C_454_89, V2C_688_89, V2C_752_89, V2C_806_89, V2C_884_89, V2C_932_89, V2C_975_89, V2C_1027_89, V2C_1076_89, V2C_1124_89, V2C_1240_89, V2C_1241_89, V2C_44_90, V2C_68_90, V2C_108_90, V2C_176_90, V2C_210_90, V2C_241_90, V2C_294_90, V2C_446_90, V2C_543_90, V2C_624_90, V2C_780_90, V2C_856_90, V2C_889_90, V2C_951_90, V2C_986_90, V2C_1053_90, V2C_1069_90, V2C_1119_90, V2C_1241_90, V2C_1242_90, V2C_20_91, V2C_56_91, V2C_124_91, V2C_185_91, V2C_199_91, V2C_242_91, V2C_342_91, V2C_396_91, V2C_493_91, V2C_729_91, V2C_777_91, V2C_825_91, V2C_866_91, V2C_955_91, V2C_989_91, V2C_1028_91, V2C_1102_91, V2C_1113_91, V2C_1242_91, V2C_1243_91, V2C_29_92, V2C_78_92, V2C_134_92, V2C_182_92, V2C_211_92, V2C_280_92, V2C_331_92, V2C_390_92, V2C_527_92, V2C_639_92, V2C_700_92, V2C_820_92, V2C_910_92, V2C_925_92, V2C_1004_92, V2C_1036_92, V2C_1103_92, V2C_1134_92, V2C_1243_92, V2C_1244_92, V2C_24_93, V2C_51_93, V2C_116_93, V2C_150_93, V2C_216_93, V2C_283_93, V2C_380_93, V2C_387_93, V2C_546_93, V2C_603_93, V2C_631_93, V2C_735_93, V2C_866_93, V2C_958_93, V2C_983_93, V2C_1043_93, V2C_1073_93, V2C_1118_93, V2C_1244_93, V2C_1245_93, V2C_43_94, V2C_54_94, V2C_141_94, V2C_149_94, V2C_214_94, V2C_268_94, V2C_444_94, V2C_484_94, V2C_568_94, V2C_582_94, V2C_655_94, V2C_701_94, V2C_870_94, V2C_942_94, V2C_978_94, V2C_1056_94, V2C_1083_94, V2C_1147_94, V2C_1245_94, V2C_1246_94, V2C_14_95, V2C_72_95, V2C_107_95, V2C_178_95, V2C_194_95, V2C_260_95, V2C_309_95, V2C_376_95, V2C_455_95, V2C_689_95, V2C_753_95, V2C_807_95, V2C_885_95, V2C_933_95, V2C_976_95, V2C_1028_95, V2C_1077_95, V2C_1125_95, V2C_1246_95, V2C_1247_95, V2C_45_96, V2C_69_96, V2C_109_96, V2C_177_96, V2C_211_96, V2C_242_96, V2C_295_96, V2C_447_96, V2C_544_96, V2C_577_96, V2C_781_96, V2C_857_96, V2C_890_96, V2C_952_96, V2C_987_96, V2C_1054_96, V2C_1070_96, V2C_1120_96, V2C_1247_96, V2C_1248_96, V2C_21_97, V2C_57_97, V2C_125_97, V2C_186_97, V2C_200_97, V2C_243_97, V2C_343_97, V2C_397_97, V2C_494_97, V2C_730_97, V2C_778_97, V2C_826_97, V2C_867_97, V2C_956_97, V2C_990_97, V2C_1029_97, V2C_1103_97, V2C_1114_97, V2C_1248_97, V2C_1249_97, V2C_30_98, V2C_79_98, V2C_135_98, V2C_183_98, V2C_212_98, V2C_281_98, V2C_332_98, V2C_391_98, V2C_528_98, V2C_640_98, V2C_701_98, V2C_821_98, V2C_911_98, V2C_926_98, V2C_1005_98, V2C_1037_98, V2C_1104_98, V2C_1135_98, V2C_1249_98, V2C_1250_98, V2C_25_99, V2C_52_99, V2C_117_99, V2C_151_99, V2C_217_99, V2C_284_99, V2C_381_99, V2C_388_99, V2C_547_99, V2C_604_99, V2C_632_99, V2C_736_99, V2C_867_99, V2C_959_99, V2C_984_99, V2C_1044_99, V2C_1074_99, V2C_1119_99, V2C_1250_99, V2C_1251_99, V2C_44_100, V2C_55_100, V2C_142_100, V2C_150_100, V2C_215_100, V2C_269_100, V2C_445_100, V2C_485_100, V2C_569_100, V2C_583_100, V2C_656_100, V2C_702_100, V2C_871_100, V2C_943_100, V2C_979_100, V2C_1009_100, V2C_1084_100, V2C_1148_100, V2C_1251_100, V2C_1252_100, V2C_15_101, V2C_73_101, V2C_108_101, V2C_179_101, V2C_195_101, V2C_261_101, V2C_310_101, V2C_377_101, V2C_456_101, V2C_690_101, V2C_754_101, V2C_808_101, V2C_886_101, V2C_934_101, V2C_977_101, V2C_1029_101, V2C_1078_101, V2C_1126_101, V2C_1252_101, V2C_1253_101, V2C_46_102, V2C_70_102, V2C_110_102, V2C_178_102, V2C_212_102, V2C_243_102, V2C_296_102, V2C_448_102, V2C_545_102, V2C_578_102, V2C_782_102, V2C_858_102, V2C_891_102, V2C_953_102, V2C_988_102, V2C_1055_102, V2C_1071_102, V2C_1121_102, V2C_1253_102, V2C_1254_102, V2C_22_103, V2C_58_103, V2C_126_103, V2C_187_103, V2C_201_103, V2C_244_103, V2C_344_103, V2C_398_103, V2C_495_103, V2C_731_103, V2C_779_103, V2C_827_103, V2C_868_103, V2C_957_103, V2C_991_103, V2C_1030_103, V2C_1104_103, V2C_1115_103, V2C_1254_103, V2C_1255_103, V2C_31_104, V2C_80_104, V2C_136_104, V2C_184_104, V2C_213_104, V2C_282_104, V2C_333_104, V2C_392_104, V2C_481_104, V2C_641_104, V2C_702_104, V2C_822_104, V2C_912_104, V2C_927_104, V2C_1006_104, V2C_1038_104, V2C_1057_104, V2C_1136_104, V2C_1255_104, V2C_1256_104, V2C_26_105, V2C_53_105, V2C_118_105, V2C_152_105, V2C_218_105, V2C_285_105, V2C_382_105, V2C_389_105, V2C_548_105, V2C_605_105, V2C_633_105, V2C_737_105, V2C_868_105, V2C_960_105, V2C_985_105, V2C_1045_105, V2C_1075_105, V2C_1120_105, V2C_1256_105, V2C_1257_105, V2C_45_106, V2C_56_106, V2C_143_106, V2C_151_106, V2C_216_106, V2C_270_106, V2C_446_106, V2C_486_106, V2C_570_106, V2C_584_106, V2C_657_106, V2C_703_106, V2C_872_106, V2C_944_106, V2C_980_106, V2C_1010_106, V2C_1085_106, V2C_1149_106, V2C_1257_106, V2C_1258_106, V2C_16_107, V2C_74_107, V2C_109_107, V2C_180_107, V2C_196_107, V2C_262_107, V2C_311_107, V2C_378_107, V2C_457_107, V2C_691_107, V2C_755_107, V2C_809_107, V2C_887_107, V2C_935_107, V2C_978_107, V2C_1030_107, V2C_1079_107, V2C_1127_107, V2C_1258_107, V2C_1259_107, V2C_47_108, V2C_71_108, V2C_111_108, V2C_179_108, V2C_213_108, V2C_244_108, V2C_297_108, V2C_449_108, V2C_546_108, V2C_579_108, V2C_783_108, V2C_859_108, V2C_892_108, V2C_954_108, V2C_989_108, V2C_1056_108, V2C_1072_108, V2C_1122_108, V2C_1259_108, V2C_1260_108, V2C_23_109, V2C_59_109, V2C_127_109, V2C_188_109, V2C_202_109, V2C_245_109, V2C_345_109, V2C_399_109, V2C_496_109, V2C_732_109, V2C_780_109, V2C_828_109, V2C_869_109, V2C_958_109, V2C_992_109, V2C_1031_109, V2C_1057_109, V2C_1116_109, V2C_1260_109, V2C_1261_109, V2C_32_110, V2C_81_110, V2C_137_110, V2C_185_110, V2C_214_110, V2C_283_110, V2C_334_110, V2C_393_110, V2C_482_110, V2C_642_110, V2C_703_110, V2C_823_110, V2C_865_110, V2C_928_110, V2C_1007_110, V2C_1039_110, V2C_1058_110, V2C_1137_110, V2C_1261_110, V2C_1262_110, V2C_27_111, V2C_54_111, V2C_119_111, V2C_153_111, V2C_219_111, V2C_286_111, V2C_383_111, V2C_390_111, V2C_549_111, V2C_606_111, V2C_634_111, V2C_738_111, V2C_869_111, V2C_913_111, V2C_986_111, V2C_1046_111, V2C_1076_111, V2C_1121_111, V2C_1262_111, V2C_1263_111, V2C_46_112, V2C_57_112, V2C_144_112, V2C_152_112, V2C_217_112, V2C_271_112, V2C_447_112, V2C_487_112, V2C_571_112, V2C_585_112, V2C_658_112, V2C_704_112, V2C_873_112, V2C_945_112, V2C_981_112, V2C_1011_112, V2C_1086_112, V2C_1150_112, V2C_1263_112, V2C_1264_112, V2C_17_113, V2C_75_113, V2C_110_113, V2C_181_113, V2C_197_113, V2C_263_113, V2C_312_113, V2C_379_113, V2C_458_113, V2C_692_113, V2C_756_113, V2C_810_113, V2C_888_113, V2C_936_113, V2C_979_113, V2C_1031_113, V2C_1080_113, V2C_1128_113, V2C_1264_113, V2C_1265_113, V2C_48_114, V2C_72_114, V2C_112_114, V2C_180_114, V2C_214_114, V2C_245_114, V2C_298_114, V2C_450_114, V2C_547_114, V2C_580_114, V2C_784_114, V2C_860_114, V2C_893_114, V2C_955_114, V2C_990_114, V2C_1009_114, V2C_1073_114, V2C_1123_114, V2C_1265_114, V2C_1266_114, V2C_24_115, V2C_60_115, V2C_128_115, V2C_189_115, V2C_203_115, V2C_246_115, V2C_346_115, V2C_400_115, V2C_497_115, V2C_733_115, V2C_781_115, V2C_829_115, V2C_870_115, V2C_959_115, V2C_993_115, V2C_1032_115, V2C_1058_115, V2C_1117_115, V2C_1266_115, V2C_1267_115, V2C_33_116, V2C_82_116, V2C_138_116, V2C_186_116, V2C_215_116, V2C_284_116, V2C_335_116, V2C_394_116, V2C_483_116, V2C_643_116, V2C_704_116, V2C_824_116, V2C_866_116, V2C_929_116, V2C_1008_116, V2C_1040_116, V2C_1059_116, V2C_1138_116, V2C_1267_116, V2C_1268_116, V2C_28_117, V2C_55_117, V2C_120_117, V2C_154_117, V2C_220_117, V2C_287_117, V2C_384_117, V2C_391_117, V2C_550_117, V2C_607_117, V2C_635_117, V2C_739_117, V2C_870_117, V2C_914_117, V2C_987_117, V2C_1047_117, V2C_1077_117, V2C_1122_117, V2C_1268_117, V2C_1269_117, V2C_47_118, V2C_58_118, V2C_97_118, V2C_153_118, V2C_218_118, V2C_272_118, V2C_448_118, V2C_488_118, V2C_572_118, V2C_586_118, V2C_659_118, V2C_705_118, V2C_874_118, V2C_946_118, V2C_982_118, V2C_1012_118, V2C_1087_118, V2C_1151_118, V2C_1269_118, V2C_1270_118, V2C_18_119, V2C_76_119, V2C_111_119, V2C_182_119, V2C_198_119, V2C_264_119, V2C_313_119, V2C_380_119, V2C_459_119, V2C_693_119, V2C_757_119, V2C_811_119, V2C_889_119, V2C_937_119, V2C_980_119, V2C_1032_119, V2C_1081_119, V2C_1129_119, V2C_1270_119, V2C_1271_119, V2C_1_120, V2C_73_120, V2C_113_120, V2C_181_120, V2C_215_120, V2C_246_120, V2C_299_120, V2C_451_120, V2C_548_120, V2C_581_120, V2C_785_120, V2C_861_120, V2C_894_120, V2C_956_120, V2C_991_120, V2C_1010_120, V2C_1074_120, V2C_1124_120, V2C_1271_120, V2C_1272_120, V2C_25_121, V2C_61_121, V2C_129_121, V2C_190_121, V2C_204_121, V2C_247_121, V2C_347_121, V2C_401_121, V2C_498_121, V2C_734_121, V2C_782_121, V2C_830_121, V2C_871_121, V2C_960_121, V2C_994_121, V2C_1033_121, V2C_1059_121, V2C_1118_121, V2C_1272_121, V2C_1273_121, V2C_34_122, V2C_83_122, V2C_139_122, V2C_187_122, V2C_216_122, V2C_285_122, V2C_336_122, V2C_395_122, V2C_484_122, V2C_644_122, V2C_705_122, V2C_825_122, V2C_867_122, V2C_930_122, V2C_961_122, V2C_1041_122, V2C_1060_122, V2C_1139_122, V2C_1273_122, V2C_1274_122, V2C_29_123, V2C_56_123, V2C_121_123, V2C_155_123, V2C_221_123, V2C_288_123, V2C_337_123, V2C_392_123, V2C_551_123, V2C_608_123, V2C_636_123, V2C_740_123, V2C_871_123, V2C_915_123, V2C_988_123, V2C_1048_123, V2C_1078_123, V2C_1123_123, V2C_1274_123, V2C_1275_123, V2C_48_124, V2C_59_124, V2C_98_124, V2C_154_124, V2C_219_124, V2C_273_124, V2C_449_124, V2C_489_124, V2C_573_124, V2C_587_124, V2C_660_124, V2C_706_124, V2C_875_124, V2C_947_124, V2C_983_124, V2C_1013_124, V2C_1088_124, V2C_1152_124, V2C_1275_124, V2C_1276_124, V2C_19_125, V2C_77_125, V2C_112_125, V2C_183_125, V2C_199_125, V2C_265_125, V2C_314_125, V2C_381_125, V2C_460_125, V2C_694_125, V2C_758_125, V2C_812_125, V2C_890_125, V2C_938_125, V2C_981_125, V2C_1033_125, V2C_1082_125, V2C_1130_125, V2C_1276_125, V2C_1277_125, V2C_2_126, V2C_74_126, V2C_114_126, V2C_182_126, V2C_216_126, V2C_247_126, V2C_300_126, V2C_452_126, V2C_549_126, V2C_582_126, V2C_786_126, V2C_862_126, V2C_895_126, V2C_957_126, V2C_992_126, V2C_1011_126, V2C_1075_126, V2C_1125_126, V2C_1277_126, V2C_1278_126, V2C_26_127, V2C_62_127, V2C_130_127, V2C_191_127, V2C_205_127, V2C_248_127, V2C_348_127, V2C_402_127, V2C_499_127, V2C_735_127, V2C_783_127, V2C_831_127, V2C_872_127, V2C_913_127, V2C_995_127, V2C_1034_127, V2C_1060_127, V2C_1119_127, V2C_1278_127, V2C_1279_127, V2C_35_128, V2C_84_128, V2C_140_128, V2C_188_128, V2C_217_128, V2C_286_128, V2C_289_128, V2C_396_128, V2C_485_128, V2C_645_128, V2C_706_128, V2C_826_128, V2C_868_128, V2C_931_128, V2C_962_128, V2C_1042_128, V2C_1061_128, V2C_1140_128, V2C_1279_128, V2C_1280_128, V2C_30_129, V2C_57_129, V2C_122_129, V2C_156_129, V2C_222_129, V2C_241_129, V2C_338_129, V2C_393_129, V2C_552_129, V2C_609_129, V2C_637_129, V2C_741_129, V2C_872_129, V2C_916_129, V2C_989_129, V2C_1049_129, V2C_1079_129, V2C_1124_129, V2C_1280_129, V2C_1281_129, V2C_1_130, V2C_60_130, V2C_99_130, V2C_155_130, V2C_220_130, V2C_274_130, V2C_450_130, V2C_490_130, V2C_574_130, V2C_588_130, V2C_661_130, V2C_707_130, V2C_876_130, V2C_948_130, V2C_984_130, V2C_1014_130, V2C_1089_130, V2C_1105_130, V2C_1281_130, V2C_1282_130, V2C_20_131, V2C_78_131, V2C_113_131, V2C_184_131, V2C_200_131, V2C_266_131, V2C_315_131, V2C_382_131, V2C_461_131, V2C_695_131, V2C_759_131, V2C_813_131, V2C_891_131, V2C_939_131, V2C_982_131, V2C_1034_131, V2C_1083_131, V2C_1131_131, V2C_1282_131, V2C_1283_131, V2C_3_132, V2C_75_132, V2C_115_132, V2C_183_132, V2C_217_132, V2C_248_132, V2C_301_132, V2C_453_132, V2C_550_132, V2C_583_132, V2C_787_132, V2C_863_132, V2C_896_132, V2C_958_132, V2C_993_132, V2C_1012_132, V2C_1076_132, V2C_1126_132, V2C_1283_132, V2C_1284_132, V2C_27_133, V2C_63_133, V2C_131_133, V2C_192_133, V2C_206_133, V2C_249_133, V2C_349_133, V2C_403_133, V2C_500_133, V2C_736_133, V2C_784_133, V2C_832_133, V2C_873_133, V2C_914_133, V2C_996_133, V2C_1035_133, V2C_1061_133, V2C_1120_133, V2C_1284_133, V2C_1285_133, V2C_36_134, V2C_85_134, V2C_141_134, V2C_189_134, V2C_218_134, V2C_287_134, V2C_290_134, V2C_397_134, V2C_486_134, V2C_646_134, V2C_707_134, V2C_827_134, V2C_869_134, V2C_932_134, V2C_963_134, V2C_1043_134, V2C_1062_134, V2C_1141_134, V2C_1285_134, V2C_1286_134, V2C_31_135, V2C_58_135, V2C_123_135, V2C_157_135, V2C_223_135, V2C_242_135, V2C_339_135, V2C_394_135, V2C_553_135, V2C_610_135, V2C_638_135, V2C_742_135, V2C_873_135, V2C_917_135, V2C_990_135, V2C_1050_135, V2C_1080_135, V2C_1125_135, V2C_1286_135, V2C_1287_135, V2C_2_136, V2C_61_136, V2C_100_136, V2C_156_136, V2C_221_136, V2C_275_136, V2C_451_136, V2C_491_136, V2C_575_136, V2C_589_136, V2C_662_136, V2C_708_136, V2C_877_136, V2C_949_136, V2C_985_136, V2C_1015_136, V2C_1090_136, V2C_1106_136, V2C_1287_136, V2C_1288_136, V2C_21_137, V2C_79_137, V2C_114_137, V2C_185_137, V2C_201_137, V2C_267_137, V2C_316_137, V2C_383_137, V2C_462_137, V2C_696_137, V2C_760_137, V2C_814_137, V2C_892_137, V2C_940_137, V2C_983_137, V2C_1035_137, V2C_1084_137, V2C_1132_137, V2C_1288_137, V2C_1289_137, V2C_4_138, V2C_76_138, V2C_116_138, V2C_184_138, V2C_218_138, V2C_249_138, V2C_302_138, V2C_454_138, V2C_551_138, V2C_584_138, V2C_788_138, V2C_864_138, V2C_897_138, V2C_959_138, V2C_994_138, V2C_1013_138, V2C_1077_138, V2C_1127_138, V2C_1289_138, V2C_1290_138, V2C_28_139, V2C_64_139, V2C_132_139, V2C_145_139, V2C_207_139, V2C_250_139, V2C_350_139, V2C_404_139, V2C_501_139, V2C_737_139, V2C_785_139, V2C_833_139, V2C_874_139, V2C_915_139, V2C_997_139, V2C_1036_139, V2C_1062_139, V2C_1121_139, V2C_1290_139, V2C_1291_139, V2C_37_140, V2C_86_140, V2C_142_140, V2C_190_140, V2C_219_140, V2C_288_140, V2C_291_140, V2C_398_140, V2C_487_140, V2C_647_140, V2C_708_140, V2C_828_140, V2C_870_140, V2C_933_140, V2C_964_140, V2C_1044_140, V2C_1063_140, V2C_1142_140, V2C_1291_140, V2C_1292_140, V2C_32_141, V2C_59_141, V2C_124_141, V2C_158_141, V2C_224_141, V2C_243_141, V2C_340_141, V2C_395_141, V2C_554_141, V2C_611_141, V2C_639_141, V2C_743_141, V2C_874_141, V2C_918_141, V2C_991_141, V2C_1051_141, V2C_1081_141, V2C_1126_141, V2C_1292_141, V2C_1293_141, V2C_3_142, V2C_62_142, V2C_101_142, V2C_157_142, V2C_222_142, V2C_276_142, V2C_452_142, V2C_492_142, V2C_576_142, V2C_590_142, V2C_663_142, V2C_709_142, V2C_878_142, V2C_950_142, V2C_986_142, V2C_1016_142, V2C_1091_142, V2C_1107_142, V2C_1293_142, V2C_1294_142, V2C_22_143, V2C_80_143, V2C_115_143, V2C_186_143, V2C_202_143, V2C_268_143, V2C_317_143, V2C_384_143, V2C_463_143, V2C_697_143, V2C_761_143, V2C_815_143, V2C_893_143, V2C_941_143, V2C_984_143, V2C_1036_143, V2C_1085_143, V2C_1133_143, V2C_1294_143, V2C_1295_143, V2C_5_144, V2C_77_144, V2C_117_144, V2C_185_144, V2C_219_144, V2C_250_144, V2C_303_144, V2C_455_144, V2C_552_144, V2C_585_144, V2C_789_144, V2C_817_144, V2C_898_144, V2C_960_144, V2C_995_144, V2C_1014_144, V2C_1078_144, V2C_1128_144, V2C_1295_144, V2C_1296_144, V2C_29_145, V2C_65_145, V2C_133_145, V2C_146_145, V2C_208_145, V2C_251_145, V2C_351_145, V2C_405_145, V2C_502_145, V2C_738_145, V2C_786_145, V2C_834_145, V2C_875_145, V2C_916_145, V2C_998_145, V2C_1037_145, V2C_1063_145, V2C_1122_145, V2C_1296_145, V2C_1297_145, V2C_38_146, V2C_87_146, V2C_143_146, V2C_191_146, V2C_220_146, V2C_241_146, V2C_292_146, V2C_399_146, V2C_488_146, V2C_648_146, V2C_709_146, V2C_829_146, V2C_871_146, V2C_934_146, V2C_965_146, V2C_1045_146, V2C_1064_146, V2C_1143_146, V2C_1297_146, V2C_1298_146, V2C_33_147, V2C_60_147, V2C_125_147, V2C_159_147, V2C_225_147, V2C_244_147, V2C_341_147, V2C_396_147, V2C_555_147, V2C_612_147, V2C_640_147, V2C_744_147, V2C_875_147, V2C_919_147, V2C_992_147, V2C_1052_147, V2C_1082_147, V2C_1127_147, V2C_1298_147, V2C_1299_147, V2C_4_148, V2C_63_148, V2C_102_148, V2C_158_148, V2C_223_148, V2C_277_148, V2C_453_148, V2C_493_148, V2C_529_148, V2C_591_148, V2C_664_148, V2C_710_148, V2C_879_148, V2C_951_148, V2C_987_148, V2C_1017_148, V2C_1092_148, V2C_1108_148, V2C_1299_148, V2C_1300_148, V2C_23_149, V2C_81_149, V2C_116_149, V2C_187_149, V2C_203_149, V2C_269_149, V2C_318_149, V2C_337_149, V2C_464_149, V2C_698_149, V2C_762_149, V2C_816_149, V2C_894_149, V2C_942_149, V2C_985_149, V2C_1037_149, V2C_1086_149, V2C_1134_149, V2C_1300_149, V2C_1301_149, V2C_6_150, V2C_78_150, V2C_118_150, V2C_186_150, V2C_220_150, V2C_251_150, V2C_304_150, V2C_456_150, V2C_553_150, V2C_586_150, V2C_790_150, V2C_818_150, V2C_899_150, V2C_913_150, V2C_996_150, V2C_1015_150, V2C_1079_150, V2C_1129_150, V2C_1301_150, V2C_1302_150, V2C_30_151, V2C_66_151, V2C_134_151, V2C_147_151, V2C_209_151, V2C_252_151, V2C_352_151, V2C_406_151, V2C_503_151, V2C_739_151, V2C_787_151, V2C_835_151, V2C_876_151, V2C_917_151, V2C_999_151, V2C_1038_151, V2C_1064_151, V2C_1123_151, V2C_1302_151, V2C_1303_151, V2C_39_152, V2C_88_152, V2C_144_152, V2C_192_152, V2C_221_152, V2C_242_152, V2C_293_152, V2C_400_152, V2C_489_152, V2C_649_152, V2C_710_152, V2C_830_152, V2C_872_152, V2C_935_152, V2C_966_152, V2C_1046_152, V2C_1065_152, V2C_1144_152, V2C_1303_152, V2C_1304_152, V2C_34_153, V2C_61_153, V2C_126_153, V2C_160_153, V2C_226_153, V2C_245_153, V2C_342_153, V2C_397_153, V2C_556_153, V2C_613_153, V2C_641_153, V2C_745_153, V2C_876_153, V2C_920_153, V2C_993_153, V2C_1053_153, V2C_1083_153, V2C_1128_153, V2C_1304_153, V2C_1305_153, V2C_5_154, V2C_64_154, V2C_103_154, V2C_159_154, V2C_224_154, V2C_278_154, V2C_454_154, V2C_494_154, V2C_530_154, V2C_592_154, V2C_665_154, V2C_711_154, V2C_880_154, V2C_952_154, V2C_988_154, V2C_1018_154, V2C_1093_154, V2C_1109_154, V2C_1305_154, V2C_1306_154, V2C_24_155, V2C_82_155, V2C_117_155, V2C_188_155, V2C_204_155, V2C_270_155, V2C_319_155, V2C_338_155, V2C_465_155, V2C_699_155, V2C_763_155, V2C_769_155, V2C_895_155, V2C_943_155, V2C_986_155, V2C_1038_155, V2C_1087_155, V2C_1135_155, V2C_1306_155, V2C_1307_155, V2C_7_156, V2C_79_156, V2C_119_156, V2C_187_156, V2C_221_156, V2C_252_156, V2C_305_156, V2C_457_156, V2C_554_156, V2C_587_156, V2C_791_156, V2C_819_156, V2C_900_156, V2C_914_156, V2C_997_156, V2C_1016_156, V2C_1080_156, V2C_1130_156, V2C_1307_156, V2C_1308_156, V2C_31_157, V2C_67_157, V2C_135_157, V2C_148_157, V2C_210_157, V2C_253_157, V2C_353_157, V2C_407_157, V2C_504_157, V2C_740_157, V2C_788_157, V2C_836_157, V2C_877_157, V2C_918_157, V2C_1000_157, V2C_1039_157, V2C_1065_157, V2C_1124_157, V2C_1308_157, V2C_1309_157, V2C_40_158, V2C_89_158, V2C_97_158, V2C_145_158, V2C_222_158, V2C_243_158, V2C_294_158, V2C_401_158, V2C_490_158, V2C_650_158, V2C_711_158, V2C_831_158, V2C_873_158, V2C_936_158, V2C_967_158, V2C_1047_158, V2C_1066_158, V2C_1145_158, V2C_1309_158, V2C_1310_158, V2C_35_159, V2C_62_159, V2C_127_159, V2C_161_159, V2C_227_159, V2C_246_159, V2C_343_159, V2C_398_159, V2C_557_159, V2C_614_159, V2C_642_159, V2C_746_159, V2C_877_159, V2C_921_159, V2C_994_159, V2C_1054_159, V2C_1084_159, V2C_1129_159, V2C_1310_159, V2C_1311_159, V2C_6_160, V2C_65_160, V2C_104_160, V2C_160_160, V2C_225_160, V2C_279_160, V2C_455_160, V2C_495_160, V2C_531_160, V2C_593_160, V2C_666_160, V2C_712_160, V2C_881_160, V2C_953_160, V2C_989_160, V2C_1019_160, V2C_1094_160, V2C_1110_160, V2C_1311_160, V2C_1312_160, V2C_25_161, V2C_83_161, V2C_118_161, V2C_189_161, V2C_205_161, V2C_271_161, V2C_320_161, V2C_339_161, V2C_466_161, V2C_700_161, V2C_764_161, V2C_770_161, V2C_896_161, V2C_944_161, V2C_987_161, V2C_1039_161, V2C_1088_161, V2C_1136_161, V2C_1312_161, V2C_1313_161, V2C_8_162, V2C_80_162, V2C_120_162, V2C_188_162, V2C_222_162, V2C_253_162, V2C_306_162, V2C_458_162, V2C_555_162, V2C_588_162, V2C_792_162, V2C_820_162, V2C_901_162, V2C_915_162, V2C_998_162, V2C_1017_162, V2C_1081_162, V2C_1131_162, V2C_1313_162, V2C_1314_162, V2C_32_163, V2C_68_163, V2C_136_163, V2C_149_163, V2C_211_163, V2C_254_163, V2C_354_163, V2C_408_163, V2C_505_163, V2C_741_163, V2C_789_163, V2C_837_163, V2C_878_163, V2C_919_163, V2C_1001_163, V2C_1040_163, V2C_1066_163, V2C_1125_163, V2C_1314_163, V2C_1315_163, V2C_41_164, V2C_90_164, V2C_98_164, V2C_146_164, V2C_223_164, V2C_244_164, V2C_295_164, V2C_402_164, V2C_491_164, V2C_651_164, V2C_712_164, V2C_832_164, V2C_874_164, V2C_937_164, V2C_968_164, V2C_1048_164, V2C_1067_164, V2C_1146_164, V2C_1315_164, V2C_1316_164, V2C_36_165, V2C_63_165, V2C_128_165, V2C_162_165, V2C_228_165, V2C_247_165, V2C_344_165, V2C_399_165, V2C_558_165, V2C_615_165, V2C_643_165, V2C_747_165, V2C_878_165, V2C_922_165, V2C_995_165, V2C_1055_165, V2C_1085_165, V2C_1130_165, V2C_1316_165, V2C_1317_165, V2C_7_166, V2C_66_166, V2C_105_166, V2C_161_166, V2C_226_166, V2C_280_166, V2C_456_166, V2C_496_166, V2C_532_166, V2C_594_166, V2C_667_166, V2C_713_166, V2C_882_166, V2C_954_166, V2C_990_166, V2C_1020_166, V2C_1095_166, V2C_1111_166, V2C_1317_166, V2C_1318_166, V2C_26_167, V2C_84_167, V2C_119_167, V2C_190_167, V2C_206_167, V2C_272_167, V2C_321_167, V2C_340_167, V2C_467_167, V2C_701_167, V2C_765_167, V2C_771_167, V2C_897_167, V2C_945_167, V2C_988_167, V2C_1040_167, V2C_1089_167, V2C_1137_167, V2C_1318_167, V2C_1319_167, V2C_9_168, V2C_81_168, V2C_121_168, V2C_189_168, V2C_223_168, V2C_254_168, V2C_307_168, V2C_459_168, V2C_556_168, V2C_589_168, V2C_793_168, V2C_821_168, V2C_902_168, V2C_916_168, V2C_999_168, V2C_1018_168, V2C_1082_168, V2C_1132_168, V2C_1319_168, V2C_1320_168, V2C_33_169, V2C_69_169, V2C_137_169, V2C_150_169, V2C_212_169, V2C_255_169, V2C_355_169, V2C_409_169, V2C_506_169, V2C_742_169, V2C_790_169, V2C_838_169, V2C_879_169, V2C_920_169, V2C_1002_169, V2C_1041_169, V2C_1067_169, V2C_1126_169, V2C_1320_169, V2C_1321_169, V2C_42_170, V2C_91_170, V2C_99_170, V2C_147_170, V2C_224_170, V2C_245_170, V2C_296_170, V2C_403_170, V2C_492_170, V2C_652_170, V2C_713_170, V2C_833_170, V2C_875_170, V2C_938_170, V2C_969_170, V2C_1049_170, V2C_1068_170, V2C_1147_170, V2C_1321_170, V2C_1322_170, V2C_37_171, V2C_64_171, V2C_129_171, V2C_163_171, V2C_229_171, V2C_248_171, V2C_345_171, V2C_400_171, V2C_559_171, V2C_616_171, V2C_644_171, V2C_748_171, V2C_879_171, V2C_923_171, V2C_996_171, V2C_1056_171, V2C_1086_171, V2C_1131_171, V2C_1322_171, V2C_1323_171, V2C_8_172, V2C_67_172, V2C_106_172, V2C_162_172, V2C_227_172, V2C_281_172, V2C_457_172, V2C_497_172, V2C_533_172, V2C_595_172, V2C_668_172, V2C_714_172, V2C_883_172, V2C_955_172, V2C_991_172, V2C_1021_172, V2C_1096_172, V2C_1112_172, V2C_1323_172, V2C_1324_172, V2C_27_173, V2C_85_173, V2C_120_173, V2C_191_173, V2C_207_173, V2C_273_173, V2C_322_173, V2C_341_173, V2C_468_173, V2C_702_173, V2C_766_173, V2C_772_173, V2C_898_173, V2C_946_173, V2C_989_173, V2C_1041_173, V2C_1090_173, V2C_1138_173, V2C_1324_173, V2C_1325_173, V2C_10_174, V2C_82_174, V2C_122_174, V2C_190_174, V2C_224_174, V2C_255_174, V2C_308_174, V2C_460_174, V2C_557_174, V2C_590_174, V2C_794_174, V2C_822_174, V2C_903_174, V2C_917_174, V2C_1000_174, V2C_1019_174, V2C_1083_174, V2C_1133_174, V2C_1325_174, V2C_1326_174, V2C_34_175, V2C_70_175, V2C_138_175, V2C_151_175, V2C_213_175, V2C_256_175, V2C_356_175, V2C_410_175, V2C_507_175, V2C_743_175, V2C_791_175, V2C_839_175, V2C_880_175, V2C_921_175, V2C_1003_175, V2C_1042_175, V2C_1068_175, V2C_1127_175, V2C_1326_175, V2C_1327_175, V2C_43_176, V2C_92_176, V2C_100_176, V2C_148_176, V2C_225_176, V2C_246_176, V2C_297_176, V2C_404_176, V2C_493_176, V2C_653_176, V2C_714_176, V2C_834_176, V2C_876_176, V2C_939_176, V2C_970_176, V2C_1050_176, V2C_1069_176, V2C_1148_176, V2C_1327_176, V2C_1328_176, V2C_38_177, V2C_65_177, V2C_130_177, V2C_164_177, V2C_230_177, V2C_249_177, V2C_346_177, V2C_401_177, V2C_560_177, V2C_617_177, V2C_645_177, V2C_749_177, V2C_880_177, V2C_924_177, V2C_997_177, V2C_1009_177, V2C_1087_177, V2C_1132_177, V2C_1328_177, V2C_1329_177, V2C_9_178, V2C_68_178, V2C_107_178, V2C_163_178, V2C_228_178, V2C_282_178, V2C_458_178, V2C_498_178, V2C_534_178, V2C_596_178, V2C_669_178, V2C_715_178, V2C_884_178, V2C_956_178, V2C_992_178, V2C_1022_178, V2C_1097_178, V2C_1113_178, V2C_1329_178, V2C_1330_178, V2C_28_179, V2C_86_179, V2C_121_179, V2C_192_179, V2C_208_179, V2C_274_179, V2C_323_179, V2C_342_179, V2C_469_179, V2C_703_179, V2C_767_179, V2C_773_179, V2C_899_179, V2C_947_179, V2C_990_179, V2C_1042_179, V2C_1091_179, V2C_1139_179, V2C_1330_179, V2C_1331_179, V2C_11_180, V2C_83_180, V2C_123_180, V2C_191_180, V2C_225_180, V2C_256_180, V2C_309_180, V2C_461_180, V2C_558_180, V2C_591_180, V2C_795_180, V2C_823_180, V2C_904_180, V2C_918_180, V2C_1001_180, V2C_1020_180, V2C_1084_180, V2C_1134_180, V2C_1331_180, V2C_1332_180, V2C_35_181, V2C_71_181, V2C_139_181, V2C_152_181, V2C_214_181, V2C_257_181, V2C_357_181, V2C_411_181, V2C_508_181, V2C_744_181, V2C_792_181, V2C_840_181, V2C_881_181, V2C_922_181, V2C_1004_181, V2C_1043_181, V2C_1069_181, V2C_1128_181, V2C_1332_181, V2C_1333_181, V2C_44_182, V2C_93_182, V2C_101_182, V2C_149_182, V2C_226_182, V2C_247_182, V2C_298_182, V2C_405_182, V2C_494_182, V2C_654_182, V2C_715_182, V2C_835_182, V2C_877_182, V2C_940_182, V2C_971_182, V2C_1051_182, V2C_1070_182, V2C_1149_182, V2C_1333_182, V2C_1334_182, V2C_39_183, V2C_66_183, V2C_131_183, V2C_165_183, V2C_231_183, V2C_250_183, V2C_347_183, V2C_402_183, V2C_561_183, V2C_618_183, V2C_646_183, V2C_750_183, V2C_881_183, V2C_925_183, V2C_998_183, V2C_1010_183, V2C_1088_183, V2C_1133_183, V2C_1334_183, V2C_1335_183, V2C_10_184, V2C_69_184, V2C_108_184, V2C_164_184, V2C_229_184, V2C_283_184, V2C_459_184, V2C_499_184, V2C_535_184, V2C_597_184, V2C_670_184, V2C_716_184, V2C_885_184, V2C_957_184, V2C_993_184, V2C_1023_184, V2C_1098_184, V2C_1114_184, V2C_1335_184, V2C_1336_184, V2C_29_185, V2C_87_185, V2C_122_185, V2C_145_185, V2C_209_185, V2C_275_185, V2C_324_185, V2C_343_185, V2C_470_185, V2C_704_185, V2C_768_185, V2C_774_185, V2C_900_185, V2C_948_185, V2C_991_185, V2C_1043_185, V2C_1092_185, V2C_1140_185, V2C_1336_185, V2C_1337_185, V2C_12_186, V2C_84_186, V2C_124_186, V2C_192_186, V2C_226_186, V2C_257_186, V2C_310_186, V2C_462_186, V2C_559_186, V2C_592_186, V2C_796_186, V2C_824_186, V2C_905_186, V2C_919_186, V2C_1002_186, V2C_1021_186, V2C_1085_186, V2C_1135_186, V2C_1337_186, V2C_1338_186, V2C_36_187, V2C_72_187, V2C_140_187, V2C_153_187, V2C_215_187, V2C_258_187, V2C_358_187, V2C_412_187, V2C_509_187, V2C_745_187, V2C_793_187, V2C_841_187, V2C_882_187, V2C_923_187, V2C_1005_187, V2C_1044_187, V2C_1070_187, V2C_1129_187, V2C_1338_187, V2C_1339_187, V2C_45_188, V2C_94_188, V2C_102_188, V2C_150_188, V2C_227_188, V2C_248_188, V2C_299_188, V2C_406_188, V2C_495_188, V2C_655_188, V2C_716_188, V2C_836_188, V2C_878_188, V2C_941_188, V2C_972_188, V2C_1052_188, V2C_1071_188, V2C_1150_188, V2C_1339_188, V2C_1340_188, V2C_40_189, V2C_67_189, V2C_132_189, V2C_166_189, V2C_232_189, V2C_251_189, V2C_348_189, V2C_403_189, V2C_562_189, V2C_619_189, V2C_647_189, V2C_751_189, V2C_882_189, V2C_926_189, V2C_999_189, V2C_1011_189, V2C_1089_189, V2C_1134_189, V2C_1340_189, V2C_1341_189, V2C_11_190, V2C_70_190, V2C_109_190, V2C_165_190, V2C_230_190, V2C_284_190, V2C_460_190, V2C_500_190, V2C_536_190, V2C_598_190, V2C_671_190, V2C_717_190, V2C_886_190, V2C_958_190, V2C_994_190, V2C_1024_190, V2C_1099_190, V2C_1115_190, V2C_1341_190, V2C_1342_190, V2C_30_191, V2C_88_191, V2C_123_191, V2C_146_191, V2C_210_191, V2C_276_191, V2C_325_191, V2C_344_191, V2C_471_191, V2C_705_191, V2C_721_191, V2C_775_191, V2C_901_191, V2C_949_191, V2C_992_191, V2C_1044_191, V2C_1093_191, V2C_1141_191, V2C_1342_191, V2C_1343_191, V2C_13_192, V2C_85_192, V2C_125_192, V2C_145_192, V2C_227_192, V2C_258_192, V2C_311_192, V2C_463_192, V2C_560_192, V2C_593_192, V2C_797_192, V2C_825_192, V2C_906_192, V2C_920_192, V2C_1003_192, V2C_1022_192, V2C_1086_192, V2C_1136_192, V2C_1343_192, V2C_1344_192, V2C_37_193, V2C_73_193, V2C_141_193, V2C_154_193, V2C_216_193, V2C_259_193, V2C_359_193, V2C_413_193, V2C_510_193, V2C_746_193, V2C_794_193, V2C_842_193, V2C_883_193, V2C_924_193, V2C_1006_193, V2C_1045_193, V2C_1071_193, V2C_1130_193, V2C_1344_193, V2C_1345_193, V2C_46_194, V2C_95_194, V2C_103_194, V2C_151_194, V2C_228_194, V2C_249_194, V2C_300_194, V2C_407_194, V2C_496_194, V2C_656_194, V2C_717_194, V2C_837_194, V2C_879_194, V2C_942_194, V2C_973_194, V2C_1053_194, V2C_1072_194, V2C_1151_194, V2C_1345_194, V2C_1346_194, V2C_41_195, V2C_68_195, V2C_133_195, V2C_167_195, V2C_233_195, V2C_252_195, V2C_349_195, V2C_404_195, V2C_563_195, V2C_620_195, V2C_648_195, V2C_752_195, V2C_883_195, V2C_927_195, V2C_1000_195, V2C_1012_195, V2C_1090_195, V2C_1135_195, V2C_1346_195, V2C_1347_195, V2C_12_196, V2C_71_196, V2C_110_196, V2C_166_196, V2C_231_196, V2C_285_196, V2C_461_196, V2C_501_196, V2C_537_196, V2C_599_196, V2C_672_196, V2C_718_196, V2C_887_196, V2C_959_196, V2C_995_196, V2C_1025_196, V2C_1100_196, V2C_1116_196, V2C_1347_196, V2C_1348_196, V2C_31_197, V2C_89_197, V2C_124_197, V2C_147_197, V2C_211_197, V2C_277_197, V2C_326_197, V2C_345_197, V2C_472_197, V2C_706_197, V2C_722_197, V2C_776_197, V2C_902_197, V2C_950_197, V2C_993_197, V2C_1045_197, V2C_1094_197, V2C_1142_197, V2C_1348_197, V2C_1349_197, V2C_14_198, V2C_86_198, V2C_126_198, V2C_146_198, V2C_228_198, V2C_259_198, V2C_312_198, V2C_464_198, V2C_561_198, V2C_594_198, V2C_798_198, V2C_826_198, V2C_907_198, V2C_921_198, V2C_1004_198, V2C_1023_198, V2C_1087_198, V2C_1137_198, V2C_1349_198, V2C_1350_198, V2C_38_199, V2C_74_199, V2C_142_199, V2C_155_199, V2C_217_199, V2C_260_199, V2C_360_199, V2C_414_199, V2C_511_199, V2C_747_199, V2C_795_199, V2C_843_199, V2C_884_199, V2C_925_199, V2C_1007_199, V2C_1046_199, V2C_1072_199, V2C_1131_199, V2C_1350_199, V2C_1351_199, V2C_47_200, V2C_96_200, V2C_104_200, V2C_152_200, V2C_229_200, V2C_250_200, V2C_301_200, V2C_408_200, V2C_497_200, V2C_657_200, V2C_718_200, V2C_838_200, V2C_880_200, V2C_943_200, V2C_974_200, V2C_1054_200, V2C_1073_200, V2C_1152_200, V2C_1351_200, V2C_1352_200, V2C_42_201, V2C_69_201, V2C_134_201, V2C_168_201, V2C_234_201, V2C_253_201, V2C_350_201, V2C_405_201, V2C_564_201, V2C_621_201, V2C_649_201, V2C_753_201, V2C_884_201, V2C_928_201, V2C_1001_201, V2C_1013_201, V2C_1091_201, V2C_1136_201, V2C_1352_201, V2C_1353_201, V2C_13_202, V2C_72_202, V2C_111_202, V2C_167_202, V2C_232_202, V2C_286_202, V2C_462_202, V2C_502_202, V2C_538_202, V2C_600_202, V2C_625_202, V2C_719_202, V2C_888_202, V2C_960_202, V2C_996_202, V2C_1026_202, V2C_1101_202, V2C_1117_202, V2C_1353_202, V2C_1354_202, V2C_32_203, V2C_90_203, V2C_125_203, V2C_148_203, V2C_212_203, V2C_278_203, V2C_327_203, V2C_346_203, V2C_473_203, V2C_707_203, V2C_723_203, V2C_777_203, V2C_903_203, V2C_951_203, V2C_994_203, V2C_1046_203, V2C_1095_203, V2C_1143_203, V2C_1354_203, V2C_1355_203, V2C_15_204, V2C_87_204, V2C_127_204, V2C_147_204, V2C_229_204, V2C_260_204, V2C_313_204, V2C_465_204, V2C_562_204, V2C_595_204, V2C_799_204, V2C_827_204, V2C_908_204, V2C_922_204, V2C_1005_204, V2C_1024_204, V2C_1088_204, V2C_1138_204, V2C_1355_204, V2C_1356_204, V2C_39_205, V2C_75_205, V2C_143_205, V2C_156_205, V2C_218_205, V2C_261_205, V2C_361_205, V2C_415_205, V2C_512_205, V2C_748_205, V2C_796_205, V2C_844_205, V2C_885_205, V2C_926_205, V2C_1008_205, V2C_1047_205, V2C_1073_205, V2C_1132_205, V2C_1356_205, V2C_1357_205, V2C_48_206, V2C_49_206, V2C_105_206, V2C_153_206, V2C_230_206, V2C_251_206, V2C_302_206, V2C_409_206, V2C_498_206, V2C_658_206, V2C_719_206, V2C_839_206, V2C_881_206, V2C_944_206, V2C_975_206, V2C_1055_206, V2C_1074_206, V2C_1105_206, V2C_1357_206, V2C_1358_206, V2C_43_207, V2C_70_207, V2C_135_207, V2C_169_207, V2C_235_207, V2C_254_207, V2C_351_207, V2C_406_207, V2C_565_207, V2C_622_207, V2C_650_207, V2C_754_207, V2C_885_207, V2C_929_207, V2C_1002_207, V2C_1014_207, V2C_1092_207, V2C_1137_207, V2C_1358_207, V2C_1359_207, V2C_14_208, V2C_73_208, V2C_112_208, V2C_168_208, V2C_233_208, V2C_287_208, V2C_463_208, V2C_503_208, V2C_539_208, V2C_601_208, V2C_626_208, V2C_720_208, V2C_889_208, V2C_913_208, V2C_997_208, V2C_1027_208, V2C_1102_208, V2C_1118_208, V2C_1359_208, V2C_1360_208, V2C_33_209, V2C_91_209, V2C_126_209, V2C_149_209, V2C_213_209, V2C_279_209, V2C_328_209, V2C_347_209, V2C_474_209, V2C_708_209, V2C_724_209, V2C_778_209, V2C_904_209, V2C_952_209, V2C_995_209, V2C_1047_209, V2C_1096_209, V2C_1144_209, V2C_1360_209, V2C_1361_209, V2C_16_210, V2C_88_210, V2C_128_210, V2C_148_210, V2C_230_210, V2C_261_210, V2C_314_210, V2C_466_210, V2C_563_210, V2C_596_210, V2C_800_210, V2C_828_210, V2C_909_210, V2C_923_210, V2C_1006_210, V2C_1025_210, V2C_1089_210, V2C_1139_210, V2C_1361_210, V2C_1362_210, V2C_40_211, V2C_76_211, V2C_144_211, V2C_157_211, V2C_219_211, V2C_262_211, V2C_362_211, V2C_416_211, V2C_513_211, V2C_749_211, V2C_797_211, V2C_845_211, V2C_886_211, V2C_927_211, V2C_961_211, V2C_1048_211, V2C_1074_211, V2C_1133_211, V2C_1362_211, V2C_1363_211, V2C_1_212, V2C_50_212, V2C_106_212, V2C_154_212, V2C_231_212, V2C_252_212, V2C_303_212, V2C_410_212, V2C_499_212, V2C_659_212, V2C_720_212, V2C_840_212, V2C_882_212, V2C_945_212, V2C_976_212, V2C_1056_212, V2C_1075_212, V2C_1106_212, V2C_1363_212, V2C_1364_212, V2C_44_213, V2C_71_213, V2C_136_213, V2C_170_213, V2C_236_213, V2C_255_213, V2C_352_213, V2C_407_213, V2C_566_213, V2C_623_213, V2C_651_213, V2C_755_213, V2C_886_213, V2C_930_213, V2C_1003_213, V2C_1015_213, V2C_1093_213, V2C_1138_213, V2C_1364_213, V2C_1365_213, V2C_15_214, V2C_74_214, V2C_113_214, V2C_169_214, V2C_234_214, V2C_288_214, V2C_464_214, V2C_504_214, V2C_540_214, V2C_602_214, V2C_627_214, V2C_673_214, V2C_890_214, V2C_914_214, V2C_998_214, V2C_1028_214, V2C_1103_214, V2C_1119_214, V2C_1365_214, V2C_1366_214, V2C_34_215, V2C_92_215, V2C_127_215, V2C_150_215, V2C_214_215, V2C_280_215, V2C_329_215, V2C_348_215, V2C_475_215, V2C_709_215, V2C_725_215, V2C_779_215, V2C_905_215, V2C_953_215, V2C_996_215, V2C_1048_215, V2C_1097_215, V2C_1145_215, V2C_1366_215, V2C_1367_215, V2C_17_216, V2C_89_216, V2C_129_216, V2C_149_216, V2C_231_216, V2C_262_216, V2C_315_216, V2C_467_216, V2C_564_216, V2C_597_216, V2C_801_216, V2C_829_216, V2C_910_216, V2C_924_216, V2C_1007_216, V2C_1026_216, V2C_1090_216, V2C_1140_216, V2C_1367_216, V2C_1368_216, V2C_41_217, V2C_77_217, V2C_97_217, V2C_158_217, V2C_220_217, V2C_263_217, V2C_363_217, V2C_417_217, V2C_514_217, V2C_750_217, V2C_798_217, V2C_846_217, V2C_887_217, V2C_928_217, V2C_962_217, V2C_1049_217, V2C_1075_217, V2C_1134_217, V2C_1368_217, V2C_1369_217, V2C_2_218, V2C_51_218, V2C_107_218, V2C_155_218, V2C_232_218, V2C_253_218, V2C_304_218, V2C_411_218, V2C_500_218, V2C_660_218, V2C_673_218, V2C_841_218, V2C_883_218, V2C_946_218, V2C_977_218, V2C_1009_218, V2C_1076_218, V2C_1107_218, V2C_1369_218, V2C_1370_218, V2C_45_219, V2C_72_219, V2C_137_219, V2C_171_219, V2C_237_219, V2C_256_219, V2C_353_219, V2C_408_219, V2C_567_219, V2C_624_219, V2C_652_219, V2C_756_219, V2C_887_219, V2C_931_219, V2C_1004_219, V2C_1016_219, V2C_1094_219, V2C_1139_219, V2C_1370_219, V2C_1371_219, V2C_16_220, V2C_75_220, V2C_114_220, V2C_170_220, V2C_235_220, V2C_241_220, V2C_465_220, V2C_505_220, V2C_541_220, V2C_603_220, V2C_628_220, V2C_674_220, V2C_891_220, V2C_915_220, V2C_999_220, V2C_1029_220, V2C_1104_220, V2C_1120_220, V2C_1371_220, V2C_1372_220, V2C_35_221, V2C_93_221, V2C_128_221, V2C_151_221, V2C_215_221, V2C_281_221, V2C_330_221, V2C_349_221, V2C_476_221, V2C_710_221, V2C_726_221, V2C_780_221, V2C_906_221, V2C_954_221, V2C_997_221, V2C_1049_221, V2C_1098_221, V2C_1146_221, V2C_1372_221, V2C_1373_221, V2C_18_222, V2C_90_222, V2C_130_222, V2C_150_222, V2C_232_222, V2C_263_222, V2C_316_222, V2C_468_222, V2C_565_222, V2C_598_222, V2C_802_222, V2C_830_222, V2C_911_222, V2C_925_222, V2C_1008_222, V2C_1027_222, V2C_1091_222, V2C_1141_222, V2C_1373_222, V2C_1374_222, V2C_42_223, V2C_78_223, V2C_98_223, V2C_159_223, V2C_221_223, V2C_264_223, V2C_364_223, V2C_418_223, V2C_515_223, V2C_751_223, V2C_799_223, V2C_847_223, V2C_888_223, V2C_929_223, V2C_963_223, V2C_1050_223, V2C_1076_223, V2C_1135_223, V2C_1374_223, V2C_1375_223, V2C_3_224, V2C_52_224, V2C_108_224, V2C_156_224, V2C_233_224, V2C_254_224, V2C_305_224, V2C_412_224, V2C_501_224, V2C_661_224, V2C_674_224, V2C_842_224, V2C_884_224, V2C_947_224, V2C_978_224, V2C_1010_224, V2C_1077_224, V2C_1108_224, V2C_1375_224, V2C_1376_224, V2C_46_225, V2C_73_225, V2C_138_225, V2C_172_225, V2C_238_225, V2C_257_225, V2C_354_225, V2C_409_225, V2C_568_225, V2C_577_225, V2C_653_225, V2C_757_225, V2C_888_225, V2C_932_225, V2C_1005_225, V2C_1017_225, V2C_1095_225, V2C_1140_225, V2C_1376_225, V2C_1377_225, V2C_17_226, V2C_76_226, V2C_115_226, V2C_171_226, V2C_236_226, V2C_242_226, V2C_466_226, V2C_506_226, V2C_542_226, V2C_604_226, V2C_629_226, V2C_675_226, V2C_892_226, V2C_916_226, V2C_1000_226, V2C_1030_226, V2C_1057_226, V2C_1121_226, V2C_1377_226, V2C_1378_226, V2C_36_227, V2C_94_227, V2C_129_227, V2C_152_227, V2C_216_227, V2C_282_227, V2C_331_227, V2C_350_227, V2C_477_227, V2C_711_227, V2C_727_227, V2C_781_227, V2C_907_227, V2C_955_227, V2C_998_227, V2C_1050_227, V2C_1099_227, V2C_1147_227, V2C_1378_227, V2C_1379_227, V2C_19_228, V2C_91_228, V2C_131_228, V2C_151_228, V2C_233_228, V2C_264_228, V2C_317_228, V2C_469_228, V2C_566_228, V2C_599_228, V2C_803_228, V2C_831_228, V2C_912_228, V2C_926_228, V2C_961_228, V2C_1028_228, V2C_1092_228, V2C_1142_228, V2C_1379_228, V2C_1380_228, V2C_43_229, V2C_79_229, V2C_99_229, V2C_160_229, V2C_222_229, V2C_265_229, V2C_365_229, V2C_419_229, V2C_516_229, V2C_752_229, V2C_800_229, V2C_848_229, V2C_889_229, V2C_930_229, V2C_964_229, V2C_1051_229, V2C_1077_229, V2C_1136_229, V2C_1380_229, V2C_1381_229, V2C_4_230, V2C_53_230, V2C_109_230, V2C_157_230, V2C_234_230, V2C_255_230, V2C_306_230, V2C_413_230, V2C_502_230, V2C_662_230, V2C_675_230, V2C_843_230, V2C_885_230, V2C_948_230, V2C_979_230, V2C_1011_230, V2C_1078_230, V2C_1109_230, V2C_1381_230, V2C_1382_230, V2C_47_231, V2C_74_231, V2C_139_231, V2C_173_231, V2C_239_231, V2C_258_231, V2C_355_231, V2C_410_231, V2C_569_231, V2C_578_231, V2C_654_231, V2C_758_231, V2C_889_231, V2C_933_231, V2C_1006_231, V2C_1018_231, V2C_1096_231, V2C_1141_231, V2C_1382_231, V2C_1383_231, V2C_18_232, V2C_77_232, V2C_116_232, V2C_172_232, V2C_237_232, V2C_243_232, V2C_467_232, V2C_507_232, V2C_543_232, V2C_605_232, V2C_630_232, V2C_676_232, V2C_893_232, V2C_917_232, V2C_1001_232, V2C_1031_232, V2C_1058_232, V2C_1122_232, V2C_1383_232, V2C_1384_232, V2C_37_233, V2C_95_233, V2C_130_233, V2C_153_233, V2C_217_233, V2C_283_233, V2C_332_233, V2C_351_233, V2C_478_233, V2C_712_233, V2C_728_233, V2C_782_233, V2C_908_233, V2C_956_233, V2C_999_233, V2C_1051_233, V2C_1100_233, V2C_1148_233, V2C_1384_233, V2C_1385_233, V2C_20_234, V2C_92_234, V2C_132_234, V2C_152_234, V2C_234_234, V2C_265_234, V2C_318_234, V2C_470_234, V2C_567_234, V2C_600_234, V2C_804_234, V2C_832_234, V2C_865_234, V2C_927_234, V2C_962_234, V2C_1029_234, V2C_1093_234, V2C_1143_234, V2C_1385_234, V2C_1386_234, V2C_44_235, V2C_80_235, V2C_100_235, V2C_161_235, V2C_223_235, V2C_266_235, V2C_366_235, V2C_420_235, V2C_517_235, V2C_753_235, V2C_801_235, V2C_849_235, V2C_890_235, V2C_931_235, V2C_965_235, V2C_1052_235, V2C_1078_235, V2C_1137_235, V2C_1386_235, V2C_1387_235, V2C_5_236, V2C_54_236, V2C_110_236, V2C_158_236, V2C_235_236, V2C_256_236, V2C_307_236, V2C_414_236, V2C_503_236, V2C_663_236, V2C_676_236, V2C_844_236, V2C_886_236, V2C_949_236, V2C_980_236, V2C_1012_236, V2C_1079_236, V2C_1110_236, V2C_1387_236, V2C_1388_236, V2C_48_237, V2C_75_237, V2C_140_237, V2C_174_237, V2C_240_237, V2C_259_237, V2C_356_237, V2C_411_237, V2C_570_237, V2C_579_237, V2C_655_237, V2C_759_237, V2C_890_237, V2C_934_237, V2C_1007_237, V2C_1019_237, V2C_1097_237, V2C_1142_237, V2C_1388_237, V2C_1389_237, V2C_19_238, V2C_78_238, V2C_117_238, V2C_173_238, V2C_238_238, V2C_244_238, V2C_468_238, V2C_508_238, V2C_544_238, V2C_606_238, V2C_631_238, V2C_677_238, V2C_894_238, V2C_918_238, V2C_1002_238, V2C_1032_238, V2C_1059_238, V2C_1123_238, V2C_1389_238, V2C_1390_238, V2C_38_239, V2C_96_239, V2C_131_239, V2C_154_239, V2C_218_239, V2C_284_239, V2C_333_239, V2C_352_239, V2C_479_239, V2C_713_239, V2C_729_239, V2C_783_239, V2C_909_239, V2C_957_239, V2C_1000_239, V2C_1052_239, V2C_1101_239, V2C_1149_239, V2C_1390_239, V2C_1391_239, V2C_21_240, V2C_93_240, V2C_133_240, V2C_153_240, V2C_235_240, V2C_266_240, V2C_319_240, V2C_471_240, V2C_568_240, V2C_601_240, V2C_805_240, V2C_833_240, V2C_866_240, V2C_928_240, V2C_963_240, V2C_1030_240, V2C_1094_240, V2C_1144_240, V2C_1391_240, V2C_1392_240, V2C_45_241, V2C_81_241, V2C_101_241, V2C_162_241, V2C_224_241, V2C_267_241, V2C_367_241, V2C_421_241, V2C_518_241, V2C_754_241, V2C_802_241, V2C_850_241, V2C_891_241, V2C_932_241, V2C_966_241, V2C_1053_241, V2C_1079_241, V2C_1138_241, V2C_1392_241, V2C_1393_241, V2C_6_242, V2C_55_242, V2C_111_242, V2C_159_242, V2C_236_242, V2C_257_242, V2C_308_242, V2C_415_242, V2C_504_242, V2C_664_242, V2C_677_242, V2C_845_242, V2C_887_242, V2C_950_242, V2C_981_242, V2C_1013_242, V2C_1080_242, V2C_1111_242, V2C_1393_242, V2C_1394_242, V2C_1_243, V2C_76_243, V2C_141_243, V2C_175_243, V2C_193_243, V2C_260_243, V2C_357_243, V2C_412_243, V2C_571_243, V2C_580_243, V2C_656_243, V2C_760_243, V2C_891_243, V2C_935_243, V2C_1008_243, V2C_1020_243, V2C_1098_243, V2C_1143_243, V2C_1394_243, V2C_1395_243, V2C_20_244, V2C_79_244, V2C_118_244, V2C_174_244, V2C_239_244, V2C_245_244, V2C_469_244, V2C_509_244, V2C_545_244, V2C_607_244, V2C_632_244, V2C_678_244, V2C_895_244, V2C_919_244, V2C_1003_244, V2C_1033_244, V2C_1060_244, V2C_1124_244, V2C_1395_244, V2C_1396_244, V2C_39_245, V2C_49_245, V2C_132_245, V2C_155_245, V2C_219_245, V2C_285_245, V2C_334_245, V2C_353_245, V2C_480_245, V2C_714_245, V2C_730_245, V2C_784_245, V2C_910_245, V2C_958_245, V2C_1001_245, V2C_1053_245, V2C_1102_245, V2C_1150_245, V2C_1396_245, V2C_1397_245, V2C_22_246, V2C_94_246, V2C_134_246, V2C_154_246, V2C_236_246, V2C_267_246, V2C_320_246, V2C_472_246, V2C_569_246, V2C_602_246, V2C_806_246, V2C_834_246, V2C_867_246, V2C_929_246, V2C_964_246, V2C_1031_246, V2C_1095_246, V2C_1145_246, V2C_1397_246, V2C_1398_246, V2C_46_247, V2C_82_247, V2C_102_247, V2C_163_247, V2C_225_247, V2C_268_247, V2C_368_247, V2C_422_247, V2C_519_247, V2C_755_247, V2C_803_247, V2C_851_247, V2C_892_247, V2C_933_247, V2C_967_247, V2C_1054_247, V2C_1080_247, V2C_1139_247, V2C_1398_247, V2C_1399_247, V2C_7_248, V2C_56_248, V2C_112_248, V2C_160_248, V2C_237_248, V2C_258_248, V2C_309_248, V2C_416_248, V2C_505_248, V2C_665_248, V2C_678_248, V2C_846_248, V2C_888_248, V2C_951_248, V2C_982_248, V2C_1014_248, V2C_1081_248, V2C_1112_248, V2C_1399_248, V2C_1400_248, V2C_2_249, V2C_77_249, V2C_142_249, V2C_176_249, V2C_194_249, V2C_261_249, V2C_358_249, V2C_413_249, V2C_572_249, V2C_581_249, V2C_657_249, V2C_761_249, V2C_892_249, V2C_936_249, V2C_961_249, V2C_1021_249, V2C_1099_249, V2C_1144_249, V2C_1400_249, V2C_1401_249, V2C_21_250, V2C_80_250, V2C_119_250, V2C_175_250, V2C_240_250, V2C_246_250, V2C_470_250, V2C_510_250, V2C_546_250, V2C_608_250, V2C_633_250, V2C_679_250, V2C_896_250, V2C_920_250, V2C_1004_250, V2C_1034_250, V2C_1061_250, V2C_1125_250, V2C_1401_250, V2C_1402_250, V2C_40_251, V2C_50_251, V2C_133_251, V2C_156_251, V2C_220_251, V2C_286_251, V2C_335_251, V2C_354_251, V2C_433_251, V2C_715_251, V2C_731_251, V2C_785_251, V2C_911_251, V2C_959_251, V2C_1002_251, V2C_1054_251, V2C_1103_251, V2C_1151_251, V2C_1402_251, V2C_1403_251, V2C_23_252, V2C_95_252, V2C_135_252, V2C_155_252, V2C_237_252, V2C_268_252, V2C_321_252, V2C_473_252, V2C_570_252, V2C_603_252, V2C_807_252, V2C_835_252, V2C_868_252, V2C_930_252, V2C_965_252, V2C_1032_252, V2C_1096_252, V2C_1146_252, V2C_1403_252, V2C_1404_252, V2C_47_253, V2C_83_253, V2C_103_253, V2C_164_253, V2C_226_253, V2C_269_253, V2C_369_253, V2C_423_253, V2C_520_253, V2C_756_253, V2C_804_253, V2C_852_253, V2C_893_253, V2C_934_253, V2C_968_253, V2C_1055_253, V2C_1081_253, V2C_1140_253, V2C_1404_253, V2C_1405_253, V2C_8_254, V2C_57_254, V2C_113_254, V2C_161_254, V2C_238_254, V2C_259_254, V2C_310_254, V2C_417_254, V2C_506_254, V2C_666_254, V2C_679_254, V2C_847_254, V2C_889_254, V2C_952_254, V2C_983_254, V2C_1015_254, V2C_1082_254, V2C_1113_254, V2C_1405_254, V2C_1406_254, V2C_3_255, V2C_78_255, V2C_143_255, V2C_177_255, V2C_195_255, V2C_262_255, V2C_359_255, V2C_414_255, V2C_573_255, V2C_582_255, V2C_658_255, V2C_762_255, V2C_893_255, V2C_937_255, V2C_962_255, V2C_1022_255, V2C_1100_255, V2C_1145_255, V2C_1406_255, V2C_1407_255, V2C_22_256, V2C_81_256, V2C_120_256, V2C_176_256, V2C_193_256, V2C_247_256, V2C_471_256, V2C_511_256, V2C_547_256, V2C_609_256, V2C_634_256, V2C_680_256, V2C_897_256, V2C_921_256, V2C_1005_256, V2C_1035_256, V2C_1062_256, V2C_1126_256, V2C_1407_256, V2C_1408_256, V2C_41_257, V2C_51_257, V2C_134_257, V2C_157_257, V2C_221_257, V2C_287_257, V2C_336_257, V2C_355_257, V2C_434_257, V2C_716_257, V2C_732_257, V2C_786_257, V2C_912_257, V2C_960_257, V2C_1003_257, V2C_1055_257, V2C_1104_257, V2C_1152_257, V2C_1408_257, V2C_1409_257, V2C_24_258, V2C_96_258, V2C_136_258, V2C_156_258, V2C_238_258, V2C_269_258, V2C_322_258, V2C_474_258, V2C_571_258, V2C_604_258, V2C_808_258, V2C_836_258, V2C_869_258, V2C_931_258, V2C_966_258, V2C_1033_258, V2C_1097_258, V2C_1147_258, V2C_1409_258, V2C_1410_258, V2C_48_259, V2C_84_259, V2C_104_259, V2C_165_259, V2C_227_259, V2C_270_259, V2C_370_259, V2C_424_259, V2C_521_259, V2C_757_259, V2C_805_259, V2C_853_259, V2C_894_259, V2C_935_259, V2C_969_259, V2C_1056_259, V2C_1082_259, V2C_1141_259, V2C_1410_259, V2C_1411_259, V2C_9_260, V2C_58_260, V2C_114_260, V2C_162_260, V2C_239_260, V2C_260_260, V2C_311_260, V2C_418_260, V2C_507_260, V2C_667_260, V2C_680_260, V2C_848_260, V2C_890_260, V2C_953_260, V2C_984_260, V2C_1016_260, V2C_1083_260, V2C_1114_260, V2C_1411_260, V2C_1412_260, V2C_4_261, V2C_79_261, V2C_144_261, V2C_178_261, V2C_196_261, V2C_263_261, V2C_360_261, V2C_415_261, V2C_574_261, V2C_583_261, V2C_659_261, V2C_763_261, V2C_894_261, V2C_938_261, V2C_963_261, V2C_1023_261, V2C_1101_261, V2C_1146_261, V2C_1412_261, V2C_1413_261, V2C_23_262, V2C_82_262, V2C_121_262, V2C_177_262, V2C_194_262, V2C_248_262, V2C_472_262, V2C_512_262, V2C_548_262, V2C_610_262, V2C_635_262, V2C_681_262, V2C_898_262, V2C_922_262, V2C_1006_262, V2C_1036_262, V2C_1063_262, V2C_1127_262, V2C_1413_262, V2C_1414_262, V2C_42_263, V2C_52_263, V2C_135_263, V2C_158_263, V2C_222_263, V2C_288_263, V2C_289_263, V2C_356_263, V2C_435_263, V2C_717_263, V2C_733_263, V2C_787_263, V2C_865_263, V2C_913_263, V2C_1004_263, V2C_1056_263, V2C_1057_263, V2C_1105_263, V2C_1414_263, V2C_1415_263, V2C_25_264, V2C_49_264, V2C_137_264, V2C_157_264, V2C_239_264, V2C_270_264, V2C_323_264, V2C_475_264, V2C_572_264, V2C_605_264, V2C_809_264, V2C_837_264, V2C_870_264, V2C_932_264, V2C_967_264, V2C_1034_264, V2C_1098_264, V2C_1148_264, V2C_1415_264, V2C_1416_264, V2C_1_265, V2C_85_265, V2C_105_265, V2C_166_265, V2C_228_265, V2C_271_265, V2C_371_265, V2C_425_265, V2C_522_265, V2C_758_265, V2C_806_265, V2C_854_265, V2C_895_265, V2C_936_265, V2C_970_265, V2C_1009_265, V2C_1083_265, V2C_1142_265, V2C_1416_265, V2C_1417_265, V2C_10_266, V2C_59_266, V2C_115_266, V2C_163_266, V2C_240_266, V2C_261_266, V2C_312_266, V2C_419_266, V2C_508_266, V2C_668_266, V2C_681_266, V2C_849_266, V2C_891_266, V2C_954_266, V2C_985_266, V2C_1017_266, V2C_1084_266, V2C_1115_266, V2C_1417_266, V2C_1418_266, V2C_5_267, V2C_80_267, V2C_97_267, V2C_179_267, V2C_197_267, V2C_264_267, V2C_361_267, V2C_416_267, V2C_575_267, V2C_584_267, V2C_660_267, V2C_764_267, V2C_895_267, V2C_939_267, V2C_964_267, V2C_1024_267, V2C_1102_267, V2C_1147_267, V2C_1418_267, V2C_1419_267, V2C_24_268, V2C_83_268, V2C_122_268, V2C_178_268, V2C_195_268, V2C_249_268, V2C_473_268, V2C_513_268, V2C_549_268, V2C_611_268, V2C_636_268, V2C_682_268, V2C_899_268, V2C_923_268, V2C_1007_268, V2C_1037_268, V2C_1064_268, V2C_1128_268, V2C_1419_268, V2C_1420_268, V2C_43_269, V2C_53_269, V2C_136_269, V2C_159_269, V2C_223_269, V2C_241_269, V2C_290_269, V2C_357_269, V2C_436_269, V2C_718_269, V2C_734_269, V2C_788_269, V2C_866_269, V2C_914_269, V2C_1005_269, V2C_1009_269, V2C_1058_269, V2C_1106_269, V2C_1420_269, V2C_1421_269, V2C_26_270, V2C_50_270, V2C_138_270, V2C_158_270, V2C_240_270, V2C_271_270, V2C_324_270, V2C_476_270, V2C_573_270, V2C_606_270, V2C_810_270, V2C_838_270, V2C_871_270, V2C_933_270, V2C_968_270, V2C_1035_270, V2C_1099_270, V2C_1149_270, V2C_1421_270, V2C_1422_270, V2C_2_271, V2C_86_271, V2C_106_271, V2C_167_271, V2C_229_271, V2C_272_271, V2C_372_271, V2C_426_271, V2C_523_271, V2C_759_271, V2C_807_271, V2C_855_271, V2C_896_271, V2C_937_271, V2C_971_271, V2C_1010_271, V2C_1084_271, V2C_1143_271, V2C_1422_271, V2C_1423_271, V2C_11_272, V2C_60_272, V2C_116_272, V2C_164_272, V2C_193_272, V2C_262_272, V2C_313_272, V2C_420_272, V2C_509_272, V2C_669_272, V2C_682_272, V2C_850_272, V2C_892_272, V2C_955_272, V2C_986_272, V2C_1018_272, V2C_1085_272, V2C_1116_272, V2C_1423_272, V2C_1424_272, V2C_6_273, V2C_81_273, V2C_98_273, V2C_180_273, V2C_198_273, V2C_265_273, V2C_362_273, V2C_417_273, V2C_576_273, V2C_585_273, V2C_661_273, V2C_765_273, V2C_896_273, V2C_940_273, V2C_965_273, V2C_1025_273, V2C_1103_273, V2C_1148_273, V2C_1424_273, V2C_1425_273, V2C_25_274, V2C_84_274, V2C_123_274, V2C_179_274, V2C_196_274, V2C_250_274, V2C_474_274, V2C_514_274, V2C_550_274, V2C_612_274, V2C_637_274, V2C_683_274, V2C_900_274, V2C_924_274, V2C_1008_274, V2C_1038_274, V2C_1065_274, V2C_1129_274, V2C_1425_274, V2C_1426_274, V2C_44_275, V2C_54_275, V2C_137_275, V2C_160_275, V2C_224_275, V2C_242_275, V2C_291_275, V2C_358_275, V2C_437_275, V2C_719_275, V2C_735_275, V2C_789_275, V2C_867_275, V2C_915_275, V2C_1006_275, V2C_1010_275, V2C_1059_275, V2C_1107_275, V2C_1426_275, V2C_1427_275, V2C_27_276, V2C_51_276, V2C_139_276, V2C_159_276, V2C_193_276, V2C_272_276, V2C_325_276, V2C_477_276, V2C_574_276, V2C_607_276, V2C_811_276, V2C_839_276, V2C_872_276, V2C_934_276, V2C_969_276, V2C_1036_276, V2C_1100_276, V2C_1150_276, V2C_1427_276, V2C_1428_276, V2C_3_277, V2C_87_277, V2C_107_277, V2C_168_277, V2C_230_277, V2C_273_277, V2C_373_277, V2C_427_277, V2C_524_277, V2C_760_277, V2C_808_277, V2C_856_277, V2C_897_277, V2C_938_277, V2C_972_277, V2C_1011_277, V2C_1085_277, V2C_1144_277, V2C_1428_277, V2C_1429_277, V2C_12_278, V2C_61_278, V2C_117_278, V2C_165_278, V2C_194_278, V2C_263_278, V2C_314_278, V2C_421_278, V2C_510_278, V2C_670_278, V2C_683_278, V2C_851_278, V2C_893_278, V2C_956_278, V2C_987_278, V2C_1019_278, V2C_1086_278, V2C_1117_278, V2C_1429_278, V2C_1430_278, V2C_7_279, V2C_82_279, V2C_99_279, V2C_181_279, V2C_199_279, V2C_266_279, V2C_363_279, V2C_418_279, V2C_529_279, V2C_586_279, V2C_662_279, V2C_766_279, V2C_897_279, V2C_941_279, V2C_966_279, V2C_1026_279, V2C_1104_279, V2C_1149_279, V2C_1430_279, V2C_1431_279, V2C_26_280, V2C_85_280, V2C_124_280, V2C_180_280, V2C_197_280, V2C_251_280, V2C_475_280, V2C_515_280, V2C_551_280, V2C_613_280, V2C_638_280, V2C_684_280, V2C_901_280, V2C_925_280, V2C_961_280, V2C_1039_280, V2C_1066_280, V2C_1130_280, V2C_1431_280, V2C_1432_280, V2C_45_281, V2C_55_281, V2C_138_281, V2C_161_281, V2C_225_281, V2C_243_281, V2C_292_281, V2C_359_281, V2C_438_281, V2C_720_281, V2C_736_281, V2C_790_281, V2C_868_281, V2C_916_281, V2C_1007_281, V2C_1011_281, V2C_1060_281, V2C_1108_281, V2C_1432_281, V2C_1433_281, V2C_28_282, V2C_52_282, V2C_140_282, V2C_160_282, V2C_194_282, V2C_273_282, V2C_326_282, V2C_478_282, V2C_575_282, V2C_608_282, V2C_812_282, V2C_840_282, V2C_873_282, V2C_935_282, V2C_970_282, V2C_1037_282, V2C_1101_282, V2C_1151_282, V2C_1433_282, V2C_1434_282, V2C_4_283, V2C_88_283, V2C_108_283, V2C_169_283, V2C_231_283, V2C_274_283, V2C_374_283, V2C_428_283, V2C_525_283, V2C_761_283, V2C_809_283, V2C_857_283, V2C_898_283, V2C_939_283, V2C_973_283, V2C_1012_283, V2C_1086_283, V2C_1145_283, V2C_1434_283, V2C_1435_283, V2C_13_284, V2C_62_284, V2C_118_284, V2C_166_284, V2C_195_284, V2C_264_284, V2C_315_284, V2C_422_284, V2C_511_284, V2C_671_284, V2C_684_284, V2C_852_284, V2C_894_284, V2C_957_284, V2C_988_284, V2C_1020_284, V2C_1087_284, V2C_1118_284, V2C_1435_284, V2C_1436_284, V2C_8_285, V2C_83_285, V2C_100_285, V2C_182_285, V2C_200_285, V2C_267_285, V2C_364_285, V2C_419_285, V2C_530_285, V2C_587_285, V2C_663_285, V2C_767_285, V2C_898_285, V2C_942_285, V2C_967_285, V2C_1027_285, V2C_1057_285, V2C_1150_285, V2C_1436_285, V2C_1437_285, V2C_27_286, V2C_86_286, V2C_125_286, V2C_181_286, V2C_198_286, V2C_252_286, V2C_476_286, V2C_516_286, V2C_552_286, V2C_614_286, V2C_639_286, V2C_685_286, V2C_902_286, V2C_926_286, V2C_962_286, V2C_1040_286, V2C_1067_286, V2C_1131_286, V2C_1437_286, V2C_1438_286, V2C_46_287, V2C_56_287, V2C_139_287, V2C_162_287, V2C_226_287, V2C_244_287, V2C_293_287, V2C_360_287, V2C_439_287, V2C_673_287, V2C_737_287, V2C_791_287, V2C_869_287, V2C_917_287, V2C_1008_287, V2C_1012_287, V2C_1061_287, V2C_1109_287, V2C_1438_287, V2C_1439_287, V2C_29_288, V2C_53_288, V2C_141_288, V2C_161_288, V2C_195_288, V2C_274_288, V2C_327_288, V2C_479_288, V2C_576_288, V2C_609_288, V2C_813_288, V2C_841_288, V2C_874_288, V2C_936_288, V2C_971_288, V2C_1038_288, V2C_1102_288, V2C_1152_288, V2C_1439_288, V2C_1440_288, V2C_0_0;
wire [quan_width - 1:0] V_1, V_2, V_3, V_4, V_5, V_6, V_7, V_8, V_9, V_10, V_11, V_12, V_13, V_14, V_15, V_16, V_17, V_18, V_19, V_20, V_21, V_22, V_23, V_24, V_25, V_26, V_27, V_28, V_29, V_30, V_31, V_32, V_33, V_34, V_35, V_36, V_37, V_38, V_39, V_40, V_41, V_42, V_43, V_44, V_45, V_46, V_47, V_48, V_49, V_50, V_51, V_52, V_53, V_54, V_55, V_56, V_57, V_58, V_59, V_60, V_61, V_62, V_63, V_64, V_65, V_66, V_67, V_68, V_69, V_70, V_71, V_72, V_73, V_74, V_75, V_76, V_77, V_78, V_79, V_80, V_81, V_82, V_83, V_84, V_85, V_86, V_87, V_88, V_89, V_90, V_91, V_92, V_93, V_94, V_95, V_96, V_97, V_98, V_99, V_100, V_101, V_102, V_103, V_104, V_105, V_106, V_107, V_108, V_109, V_110, V_111, V_112, V_113, V_114, V_115, V_116, V_117, V_118, V_119, V_120, V_121, V_122, V_123, V_124, V_125, V_126, V_127, V_128, V_129, V_130, V_131, V_132, V_133, V_134, V_135, V_136, V_137, V_138, V_139, V_140, V_141, V_142, V_143, V_144, V_145, V_146, V_147, V_148, V_149, V_150, V_151, V_152, V_153, V_154, V_155, V_156, V_157, V_158, V_159, V_160, V_161, V_162, V_163, V_164, V_165, V_166, V_167, V_168, V_169, V_170, V_171, V_172, V_173, V_174, V_175, V_176, V_177, V_178, V_179, V_180, V_181, V_182, V_183, V_184, V_185, V_186, V_187, V_188, V_189, V_190, V_191, V_192, V_193, V_194, V_195, V_196, V_197, V_198, V_199, V_200, V_201, V_202, V_203, V_204, V_205, V_206, V_207, V_208, V_209, V_210, V_211, V_212, V_213, V_214, V_215, V_216, V_217, V_218, V_219, V_220, V_221, V_222, V_223, V_224, V_225, V_226, V_227, V_228, V_229, V_230, V_231, V_232, V_233, V_234, V_235, V_236, V_237, V_238, V_239, V_240, V_241, V_242, V_243, V_244, V_245, V_246, V_247, V_248, V_249, V_250, V_251, V_252, V_253, V_254, V_255, V_256, V_257, V_258, V_259, V_260, V_261, V_262, V_263, V_264, V_265, V_266, V_267, V_268, V_269, V_270, V_271, V_272, V_273, V_274, V_275, V_276, V_277, V_278, V_279, V_280, V_281, V_282, V_283, V_284, V_285, V_286, V_287, V_288, V_289, V_290, V_291, V_292, V_293, V_294, V_295, V_296, V_297, V_298, V_299, V_300, V_301, V_302, V_303, V_304, V_305, V_306, V_307, V_308, V_309, V_310, V_311, V_312, V_313, V_314, V_315, V_316, V_317, V_318, V_319, V_320, V_321, V_322, V_323, V_324, V_325, V_326, V_327, V_328, V_329, V_330, V_331, V_332, V_333, V_334, V_335, V_336, V_337, V_338, V_339, V_340, V_341, V_342, V_343, V_344, V_345, V_346, V_347, V_348, V_349, V_350, V_351, V_352, V_353, V_354, V_355, V_356, V_357, V_358, V_359, V_360, V_361, V_362, V_363, V_364, V_365, V_366, V_367, V_368, V_369, V_370, V_371, V_372, V_373, V_374, V_375, V_376, V_377, V_378, V_379, V_380, V_381, V_382, V_383, V_384, V_385, V_386, V_387, V_388, V_389, V_390, V_391, V_392, V_393, V_394, V_395, V_396, V_397, V_398, V_399, V_400, V_401, V_402, V_403, V_404, V_405, V_406, V_407, V_408, V_409, V_410, V_411, V_412, V_413, V_414, V_415, V_416, V_417, V_418, V_419, V_420, V_421, V_422, V_423, V_424, V_425, V_426, V_427, V_428, V_429, V_430, V_431, V_432, V_433, V_434, V_435, V_436, V_437, V_438, V_439, V_440, V_441, V_442, V_443, V_444, V_445, V_446, V_447, V_448, V_449, V_450, V_451, V_452, V_453, V_454, V_455, V_456, V_457, V_458, V_459, V_460, V_461, V_462, V_463, V_464, V_465, V_466, V_467, V_468, V_469, V_470, V_471, V_472, V_473, V_474, V_475, V_476, V_477, V_478, V_479, V_480, V_481, V_482, V_483, V_484, V_485, V_486, V_487, V_488, V_489, V_490, V_491, V_492, V_493, V_494, V_495, V_496, V_497, V_498, V_499, V_500, V_501, V_502, V_503, V_504, V_505, V_506, V_507, V_508, V_509, V_510, V_511, V_512, V_513, V_514, V_515, V_516, V_517, V_518, V_519, V_520, V_521, V_522, V_523, V_524, V_525, V_526, V_527, V_528, V_529, V_530, V_531, V_532, V_533, V_534, V_535, V_536, V_537, V_538, V_539, V_540, V_541, V_542, V_543, V_544, V_545, V_546, V_547, V_548, V_549, V_550, V_551, V_552, V_553, V_554, V_555, V_556, V_557, V_558, V_559, V_560, V_561, V_562, V_563, V_564, V_565, V_566, V_567, V_568, V_569, V_570, V_571, V_572, V_573, V_574, V_575, V_576, V_577, V_578, V_579, V_580, V_581, V_582, V_583, V_584, V_585, V_586, V_587, V_588, V_589, V_590, V_591, V_592, V_593, V_594, V_595, V_596, V_597, V_598, V_599, V_600, V_601, V_602, V_603, V_604, V_605, V_606, V_607, V_608, V_609, V_610, V_611, V_612, V_613, V_614, V_615, V_616, V_617, V_618, V_619, V_620, V_621, V_622, V_623, V_624, V_625, V_626, V_627, V_628, V_629, V_630, V_631, V_632, V_633, V_634, V_635, V_636, V_637, V_638, V_639, V_640, V_641, V_642, V_643, V_644, V_645, V_646, V_647, V_648, V_649, V_650, V_651, V_652, V_653, V_654, V_655, V_656, V_657, V_658, V_659, V_660, V_661, V_662, V_663, V_664, V_665, V_666, V_667, V_668, V_669, V_670, V_671, V_672, V_673, V_674, V_675, V_676, V_677, V_678, V_679, V_680, V_681, V_682, V_683, V_684, V_685, V_686, V_687, V_688, V_689, V_690, V_691, V_692, V_693, V_694, V_695, V_696, V_697, V_698, V_699, V_700, V_701, V_702, V_703, V_704, V_705, V_706, V_707, V_708, V_709, V_710, V_711, V_712, V_713, V_714, V_715, V_716, V_717, V_718, V_719, V_720, V_721, V_722, V_723, V_724, V_725, V_726, V_727, V_728, V_729, V_730, V_731, V_732, V_733, V_734, V_735, V_736, V_737, V_738, V_739, V_740, V_741, V_742, V_743, V_744, V_745, V_746, V_747, V_748, V_749, V_750, V_751, V_752, V_753, V_754, V_755, V_756, V_757, V_758, V_759, V_760, V_761, V_762, V_763, V_764, V_765, V_766, V_767, V_768, V_769, V_770, V_771, V_772, V_773, V_774, V_775, V_776, V_777, V_778, V_779, V_780, V_781, V_782, V_783, V_784, V_785, V_786, V_787, V_788, V_789, V_790, V_791, V_792, V_793, V_794, V_795, V_796, V_797, V_798, V_799, V_800, V_801, V_802, V_803, V_804, V_805, V_806, V_807, V_808, V_809, V_810, V_811, V_812, V_813, V_814, V_815, V_816, V_817, V_818, V_819, V_820, V_821, V_822, V_823, V_824, V_825, V_826, V_827, V_828, V_829, V_830, V_831, V_832, V_833, V_834, V_835, V_836, V_837, V_838, V_839, V_840, V_841, V_842, V_843, V_844, V_845, V_846, V_847, V_848, V_849, V_850, V_851, V_852, V_853, V_854, V_855, V_856, V_857, V_858, V_859, V_860, V_861, V_862, V_863, V_864, V_865, V_866, V_867, V_868, V_869, V_870, V_871, V_872, V_873, V_874, V_875, V_876, V_877, V_878, V_879, V_880, V_881, V_882, V_883, V_884, V_885, V_886, V_887, V_888, V_889, V_890, V_891, V_892, V_893, V_894, V_895, V_896, V_897, V_898, V_899, V_900, V_901, V_902, V_903, V_904, V_905, V_906, V_907, V_908, V_909, V_910, V_911, V_912, V_913, V_914, V_915, V_916, V_917, V_918, V_919, V_920, V_921, V_922, V_923, V_924, V_925, V_926, V_927, V_928, V_929, V_930, V_931, V_932, V_933, V_934, V_935, V_936, V_937, V_938, V_939, V_940, V_941, V_942, V_943, V_944, V_945, V_946, V_947, V_948, V_949, V_950, V_951, V_952, V_953, V_954, V_955, V_956, V_957, V_958, V_959, V_960, V_961, V_962, V_963, V_964, V_965, V_966, V_967, V_968, V_969, V_970, V_971, V_972, V_973, V_974, V_975, V_976, V_977, V_978, V_979, V_980, V_981, V_982, V_983, V_984, V_985, V_986, V_987, V_988, V_989, V_990, V_991, V_992, V_993, V_994, V_995, V_996, V_997, V_998, V_999, V_1000, V_1001, V_1002, V_1003, V_1004, V_1005, V_1006, V_1007, V_1008, V_1009, V_1010, V_1011, V_1012, V_1013, V_1014, V_1015, V_1016, V_1017, V_1018, V_1019, V_1020, V_1021, V_1022, V_1023, V_1024, V_1025, V_1026, V_1027, V_1028, V_1029, V_1030, V_1031, V_1032, V_1033, V_1034, V_1035, V_1036, V_1037, V_1038, V_1039, V_1040, V_1041, V_1042, V_1043, V_1044, V_1045, V_1046, V_1047, V_1048, V_1049, V_1050, V_1051, V_1052, V_1053, V_1054, V_1055, V_1056, V_1057, V_1058, V_1059, V_1060, V_1061, V_1062, V_1063, V_1064, V_1065, V_1066, V_1067, V_1068, V_1069, V_1070, V_1071, V_1072, V_1073, V_1074, V_1075, V_1076, V_1077, V_1078, V_1079, V_1080, V_1081, V_1082, V_1083, V_1084, V_1085, V_1086, V_1087, V_1088, V_1089, V_1090, V_1091, V_1092, V_1093, V_1094, V_1095, V_1096, V_1097, V_1098, V_1099, V_1100, V_1101, V_1102, V_1103, V_1104, V_1105, V_1106, V_1107, V_1108, V_1109, V_1110, V_1111, V_1112, V_1113, V_1114, V_1115, V_1116, V_1117, V_1118, V_1119, V_1120, V_1121, V_1122, V_1123, V_1124, V_1125, V_1126, V_1127, V_1128, V_1129, V_1130, V_1131, V_1132, V_1133, V_1134, V_1135, V_1136, V_1137, V_1138, V_1139, V_1140, V_1141, V_1142, V_1143, V_1144, V_1145, V_1146, V_1147, V_1148, V_1149, V_1150, V_1151, V_1152, V_1153, V_1154, V_1155, V_1156, V_1157, V_1158, V_1159, V_1160, V_1161, V_1162, V_1163, V_1164, V_1165, V_1166, V_1167, V_1168, V_1169, V_1170, V_1171, V_1172, V_1173, V_1174, V_1175, V_1176, V_1177, V_1178, V_1179, V_1180, V_1181, V_1182, V_1183, V_1184, V_1185, V_1186, V_1187, V_1188, V_1189, V_1190, V_1191, V_1192, V_1193, V_1194, V_1195, V_1196, V_1197, V_1198, V_1199, V_1200, V_1201, V_1202, V_1203, V_1204, V_1205, V_1206, V_1207, V_1208, V_1209, V_1210, V_1211, V_1212, V_1213, V_1214, V_1215, V_1216, V_1217, V_1218, V_1219, V_1220, V_1221, V_1222, V_1223, V_1224, V_1225, V_1226, V_1227, V_1228, V_1229, V_1230, V_1231, V_1232, V_1233, V_1234, V_1235, V_1236, V_1237, V_1238, V_1239, V_1240, V_1241, V_1242, V_1243, V_1244, V_1245, V_1246, V_1247, V_1248, V_1249, V_1250, V_1251, V_1252, V_1253, V_1254, V_1255, V_1256, V_1257, V_1258, V_1259, V_1260, V_1261, V_1262, V_1263, V_1264, V_1265, V_1266, V_1267, V_1268, V_1269, V_1270, V_1271, V_1272, V_1273, V_1274, V_1275, V_1276, V_1277, V_1278, V_1279, V_1280, V_1281, V_1282, V_1283, V_1284, V_1285, V_1286, V_1287, V_1288, V_1289, V_1290, V_1291, V_1292, V_1293, V_1294, V_1295, V_1296, V_1297, V_1298, V_1299, V_1300, V_1301, V_1302, V_1303, V_1304, V_1305, V_1306, V_1307, V_1308, V_1309, V_1310, V_1311, V_1312, V_1313, V_1314, V_1315, V_1316, V_1317, V_1318, V_1319, V_1320, V_1321, V_1322, V_1323, V_1324, V_1325, V_1326, V_1327, V_1328, V_1329, V_1330, V_1331, V_1332, V_1333, V_1334, V_1335, V_1336, V_1337, V_1338, V_1339, V_1340, V_1341, V_1342, V_1343, V_1344, V_1345, V_1346, V_1347, V_1348, V_1349, V_1350, V_1351, V_1352, V_1353, V_1354, V_1355, V_1356, V_1357, V_1358, V_1359, V_1360, V_1361, V_1362, V_1363, V_1364, V_1365, V_1366, V_1367, V_1368, V_1369, V_1370, V_1371, V_1372, V_1373, V_1374, V_1375, V_1376, V_1377, V_1378, V_1379, V_1380, V_1381, V_1382, V_1383, V_1384, V_1385, V_1386, V_1387, V_1388, V_1389, V_1390, V_1391, V_1392, V_1393, V_1394, V_1395, V_1396, V_1397, V_1398, V_1399, V_1400, V_1401, V_1402, V_1403, V_1404, V_1405, V_1406, V_1407, V_1408, V_1409, V_1410, V_1411, V_1412, V_1413, V_1414, V_1415, V_1416, V_1417, V_1418, V_1419, V_1420, V_1421, V_1422, V_1423, V_1424, V_1425, V_1426, V_1427, V_1428, V_1429, V_1430, V_1431, V_1432, V_1433, V_1434, V_1435, V_1436, V_1437, V_1438, V_1439, V_1440;

always @ (posedge clk or negedge rst) begin
if (rst && in_valid == 1) begin
	L [(in_index + 4)*quan_width-1-:4*quan_width] <= data_in;
	cnt <= 0;
end
if (rst && in_valid == 0 && cnt == 0) 
cnt <= 1;
end


always @ (posedge clk or negedge rst) begin
if (rst && out_valid == 1)
data_out <= Bit [out_index+3-:4];

if (rst && out_valid == 1) begin
if (out_index < code_length - 4)
out_index <= out_index + 4;
else begin
out_valid <= 0;
end
end
end

always @ (posedge clk or negedge rst) begin
	if (!rst) begin
		cnt <= 0;
		iter <= 0;
		out_valid <= 0;
		out_index <= 0;
		data_out <= 4'd0;
		Check_1 <= 1;
		Check_2 <= 1;
		Check_3 <= 1;
		Check_4 <= 1;
		Check_5 <= 1;
		Check_6 <= 1;
		Check_7 <= 1;
		Check_8 <= 1;
		Check_9 <= 1;
		Check_10 <= 1;
		Check_11 <= 1;
		Check_12 <= 1;
		Check_13 <= 1;
		Check_14 <= 1;
		Check_15 <= 1;
		Check_16 <= 1;
		Check_17 <= 1;
		Check_18 <= 1;
		Check_19 <= 1;
		Check_20 <= 1;
		Check_21 <= 1;
		Check_22 <= 1;
		Check_23 <= 1;
		Check_24 <= 1;
		Check_25 <= 1;
		Check_26 <= 1;
		Check_27 <= 1;
		Check_28 <= 1;
		Check_29 <= 1;
		Check_30 <= 1;
		Check_31 <= 1;
		Check_32 <= 1;
		Check_33 <= 1;
		Check_34 <= 1;
		Check_35 <= 1;
		Check_36 <= 1;
		Check_37 <= 1;
		Check_38 <= 1;
		Check_39 <= 1;
		Check_40 <= 1;
		Check_41 <= 1;
		Check_42 <= 1;
		Check_43 <= 1;
		Check_44 <= 1;
		Check_45 <= 1;
		Check_46 <= 1;
		Check_47 <= 1;
		Check_48 <= 1;
		Check_49 <= 1;
		Check_50 <= 1;
		Check_51 <= 1;
		Check_52 <= 1;
		Check_53 <= 1;
		Check_54 <= 1;
		Check_55 <= 1;
		Check_56 <= 1;
		Check_57 <= 1;
		Check_58 <= 1;
		Check_59 <= 1;
		Check_60 <= 1;
		Check_61 <= 1;
		Check_62 <= 1;
		Check_63 <= 1;
		Check_64 <= 1;
		Check_65 <= 1;
		Check_66 <= 1;
		Check_67 <= 1;
		Check_68 <= 1;
		Check_69 <= 1;
		Check_70 <= 1;
		Check_71 <= 1;
		Check_72 <= 1;
		Check_73 <= 1;
		Check_74 <= 1;
		Check_75 <= 1;
		Check_76 <= 1;
		Check_77 <= 1;
		Check_78 <= 1;
		Check_79 <= 1;
		Check_80 <= 1;
		Check_81 <= 1;
		Check_82 <= 1;
		Check_83 <= 1;
		Check_84 <= 1;
		Check_85 <= 1;
		Check_86 <= 1;
		Check_87 <= 1;
		Check_88 <= 1;
		Check_89 <= 1;
		Check_90 <= 1;
		Check_91 <= 1;
		Check_92 <= 1;
		Check_93 <= 1;
		Check_94 <= 1;
		Check_95 <= 1;
		Check_96 <= 1;
		Check_97 <= 1;
		Check_98 <= 1;
		Check_99 <= 1;
		Check_100 <= 1;
		Check_101 <= 1;
		Check_102 <= 1;
		Check_103 <= 1;
		Check_104 <= 1;
		Check_105 <= 1;
		Check_106 <= 1;
		Check_107 <= 1;
		Check_108 <= 1;
		Check_109 <= 1;
		Check_110 <= 1;
		Check_111 <= 1;
		Check_112 <= 1;
		Check_113 <= 1;
		Check_114 <= 1;
		Check_115 <= 1;
		Check_116 <= 1;
		Check_117 <= 1;
		Check_118 <= 1;
		Check_119 <= 1;
		Check_120 <= 1;
		Check_121 <= 1;
		Check_122 <= 1;
		Check_123 <= 1;
		Check_124 <= 1;
		Check_125 <= 1;
		Check_126 <= 1;
		Check_127 <= 1;
		Check_128 <= 1;
		Check_129 <= 1;
		Check_130 <= 1;
		Check_131 <= 1;
		Check_132 <= 1;
		Check_133 <= 1;
		Check_134 <= 1;
		Check_135 <= 1;
		Check_136 <= 1;
		Check_137 <= 1;
		Check_138 <= 1;
		Check_139 <= 1;
		Check_140 <= 1;
		Check_141 <= 1;
		Check_142 <= 1;
		Check_143 <= 1;
		Check_144 <= 1;
		Check_145 <= 1;
		Check_146 <= 1;
		Check_147 <= 1;
		Check_148 <= 1;
		Check_149 <= 1;
		Check_150 <= 1;
		Check_151 <= 1;
		Check_152 <= 1;
		Check_153 <= 1;
		Check_154 <= 1;
		Check_155 <= 1;
		Check_156 <= 1;
		Check_157 <= 1;
		Check_158 <= 1;
		Check_159 <= 1;
		Check_160 <= 1;
		Check_161 <= 1;
		Check_162 <= 1;
		Check_163 <= 1;
		Check_164 <= 1;
		Check_165 <= 1;
		Check_166 <= 1;
		Check_167 <= 1;
		Check_168 <= 1;
		Check_169 <= 1;
		Check_170 <= 1;
		Check_171 <= 1;
		Check_172 <= 1;
		Check_173 <= 1;
		Check_174 <= 1;
		Check_175 <= 1;
		Check_176 <= 1;
		Check_177 <= 1;
		Check_178 <= 1;
		Check_179 <= 1;
		Check_180 <= 1;
		Check_181 <= 1;
		Check_182 <= 1;
		Check_183 <= 1;
		Check_184 <= 1;
		Check_185 <= 1;
		Check_186 <= 1;
		Check_187 <= 1;
		Check_188 <= 1;
		Check_189 <= 1;
		Check_190 <= 1;
		Check_191 <= 1;
		Check_192 <= 1;
		Check_193 <= 1;
		Check_194 <= 1;
		Check_195 <= 1;
		Check_196 <= 1;
		Check_197 <= 1;
		Check_198 <= 1;
		Check_199 <= 1;
		Check_200 <= 1;
		Check_201 <= 1;
		Check_202 <= 1;
		Check_203 <= 1;
		Check_204 <= 1;
		Check_205 <= 1;
		Check_206 <= 1;
		Check_207 <= 1;
		Check_208 <= 1;
		Check_209 <= 1;
		Check_210 <= 1;
		Check_211 <= 1;
		Check_212 <= 1;
		Check_213 <= 1;
		Check_214 <= 1;
		Check_215 <= 1;
		Check_216 <= 1;
		Check_217 <= 1;
		Check_218 <= 1;
		Check_219 <= 1;
		Check_220 <= 1;
		Check_221 <= 1;
		Check_222 <= 1;
		Check_223 <= 1;
		Check_224 <= 1;
		Check_225 <= 1;
		Check_226 <= 1;
		Check_227 <= 1;
		Check_228 <= 1;
		Check_229 <= 1;
		Check_230 <= 1;
		Check_231 <= 1;
		Check_232 <= 1;
		Check_233 <= 1;
		Check_234 <= 1;
		Check_235 <= 1;
		Check_236 <= 1;
		Check_237 <= 1;
		Check_238 <= 1;
		Check_239 <= 1;
		Check_240 <= 1;
		Check_241 <= 1;
		Check_242 <= 1;
		Check_243 <= 1;
		Check_244 <= 1;
		Check_245 <= 1;
		Check_246 <= 1;
		Check_247 <= 1;
		Check_248 <= 1;
		Check_249 <= 1;
		Check_250 <= 1;
		Check_251 <= 1;
		Check_252 <= 1;
		Check_253 <= 1;
		Check_254 <= 1;
		Check_255 <= 1;
		Check_256 <= 1;
		Check_257 <= 1;
		Check_258 <= 1;
		Check_259 <= 1;
		Check_260 <= 1;
		Check_261 <= 1;
		Check_262 <= 1;
		Check_263 <= 1;
		Check_264 <= 1;
		Check_265 <= 1;
		Check_266 <= 1;
		Check_267 <= 1;
		Check_268 <= 1;
		Check_269 <= 1;
		Check_270 <= 1;
		Check_271 <= 1;
		Check_272 <= 1;
		Check_273 <= 1;
		Check_274 <= 1;
		Check_275 <= 1;
		Check_276 <= 1;
		Check_277 <= 1;
		Check_278 <= 1;
		Check_279 <= 1;
		Check_280 <= 1;
		Check_281 <= 1;
		Check_282 <= 1;
		Check_283 <= 1;
		Check_284 <= 1;
		Check_285 <= 1;
		Check_286 <= 1;
		Check_287 <= 1;
		Check_288 <= 1;
		Check_Sum <= 1;
	end
	else begin
		if (out_valid == 0) begin
			if (8'd0 < cnt && cnt < 8'd15)
			cnt <= cnt + 1;
			else if (cnt == 8'd15) begin
				Check_1 <= Bit[4] ^ Bit[88] ^ Bit[108] ^ Bit[169] ^ Bit[231] ^ Bit[274] ^ Bit[374] ^ Bit[428] ^ Bit[525] ^ Bit[761] ^ Bit[809] ^ Bit[857] ^ Bit[898] ^ Bit[939] ^ Bit[973] ^ Bit[1012] ^ Bit[1086] ^ Bit[1145] ^ Bit[1152];
				Check_2 <= Bit[13] ^ Bit[62] ^ Bit[118] ^ Bit[166] ^ Bit[195] ^ Bit[264] ^ Bit[315] ^ Bit[422] ^ Bit[511] ^ Bit[671] ^ Bit[684] ^ Bit[852] ^ Bit[894] ^ Bit[957] ^ Bit[988] ^ Bit[1020] ^ Bit[1087] ^ Bit[1118] ^ Bit[1152] ^ Bit[1153];
				Check_3 <= Bit[8] ^ Bit[83] ^ Bit[100] ^ Bit[182] ^ Bit[200] ^ Bit[267] ^ Bit[364] ^ Bit[419] ^ Bit[530] ^ Bit[587] ^ Bit[663] ^ Bit[767] ^ Bit[898] ^ Bit[942] ^ Bit[967] ^ Bit[1027] ^ Bit[1057] ^ Bit[1150] ^ Bit[1153] ^ Bit[1154];
				Check_4 <= Bit[27] ^ Bit[86] ^ Bit[125] ^ Bit[181] ^ Bit[198] ^ Bit[252] ^ Bit[476] ^ Bit[516] ^ Bit[552] ^ Bit[614] ^ Bit[639] ^ Bit[685] ^ Bit[902] ^ Bit[926] ^ Bit[962] ^ Bit[1040] ^ Bit[1067] ^ Bit[1131] ^ Bit[1154] ^ Bit[1155];
				Check_5 <= Bit[46] ^ Bit[56] ^ Bit[139] ^ Bit[162] ^ Bit[226] ^ Bit[244] ^ Bit[293] ^ Bit[360] ^ Bit[439] ^ Bit[673] ^ Bit[737] ^ Bit[791] ^ Bit[869] ^ Bit[917] ^ Bit[960] ^ Bit[1012] ^ Bit[1061] ^ Bit[1109] ^ Bit[1155] ^ Bit[1156];
				Check_6 <= Bit[29] ^ Bit[53] ^ Bit[141] ^ Bit[161] ^ Bit[195] ^ Bit[274] ^ Bit[327] ^ Bit[479] ^ Bit[528] ^ Bit[609] ^ Bit[813] ^ Bit[841] ^ Bit[874] ^ Bit[936] ^ Bit[971] ^ Bit[1038] ^ Bit[1102] ^ Bit[1104] ^ Bit[1156] ^ Bit[1157];
				Check_7 <= Bit[5] ^ Bit[89] ^ Bit[109] ^ Bit[170] ^ Bit[232] ^ Bit[275] ^ Bit[375] ^ Bit[429] ^ Bit[526] ^ Bit[762] ^ Bit[810] ^ Bit[858] ^ Bit[899] ^ Bit[940] ^ Bit[974] ^ Bit[1013] ^ Bit[1087] ^ Bit[1146] ^ Bit[1157] ^ Bit[1158];
				Check_8 <= Bit[14] ^ Bit[63] ^ Bit[119] ^ Bit[167] ^ Bit[196] ^ Bit[265] ^ Bit[316] ^ Bit[423] ^ Bit[512] ^ Bit[624] ^ Bit[685] ^ Bit[853] ^ Bit[895] ^ Bit[958] ^ Bit[989] ^ Bit[1021] ^ Bit[1088] ^ Bit[1119] ^ Bit[1158] ^ Bit[1159];
				Check_9 <= Bit[9] ^ Bit[84] ^ Bit[101] ^ Bit[183] ^ Bit[201] ^ Bit[268] ^ Bit[365] ^ Bit[420] ^ Bit[531] ^ Bit[588] ^ Bit[664] ^ Bit[720] ^ Bit[899] ^ Bit[943] ^ Bit[968] ^ Bit[1028] ^ Bit[1058] ^ Bit[1151] ^ Bit[1159] ^ Bit[1160];
				Check_10 <= Bit[28] ^ Bit[87] ^ Bit[126] ^ Bit[182] ^ Bit[199] ^ Bit[253] ^ Bit[477] ^ Bit[517] ^ Bit[553] ^ Bit[615] ^ Bit[640] ^ Bit[686] ^ Bit[903] ^ Bit[927] ^ Bit[963] ^ Bit[1041] ^ Bit[1068] ^ Bit[1132] ^ Bit[1160] ^ Bit[1161];
				Check_11 <= Bit[47] ^ Bit[57] ^ Bit[140] ^ Bit[163] ^ Bit[227] ^ Bit[245] ^ Bit[294] ^ Bit[361] ^ Bit[440] ^ Bit[674] ^ Bit[738] ^ Bit[792] ^ Bit[870] ^ Bit[918] ^ Bit[961] ^ Bit[1013] ^ Bit[1062] ^ Bit[1110] ^ Bit[1161] ^ Bit[1162];
				Check_12 <= Bit[30] ^ Bit[54] ^ Bit[142] ^ Bit[162] ^ Bit[196] ^ Bit[275] ^ Bit[328] ^ Bit[432] ^ Bit[529] ^ Bit[610] ^ Bit[814] ^ Bit[842] ^ Bit[875] ^ Bit[937] ^ Bit[972] ^ Bit[1039] ^ Bit[1103] ^ Bit[1105] ^ Bit[1162] ^ Bit[1163];
				Check_13 <= Bit[6] ^ Bit[90] ^ Bit[110] ^ Bit[171] ^ Bit[233] ^ Bit[276] ^ Bit[376] ^ Bit[430] ^ Bit[527] ^ Bit[763] ^ Bit[811] ^ Bit[859] ^ Bit[900] ^ Bit[941] ^ Bit[975] ^ Bit[1014] ^ Bit[1088] ^ Bit[1147] ^ Bit[1163] ^ Bit[1164];
				Check_14 <= Bit[15] ^ Bit[64] ^ Bit[120] ^ Bit[168] ^ Bit[197] ^ Bit[266] ^ Bit[317] ^ Bit[424] ^ Bit[513] ^ Bit[625] ^ Bit[686] ^ Bit[854] ^ Bit[896] ^ Bit[959] ^ Bit[990] ^ Bit[1022] ^ Bit[1089] ^ Bit[1120] ^ Bit[1164] ^ Bit[1165];
				Check_15 <= Bit[10] ^ Bit[85] ^ Bit[102] ^ Bit[184] ^ Bit[202] ^ Bit[269] ^ Bit[366] ^ Bit[421] ^ Bit[532] ^ Bit[589] ^ Bit[665] ^ Bit[721] ^ Bit[900] ^ Bit[944] ^ Bit[969] ^ Bit[1029] ^ Bit[1059] ^ Bit[1104] ^ Bit[1165] ^ Bit[1166];
				Check_16 <= Bit[29] ^ Bit[88] ^ Bit[127] ^ Bit[183] ^ Bit[200] ^ Bit[254] ^ Bit[478] ^ Bit[518] ^ Bit[554] ^ Bit[616] ^ Bit[641] ^ Bit[687] ^ Bit[904] ^ Bit[928] ^ Bit[964] ^ Bit[1042] ^ Bit[1069] ^ Bit[1133] ^ Bit[1166] ^ Bit[1167];
				Check_17 <= Bit[0] ^ Bit[58] ^ Bit[141] ^ Bit[164] ^ Bit[228] ^ Bit[246] ^ Bit[295] ^ Bit[362] ^ Bit[441] ^ Bit[675] ^ Bit[739] ^ Bit[793] ^ Bit[871] ^ Bit[919] ^ Bit[962] ^ Bit[1014] ^ Bit[1063] ^ Bit[1111] ^ Bit[1167] ^ Bit[1168];
				Check_18 <= Bit[31] ^ Bit[55] ^ Bit[143] ^ Bit[163] ^ Bit[197] ^ Bit[276] ^ Bit[329] ^ Bit[433] ^ Bit[530] ^ Bit[611] ^ Bit[815] ^ Bit[843] ^ Bit[876] ^ Bit[938] ^ Bit[973] ^ Bit[1040] ^ Bit[1056] ^ Bit[1106] ^ Bit[1168] ^ Bit[1169];
				Check_19 <= Bit[7] ^ Bit[91] ^ Bit[111] ^ Bit[172] ^ Bit[234] ^ Bit[277] ^ Bit[377] ^ Bit[431] ^ Bit[480] ^ Bit[764] ^ Bit[812] ^ Bit[860] ^ Bit[901] ^ Bit[942] ^ Bit[976] ^ Bit[1015] ^ Bit[1089] ^ Bit[1148] ^ Bit[1169] ^ Bit[1170];
				Check_20 <= Bit[16] ^ Bit[65] ^ Bit[121] ^ Bit[169] ^ Bit[198] ^ Bit[267] ^ Bit[318] ^ Bit[425] ^ Bit[514] ^ Bit[626] ^ Bit[687] ^ Bit[855] ^ Bit[897] ^ Bit[912] ^ Bit[991] ^ Bit[1023] ^ Bit[1090] ^ Bit[1121] ^ Bit[1170] ^ Bit[1171];
				Check_21 <= Bit[11] ^ Bit[86] ^ Bit[103] ^ Bit[185] ^ Bit[203] ^ Bit[270] ^ Bit[367] ^ Bit[422] ^ Bit[533] ^ Bit[590] ^ Bit[666] ^ Bit[722] ^ Bit[901] ^ Bit[945] ^ Bit[970] ^ Bit[1030] ^ Bit[1060] ^ Bit[1105] ^ Bit[1171] ^ Bit[1172];
				Check_22 <= Bit[30] ^ Bit[89] ^ Bit[128] ^ Bit[184] ^ Bit[201] ^ Bit[255] ^ Bit[479] ^ Bit[519] ^ Bit[555] ^ Bit[617] ^ Bit[642] ^ Bit[688] ^ Bit[905] ^ Bit[929] ^ Bit[965] ^ Bit[1043] ^ Bit[1070] ^ Bit[1134] ^ Bit[1172] ^ Bit[1173];
				Check_23 <= Bit[1] ^ Bit[59] ^ Bit[142] ^ Bit[165] ^ Bit[229] ^ Bit[247] ^ Bit[296] ^ Bit[363] ^ Bit[442] ^ Bit[676] ^ Bit[740] ^ Bit[794] ^ Bit[872] ^ Bit[920] ^ Bit[963] ^ Bit[1015] ^ Bit[1064] ^ Bit[1112] ^ Bit[1173] ^ Bit[1174];
				Check_24 <= Bit[32] ^ Bit[56] ^ Bit[96] ^ Bit[164] ^ Bit[198] ^ Bit[277] ^ Bit[330] ^ Bit[434] ^ Bit[531] ^ Bit[612] ^ Bit[768] ^ Bit[844] ^ Bit[877] ^ Bit[939] ^ Bit[974] ^ Bit[1041] ^ Bit[1057] ^ Bit[1107] ^ Bit[1174] ^ Bit[1175];
				Check_25 <= Bit[8] ^ Bit[92] ^ Bit[112] ^ Bit[173] ^ Bit[235] ^ Bit[278] ^ Bit[378] ^ Bit[384] ^ Bit[481] ^ Bit[765] ^ Bit[813] ^ Bit[861] ^ Bit[902] ^ Bit[943] ^ Bit[977] ^ Bit[1016] ^ Bit[1090] ^ Bit[1149] ^ Bit[1175] ^ Bit[1176];
				Check_26 <= Bit[17] ^ Bit[66] ^ Bit[122] ^ Bit[170] ^ Bit[199] ^ Bit[268] ^ Bit[319] ^ Bit[426] ^ Bit[515] ^ Bit[627] ^ Bit[688] ^ Bit[856] ^ Bit[898] ^ Bit[913] ^ Bit[992] ^ Bit[1024] ^ Bit[1091] ^ Bit[1122] ^ Bit[1176] ^ Bit[1177];
				Check_27 <= Bit[12] ^ Bit[87] ^ Bit[104] ^ Bit[186] ^ Bit[204] ^ Bit[271] ^ Bit[368] ^ Bit[423] ^ Bit[534] ^ Bit[591] ^ Bit[667] ^ Bit[723] ^ Bit[902] ^ Bit[946] ^ Bit[971] ^ Bit[1031] ^ Bit[1061] ^ Bit[1106] ^ Bit[1177] ^ Bit[1178];
				Check_28 <= Bit[31] ^ Bit[90] ^ Bit[129] ^ Bit[185] ^ Bit[202] ^ Bit[256] ^ Bit[432] ^ Bit[520] ^ Bit[556] ^ Bit[618] ^ Bit[643] ^ Bit[689] ^ Bit[906] ^ Bit[930] ^ Bit[966] ^ Bit[1044] ^ Bit[1071] ^ Bit[1135] ^ Bit[1178] ^ Bit[1179];
				Check_29 <= Bit[2] ^ Bit[60] ^ Bit[143] ^ Bit[166] ^ Bit[230] ^ Bit[248] ^ Bit[297] ^ Bit[364] ^ Bit[443] ^ Bit[677] ^ Bit[741] ^ Bit[795] ^ Bit[873] ^ Bit[921] ^ Bit[964] ^ Bit[1016] ^ Bit[1065] ^ Bit[1113] ^ Bit[1179] ^ Bit[1180];
				Check_30 <= Bit[33] ^ Bit[57] ^ Bit[97] ^ Bit[165] ^ Bit[199] ^ Bit[278] ^ Bit[331] ^ Bit[435] ^ Bit[532] ^ Bit[613] ^ Bit[769] ^ Bit[845] ^ Bit[878] ^ Bit[940] ^ Bit[975] ^ Bit[1042] ^ Bit[1058] ^ Bit[1108] ^ Bit[1180] ^ Bit[1181];
				Check_31 <= Bit[9] ^ Bit[93] ^ Bit[113] ^ Bit[174] ^ Bit[236] ^ Bit[279] ^ Bit[379] ^ Bit[385] ^ Bit[482] ^ Bit[766] ^ Bit[814] ^ Bit[862] ^ Bit[903] ^ Bit[944] ^ Bit[978] ^ Bit[1017] ^ Bit[1091] ^ Bit[1150] ^ Bit[1181] ^ Bit[1182];
				Check_32 <= Bit[18] ^ Bit[67] ^ Bit[123] ^ Bit[171] ^ Bit[200] ^ Bit[269] ^ Bit[320] ^ Bit[427] ^ Bit[516] ^ Bit[628] ^ Bit[689] ^ Bit[857] ^ Bit[899] ^ Bit[914] ^ Bit[993] ^ Bit[1025] ^ Bit[1092] ^ Bit[1123] ^ Bit[1182] ^ Bit[1183];
				Check_33 <= Bit[13] ^ Bit[88] ^ Bit[105] ^ Bit[187] ^ Bit[205] ^ Bit[272] ^ Bit[369] ^ Bit[424] ^ Bit[535] ^ Bit[592] ^ Bit[668] ^ Bit[724] ^ Bit[903] ^ Bit[947] ^ Bit[972] ^ Bit[1032] ^ Bit[1062] ^ Bit[1107] ^ Bit[1183] ^ Bit[1184];
				Check_34 <= Bit[32] ^ Bit[91] ^ Bit[130] ^ Bit[186] ^ Bit[203] ^ Bit[257] ^ Bit[433] ^ Bit[521] ^ Bit[557] ^ Bit[619] ^ Bit[644] ^ Bit[690] ^ Bit[907] ^ Bit[931] ^ Bit[967] ^ Bit[1045] ^ Bit[1072] ^ Bit[1136] ^ Bit[1184] ^ Bit[1185];
				Check_35 <= Bit[3] ^ Bit[61] ^ Bit[96] ^ Bit[167] ^ Bit[231] ^ Bit[249] ^ Bit[298] ^ Bit[365] ^ Bit[444] ^ Bit[678] ^ Bit[742] ^ Bit[796] ^ Bit[874] ^ Bit[922] ^ Bit[965] ^ Bit[1017] ^ Bit[1066] ^ Bit[1114] ^ Bit[1185] ^ Bit[1186];
				Check_36 <= Bit[34] ^ Bit[58] ^ Bit[98] ^ Bit[166] ^ Bit[200] ^ Bit[279] ^ Bit[332] ^ Bit[436] ^ Bit[533] ^ Bit[614] ^ Bit[770] ^ Bit[846] ^ Bit[879] ^ Bit[941] ^ Bit[976] ^ Bit[1043] ^ Bit[1059] ^ Bit[1109] ^ Bit[1186] ^ Bit[1187];
				Check_37 <= Bit[10] ^ Bit[94] ^ Bit[114] ^ Bit[175] ^ Bit[237] ^ Bit[280] ^ Bit[380] ^ Bit[386] ^ Bit[483] ^ Bit[767] ^ Bit[815] ^ Bit[863] ^ Bit[904] ^ Bit[945] ^ Bit[979] ^ Bit[1018] ^ Bit[1092] ^ Bit[1151] ^ Bit[1187] ^ Bit[1188];
				Check_38 <= Bit[19] ^ Bit[68] ^ Bit[124] ^ Bit[172] ^ Bit[201] ^ Bit[270] ^ Bit[321] ^ Bit[428] ^ Bit[517] ^ Bit[629] ^ Bit[690] ^ Bit[858] ^ Bit[900] ^ Bit[915] ^ Bit[994] ^ Bit[1026] ^ Bit[1093] ^ Bit[1124] ^ Bit[1188] ^ Bit[1189];
				Check_39 <= Bit[14] ^ Bit[89] ^ Bit[106] ^ Bit[188] ^ Bit[206] ^ Bit[273] ^ Bit[370] ^ Bit[425] ^ Bit[536] ^ Bit[593] ^ Bit[669] ^ Bit[725] ^ Bit[904] ^ Bit[948] ^ Bit[973] ^ Bit[1033] ^ Bit[1063] ^ Bit[1108] ^ Bit[1189] ^ Bit[1190];
				Check_40 <= Bit[33] ^ Bit[92] ^ Bit[131] ^ Bit[187] ^ Bit[204] ^ Bit[258] ^ Bit[434] ^ Bit[522] ^ Bit[558] ^ Bit[620] ^ Bit[645] ^ Bit[691] ^ Bit[908] ^ Bit[932] ^ Bit[968] ^ Bit[1046] ^ Bit[1073] ^ Bit[1137] ^ Bit[1190] ^ Bit[1191];
				Check_41 <= Bit[4] ^ Bit[62] ^ Bit[97] ^ Bit[168] ^ Bit[232] ^ Bit[250] ^ Bit[299] ^ Bit[366] ^ Bit[445] ^ Bit[679] ^ Bit[743] ^ Bit[797] ^ Bit[875] ^ Bit[923] ^ Bit[966] ^ Bit[1018] ^ Bit[1067] ^ Bit[1115] ^ Bit[1191] ^ Bit[1192];
				Check_42 <= Bit[35] ^ Bit[59] ^ Bit[99] ^ Bit[167] ^ Bit[201] ^ Bit[280] ^ Bit[333] ^ Bit[437] ^ Bit[534] ^ Bit[615] ^ Bit[771] ^ Bit[847] ^ Bit[880] ^ Bit[942] ^ Bit[977] ^ Bit[1044] ^ Bit[1060] ^ Bit[1110] ^ Bit[1192] ^ Bit[1193];
				Check_43 <= Bit[11] ^ Bit[95] ^ Bit[115] ^ Bit[176] ^ Bit[238] ^ Bit[281] ^ Bit[381] ^ Bit[387] ^ Bit[484] ^ Bit[720] ^ Bit[768] ^ Bit[816] ^ Bit[905] ^ Bit[946] ^ Bit[980] ^ Bit[1019] ^ Bit[1093] ^ Bit[1104] ^ Bit[1193] ^ Bit[1194];
				Check_44 <= Bit[20] ^ Bit[69] ^ Bit[125] ^ Bit[173] ^ Bit[202] ^ Bit[271] ^ Bit[322] ^ Bit[429] ^ Bit[518] ^ Bit[630] ^ Bit[691] ^ Bit[859] ^ Bit[901] ^ Bit[916] ^ Bit[995] ^ Bit[1027] ^ Bit[1094] ^ Bit[1125] ^ Bit[1194] ^ Bit[1195];
				Check_45 <= Bit[15] ^ Bit[90] ^ Bit[107] ^ Bit[189] ^ Bit[207] ^ Bit[274] ^ Bit[371] ^ Bit[426] ^ Bit[537] ^ Bit[594] ^ Bit[670] ^ Bit[726] ^ Bit[905] ^ Bit[949] ^ Bit[974] ^ Bit[1034] ^ Bit[1064] ^ Bit[1109] ^ Bit[1195] ^ Bit[1196];
				Check_46 <= Bit[34] ^ Bit[93] ^ Bit[132] ^ Bit[188] ^ Bit[205] ^ Bit[259] ^ Bit[435] ^ Bit[523] ^ Bit[559] ^ Bit[621] ^ Bit[646] ^ Bit[692] ^ Bit[909] ^ Bit[933] ^ Bit[969] ^ Bit[1047] ^ Bit[1074] ^ Bit[1138] ^ Bit[1196] ^ Bit[1197];
				Check_47 <= Bit[5] ^ Bit[63] ^ Bit[98] ^ Bit[169] ^ Bit[233] ^ Bit[251] ^ Bit[300] ^ Bit[367] ^ Bit[446] ^ Bit[680] ^ Bit[744] ^ Bit[798] ^ Bit[876] ^ Bit[924] ^ Bit[967] ^ Bit[1019] ^ Bit[1068] ^ Bit[1116] ^ Bit[1197] ^ Bit[1198];
				Check_48 <= Bit[36] ^ Bit[60] ^ Bit[100] ^ Bit[168] ^ Bit[202] ^ Bit[281] ^ Bit[334] ^ Bit[438] ^ Bit[535] ^ Bit[616] ^ Bit[772] ^ Bit[848] ^ Bit[881] ^ Bit[943] ^ Bit[978] ^ Bit[1045] ^ Bit[1061] ^ Bit[1111] ^ Bit[1198] ^ Bit[1199];
				Check_49 <= Bit[12] ^ Bit[48] ^ Bit[116] ^ Bit[177] ^ Bit[239] ^ Bit[282] ^ Bit[382] ^ Bit[388] ^ Bit[485] ^ Bit[721] ^ Bit[769] ^ Bit[817] ^ Bit[906] ^ Bit[947] ^ Bit[981] ^ Bit[1020] ^ Bit[1094] ^ Bit[1105] ^ Bit[1199] ^ Bit[1200];
				Check_50 <= Bit[21] ^ Bit[70] ^ Bit[126] ^ Bit[174] ^ Bit[203] ^ Bit[272] ^ Bit[323] ^ Bit[430] ^ Bit[519] ^ Bit[631] ^ Bit[692] ^ Bit[860] ^ Bit[902] ^ Bit[917] ^ Bit[996] ^ Bit[1028] ^ Bit[1095] ^ Bit[1126] ^ Bit[1200] ^ Bit[1201];
				Check_51 <= Bit[16] ^ Bit[91] ^ Bit[108] ^ Bit[190] ^ Bit[208] ^ Bit[275] ^ Bit[372] ^ Bit[427] ^ Bit[538] ^ Bit[595] ^ Bit[671] ^ Bit[727] ^ Bit[906] ^ Bit[950] ^ Bit[975] ^ Bit[1035] ^ Bit[1065] ^ Bit[1110] ^ Bit[1201] ^ Bit[1202];
				Check_52 <= Bit[35] ^ Bit[94] ^ Bit[133] ^ Bit[189] ^ Bit[206] ^ Bit[260] ^ Bit[436] ^ Bit[524] ^ Bit[560] ^ Bit[622] ^ Bit[647] ^ Bit[693] ^ Bit[910] ^ Bit[934] ^ Bit[970] ^ Bit[1048] ^ Bit[1075] ^ Bit[1139] ^ Bit[1202] ^ Bit[1203];
				Check_53 <= Bit[6] ^ Bit[64] ^ Bit[99] ^ Bit[170] ^ Bit[234] ^ Bit[252] ^ Bit[301] ^ Bit[368] ^ Bit[447] ^ Bit[681] ^ Bit[745] ^ Bit[799] ^ Bit[877] ^ Bit[925] ^ Bit[968] ^ Bit[1020] ^ Bit[1069] ^ Bit[1117] ^ Bit[1203] ^ Bit[1204];
				Check_54 <= Bit[37] ^ Bit[61] ^ Bit[101] ^ Bit[169] ^ Bit[203] ^ Bit[282] ^ Bit[335] ^ Bit[439] ^ Bit[536] ^ Bit[617] ^ Bit[773] ^ Bit[849] ^ Bit[882] ^ Bit[944] ^ Bit[979] ^ Bit[1046] ^ Bit[1062] ^ Bit[1112] ^ Bit[1204] ^ Bit[1205];
				Check_55 <= Bit[13] ^ Bit[49] ^ Bit[117] ^ Bit[178] ^ Bit[192] ^ Bit[283] ^ Bit[383] ^ Bit[389] ^ Bit[486] ^ Bit[722] ^ Bit[770] ^ Bit[818] ^ Bit[907] ^ Bit[948] ^ Bit[982] ^ Bit[1021] ^ Bit[1095] ^ Bit[1106] ^ Bit[1205] ^ Bit[1206];
				Check_56 <= Bit[22] ^ Bit[71] ^ Bit[127] ^ Bit[175] ^ Bit[204] ^ Bit[273] ^ Bit[324] ^ Bit[431] ^ Bit[520] ^ Bit[632] ^ Bit[693] ^ Bit[861] ^ Bit[903] ^ Bit[918] ^ Bit[997] ^ Bit[1029] ^ Bit[1096] ^ Bit[1127] ^ Bit[1206] ^ Bit[1207];
				Check_57 <= Bit[17] ^ Bit[92] ^ Bit[109] ^ Bit[191] ^ Bit[209] ^ Bit[276] ^ Bit[373] ^ Bit[428] ^ Bit[539] ^ Bit[596] ^ Bit[624] ^ Bit[728] ^ Bit[907] ^ Bit[951] ^ Bit[976] ^ Bit[1036] ^ Bit[1066] ^ Bit[1111] ^ Bit[1207] ^ Bit[1208];
				Check_58 <= Bit[36] ^ Bit[95] ^ Bit[134] ^ Bit[190] ^ Bit[207] ^ Bit[261] ^ Bit[437] ^ Bit[525] ^ Bit[561] ^ Bit[623] ^ Bit[648] ^ Bit[694] ^ Bit[911] ^ Bit[935] ^ Bit[971] ^ Bit[1049] ^ Bit[1076] ^ Bit[1140] ^ Bit[1208] ^ Bit[1209];
				Check_59 <= Bit[7] ^ Bit[65] ^ Bit[100] ^ Bit[171] ^ Bit[235] ^ Bit[253] ^ Bit[302] ^ Bit[369] ^ Bit[448] ^ Bit[682] ^ Bit[746] ^ Bit[800] ^ Bit[878] ^ Bit[926] ^ Bit[969] ^ Bit[1021] ^ Bit[1070] ^ Bit[1118] ^ Bit[1209] ^ Bit[1210];
				Check_60 <= Bit[38] ^ Bit[62] ^ Bit[102] ^ Bit[170] ^ Bit[204] ^ Bit[283] ^ Bit[288] ^ Bit[440] ^ Bit[537] ^ Bit[618] ^ Bit[774] ^ Bit[850] ^ Bit[883] ^ Bit[945] ^ Bit[980] ^ Bit[1047] ^ Bit[1063] ^ Bit[1113] ^ Bit[1210] ^ Bit[1211];
				Check_61 <= Bit[14] ^ Bit[50] ^ Bit[118] ^ Bit[179] ^ Bit[193] ^ Bit[284] ^ Bit[336] ^ Bit[390] ^ Bit[487] ^ Bit[723] ^ Bit[771] ^ Bit[819] ^ Bit[908] ^ Bit[949] ^ Bit[983] ^ Bit[1022] ^ Bit[1096] ^ Bit[1107] ^ Bit[1211] ^ Bit[1212];
				Check_62 <= Bit[23] ^ Bit[72] ^ Bit[128] ^ Bit[176] ^ Bit[205] ^ Bit[274] ^ Bit[325] ^ Bit[384] ^ Bit[521] ^ Bit[633] ^ Bit[694] ^ Bit[862] ^ Bit[904] ^ Bit[919] ^ Bit[998] ^ Bit[1030] ^ Bit[1097] ^ Bit[1128] ^ Bit[1212] ^ Bit[1213];
				Check_63 <= Bit[18] ^ Bit[93] ^ Bit[110] ^ Bit[144] ^ Bit[210] ^ Bit[277] ^ Bit[374] ^ Bit[429] ^ Bit[540] ^ Bit[597] ^ Bit[625] ^ Bit[729] ^ Bit[908] ^ Bit[952] ^ Bit[977] ^ Bit[1037] ^ Bit[1067] ^ Bit[1112] ^ Bit[1213] ^ Bit[1214];
				Check_64 <= Bit[37] ^ Bit[48] ^ Bit[135] ^ Bit[191] ^ Bit[208] ^ Bit[262] ^ Bit[438] ^ Bit[526] ^ Bit[562] ^ Bit[576] ^ Bit[649] ^ Bit[695] ^ Bit[864] ^ Bit[936] ^ Bit[972] ^ Bit[1050] ^ Bit[1077] ^ Bit[1141] ^ Bit[1214] ^ Bit[1215];
				Check_65 <= Bit[8] ^ Bit[66] ^ Bit[101] ^ Bit[172] ^ Bit[236] ^ Bit[254] ^ Bit[303] ^ Bit[370] ^ Bit[449] ^ Bit[683] ^ Bit[747] ^ Bit[801] ^ Bit[879] ^ Bit[927] ^ Bit[970] ^ Bit[1022] ^ Bit[1071] ^ Bit[1119] ^ Bit[1215] ^ Bit[1216];
				Check_66 <= Bit[39] ^ Bit[63] ^ Bit[103] ^ Bit[171] ^ Bit[205] ^ Bit[284] ^ Bit[289] ^ Bit[441] ^ Bit[538] ^ Bit[619] ^ Bit[775] ^ Bit[851] ^ Bit[884] ^ Bit[946] ^ Bit[981] ^ Bit[1048] ^ Bit[1064] ^ Bit[1114] ^ Bit[1216] ^ Bit[1217];
				Check_67 <= Bit[15] ^ Bit[51] ^ Bit[119] ^ Bit[180] ^ Bit[194] ^ Bit[285] ^ Bit[337] ^ Bit[391] ^ Bit[488] ^ Bit[724] ^ Bit[772] ^ Bit[820] ^ Bit[909] ^ Bit[950] ^ Bit[984] ^ Bit[1023] ^ Bit[1097] ^ Bit[1108] ^ Bit[1217] ^ Bit[1218];
				Check_68 <= Bit[24] ^ Bit[73] ^ Bit[129] ^ Bit[177] ^ Bit[206] ^ Bit[275] ^ Bit[326] ^ Bit[385] ^ Bit[522] ^ Bit[634] ^ Bit[695] ^ Bit[863] ^ Bit[905] ^ Bit[920] ^ Bit[999] ^ Bit[1031] ^ Bit[1098] ^ Bit[1129] ^ Bit[1218] ^ Bit[1219];
				Check_69 <= Bit[19] ^ Bit[94] ^ Bit[111] ^ Bit[145] ^ Bit[211] ^ Bit[278] ^ Bit[375] ^ Bit[430] ^ Bit[541] ^ Bit[598] ^ Bit[626] ^ Bit[730] ^ Bit[909] ^ Bit[953] ^ Bit[978] ^ Bit[1038] ^ Bit[1068] ^ Bit[1113] ^ Bit[1219] ^ Bit[1220];
				Check_70 <= Bit[38] ^ Bit[49] ^ Bit[136] ^ Bit[144] ^ Bit[209] ^ Bit[263] ^ Bit[439] ^ Bit[527] ^ Bit[563] ^ Bit[577] ^ Bit[650] ^ Bit[696] ^ Bit[865] ^ Bit[937] ^ Bit[973] ^ Bit[1051] ^ Bit[1078] ^ Bit[1142] ^ Bit[1220] ^ Bit[1221];
				Check_71 <= Bit[9] ^ Bit[67] ^ Bit[102] ^ Bit[173] ^ Bit[237] ^ Bit[255] ^ Bit[304] ^ Bit[371] ^ Bit[450] ^ Bit[684] ^ Bit[748] ^ Bit[802] ^ Bit[880] ^ Bit[928] ^ Bit[971] ^ Bit[1023] ^ Bit[1072] ^ Bit[1120] ^ Bit[1221] ^ Bit[1222];
				Check_72 <= Bit[40] ^ Bit[64] ^ Bit[104] ^ Bit[172] ^ Bit[206] ^ Bit[285] ^ Bit[290] ^ Bit[442] ^ Bit[539] ^ Bit[620] ^ Bit[776] ^ Bit[852] ^ Bit[885] ^ Bit[947] ^ Bit[982] ^ Bit[1049] ^ Bit[1065] ^ Bit[1115] ^ Bit[1222] ^ Bit[1223];
				Check_73 <= Bit[16] ^ Bit[52] ^ Bit[120] ^ Bit[181] ^ Bit[195] ^ Bit[286] ^ Bit[338] ^ Bit[392] ^ Bit[489] ^ Bit[725] ^ Bit[773] ^ Bit[821] ^ Bit[910] ^ Bit[951] ^ Bit[985] ^ Bit[1024] ^ Bit[1098] ^ Bit[1109] ^ Bit[1223] ^ Bit[1224];
				Check_74 <= Bit[25] ^ Bit[74] ^ Bit[130] ^ Bit[178] ^ Bit[207] ^ Bit[276] ^ Bit[327] ^ Bit[386] ^ Bit[523] ^ Bit[635] ^ Bit[696] ^ Bit[816] ^ Bit[906] ^ Bit[921] ^ Bit[1000] ^ Bit[1032] ^ Bit[1099] ^ Bit[1130] ^ Bit[1224] ^ Bit[1225];
				Check_75 <= Bit[20] ^ Bit[95] ^ Bit[112] ^ Bit[146] ^ Bit[212] ^ Bit[279] ^ Bit[376] ^ Bit[431] ^ Bit[542] ^ Bit[599] ^ Bit[627] ^ Bit[731] ^ Bit[910] ^ Bit[954] ^ Bit[979] ^ Bit[1039] ^ Bit[1069] ^ Bit[1114] ^ Bit[1225] ^ Bit[1226];
				Check_76 <= Bit[39] ^ Bit[50] ^ Bit[137] ^ Bit[145] ^ Bit[210] ^ Bit[264] ^ Bit[440] ^ Bit[480] ^ Bit[564] ^ Bit[578] ^ Bit[651] ^ Bit[697] ^ Bit[866] ^ Bit[938] ^ Bit[974] ^ Bit[1052] ^ Bit[1079] ^ Bit[1143] ^ Bit[1226] ^ Bit[1227];
				Check_77 <= Bit[10] ^ Bit[68] ^ Bit[103] ^ Bit[174] ^ Bit[238] ^ Bit[256] ^ Bit[305] ^ Bit[372] ^ Bit[451] ^ Bit[685] ^ Bit[749] ^ Bit[803] ^ Bit[881] ^ Bit[929] ^ Bit[972] ^ Bit[1024] ^ Bit[1073] ^ Bit[1121] ^ Bit[1227] ^ Bit[1228];
				Check_78 <= Bit[41] ^ Bit[65] ^ Bit[105] ^ Bit[173] ^ Bit[207] ^ Bit[286] ^ Bit[291] ^ Bit[443] ^ Bit[540] ^ Bit[621] ^ Bit[777] ^ Bit[853] ^ Bit[886] ^ Bit[948] ^ Bit[983] ^ Bit[1050] ^ Bit[1066] ^ Bit[1116] ^ Bit[1228] ^ Bit[1229];
				Check_79 <= Bit[17] ^ Bit[53] ^ Bit[121] ^ Bit[182] ^ Bit[196] ^ Bit[287] ^ Bit[339] ^ Bit[393] ^ Bit[490] ^ Bit[726] ^ Bit[774] ^ Bit[822] ^ Bit[911] ^ Bit[952] ^ Bit[986] ^ Bit[1025] ^ Bit[1099] ^ Bit[1110] ^ Bit[1229] ^ Bit[1230];
				Check_80 <= Bit[26] ^ Bit[75] ^ Bit[131] ^ Bit[179] ^ Bit[208] ^ Bit[277] ^ Bit[328] ^ Bit[387] ^ Bit[524] ^ Bit[636] ^ Bit[697] ^ Bit[817] ^ Bit[907] ^ Bit[922] ^ Bit[1001] ^ Bit[1033] ^ Bit[1100] ^ Bit[1131] ^ Bit[1230] ^ Bit[1231];
				Check_81 <= Bit[21] ^ Bit[48] ^ Bit[113] ^ Bit[147] ^ Bit[213] ^ Bit[280] ^ Bit[377] ^ Bit[384] ^ Bit[543] ^ Bit[600] ^ Bit[628] ^ Bit[732] ^ Bit[911] ^ Bit[955] ^ Bit[980] ^ Bit[1040] ^ Bit[1070] ^ Bit[1115] ^ Bit[1231] ^ Bit[1232];
				Check_82 <= Bit[40] ^ Bit[51] ^ Bit[138] ^ Bit[146] ^ Bit[211] ^ Bit[265] ^ Bit[441] ^ Bit[481] ^ Bit[565] ^ Bit[579] ^ Bit[652] ^ Bit[698] ^ Bit[867] ^ Bit[939] ^ Bit[975] ^ Bit[1053] ^ Bit[1080] ^ Bit[1144] ^ Bit[1232] ^ Bit[1233];
				Check_83 <= Bit[11] ^ Bit[69] ^ Bit[104] ^ Bit[175] ^ Bit[239] ^ Bit[257] ^ Bit[306] ^ Bit[373] ^ Bit[452] ^ Bit[686] ^ Bit[750] ^ Bit[804] ^ Bit[882] ^ Bit[930] ^ Bit[973] ^ Bit[1025] ^ Bit[1074] ^ Bit[1122] ^ Bit[1233] ^ Bit[1234];
				Check_84 <= Bit[42] ^ Bit[66] ^ Bit[106] ^ Bit[174] ^ Bit[208] ^ Bit[287] ^ Bit[292] ^ Bit[444] ^ Bit[541] ^ Bit[622] ^ Bit[778] ^ Bit[854] ^ Bit[887] ^ Bit[949] ^ Bit[984] ^ Bit[1051] ^ Bit[1067] ^ Bit[1117] ^ Bit[1234] ^ Bit[1235];
				Check_85 <= Bit[18] ^ Bit[54] ^ Bit[122] ^ Bit[183] ^ Bit[197] ^ Bit[240] ^ Bit[340] ^ Bit[394] ^ Bit[491] ^ Bit[727] ^ Bit[775] ^ Bit[823] ^ Bit[864] ^ Bit[953] ^ Bit[987] ^ Bit[1026] ^ Bit[1100] ^ Bit[1111] ^ Bit[1235] ^ Bit[1236];
				Check_86 <= Bit[27] ^ Bit[76] ^ Bit[132] ^ Bit[180] ^ Bit[209] ^ Bit[278] ^ Bit[329] ^ Bit[388] ^ Bit[525] ^ Bit[637] ^ Bit[698] ^ Bit[818] ^ Bit[908] ^ Bit[923] ^ Bit[1002] ^ Bit[1034] ^ Bit[1101] ^ Bit[1132] ^ Bit[1236] ^ Bit[1237];
				Check_87 <= Bit[22] ^ Bit[49] ^ Bit[114] ^ Bit[148] ^ Bit[214] ^ Bit[281] ^ Bit[378] ^ Bit[385] ^ Bit[544] ^ Bit[601] ^ Bit[629] ^ Bit[733] ^ Bit[864] ^ Bit[956] ^ Bit[981] ^ Bit[1041] ^ Bit[1071] ^ Bit[1116] ^ Bit[1237] ^ Bit[1238];
				Check_88 <= Bit[41] ^ Bit[52] ^ Bit[139] ^ Bit[147] ^ Bit[212] ^ Bit[266] ^ Bit[442] ^ Bit[482] ^ Bit[566] ^ Bit[580] ^ Bit[653] ^ Bit[699] ^ Bit[868] ^ Bit[940] ^ Bit[976] ^ Bit[1054] ^ Bit[1081] ^ Bit[1145] ^ Bit[1238] ^ Bit[1239];
				Check_89 <= Bit[12] ^ Bit[70] ^ Bit[105] ^ Bit[176] ^ Bit[192] ^ Bit[258] ^ Bit[307] ^ Bit[374] ^ Bit[453] ^ Bit[687] ^ Bit[751] ^ Bit[805] ^ Bit[883] ^ Bit[931] ^ Bit[974] ^ Bit[1026] ^ Bit[1075] ^ Bit[1123] ^ Bit[1239] ^ Bit[1240];
				Check_90 <= Bit[43] ^ Bit[67] ^ Bit[107] ^ Bit[175] ^ Bit[209] ^ Bit[240] ^ Bit[293] ^ Bit[445] ^ Bit[542] ^ Bit[623] ^ Bit[779] ^ Bit[855] ^ Bit[888] ^ Bit[950] ^ Bit[985] ^ Bit[1052] ^ Bit[1068] ^ Bit[1118] ^ Bit[1240] ^ Bit[1241];
				Check_91 <= Bit[19] ^ Bit[55] ^ Bit[123] ^ Bit[184] ^ Bit[198] ^ Bit[241] ^ Bit[341] ^ Bit[395] ^ Bit[492] ^ Bit[728] ^ Bit[776] ^ Bit[824] ^ Bit[865] ^ Bit[954] ^ Bit[988] ^ Bit[1027] ^ Bit[1101] ^ Bit[1112] ^ Bit[1241] ^ Bit[1242];
				Check_92 <= Bit[28] ^ Bit[77] ^ Bit[133] ^ Bit[181] ^ Bit[210] ^ Bit[279] ^ Bit[330] ^ Bit[389] ^ Bit[526] ^ Bit[638] ^ Bit[699] ^ Bit[819] ^ Bit[909] ^ Bit[924] ^ Bit[1003] ^ Bit[1035] ^ Bit[1102] ^ Bit[1133] ^ Bit[1242] ^ Bit[1243];
				Check_93 <= Bit[23] ^ Bit[50] ^ Bit[115] ^ Bit[149] ^ Bit[215] ^ Bit[282] ^ Bit[379] ^ Bit[386] ^ Bit[545] ^ Bit[602] ^ Bit[630] ^ Bit[734] ^ Bit[865] ^ Bit[957] ^ Bit[982] ^ Bit[1042] ^ Bit[1072] ^ Bit[1117] ^ Bit[1243] ^ Bit[1244];
				Check_94 <= Bit[42] ^ Bit[53] ^ Bit[140] ^ Bit[148] ^ Bit[213] ^ Bit[267] ^ Bit[443] ^ Bit[483] ^ Bit[567] ^ Bit[581] ^ Bit[654] ^ Bit[700] ^ Bit[869] ^ Bit[941] ^ Bit[977] ^ Bit[1055] ^ Bit[1082] ^ Bit[1146] ^ Bit[1244] ^ Bit[1245];
				Check_95 <= Bit[13] ^ Bit[71] ^ Bit[106] ^ Bit[177] ^ Bit[193] ^ Bit[259] ^ Bit[308] ^ Bit[375] ^ Bit[454] ^ Bit[688] ^ Bit[752] ^ Bit[806] ^ Bit[884] ^ Bit[932] ^ Bit[975] ^ Bit[1027] ^ Bit[1076] ^ Bit[1124] ^ Bit[1245] ^ Bit[1246];
				Check_96 <= Bit[44] ^ Bit[68] ^ Bit[108] ^ Bit[176] ^ Bit[210] ^ Bit[241] ^ Bit[294] ^ Bit[446] ^ Bit[543] ^ Bit[576] ^ Bit[780] ^ Bit[856] ^ Bit[889] ^ Bit[951] ^ Bit[986] ^ Bit[1053] ^ Bit[1069] ^ Bit[1119] ^ Bit[1246] ^ Bit[1247];
				Check_97 <= Bit[20] ^ Bit[56] ^ Bit[124] ^ Bit[185] ^ Bit[199] ^ Bit[242] ^ Bit[342] ^ Bit[396] ^ Bit[493] ^ Bit[729] ^ Bit[777] ^ Bit[825] ^ Bit[866] ^ Bit[955] ^ Bit[989] ^ Bit[1028] ^ Bit[1102] ^ Bit[1113] ^ Bit[1247] ^ Bit[1248];
				Check_98 <= Bit[29] ^ Bit[78] ^ Bit[134] ^ Bit[182] ^ Bit[211] ^ Bit[280] ^ Bit[331] ^ Bit[390] ^ Bit[527] ^ Bit[639] ^ Bit[700] ^ Bit[820] ^ Bit[910] ^ Bit[925] ^ Bit[1004] ^ Bit[1036] ^ Bit[1103] ^ Bit[1134] ^ Bit[1248] ^ Bit[1249];
				Check_99 <= Bit[24] ^ Bit[51] ^ Bit[116] ^ Bit[150] ^ Bit[216] ^ Bit[283] ^ Bit[380] ^ Bit[387] ^ Bit[546] ^ Bit[603] ^ Bit[631] ^ Bit[735] ^ Bit[866] ^ Bit[958] ^ Bit[983] ^ Bit[1043] ^ Bit[1073] ^ Bit[1118] ^ Bit[1249] ^ Bit[1250];
				Check_100 <= Bit[43] ^ Bit[54] ^ Bit[141] ^ Bit[149] ^ Bit[214] ^ Bit[268] ^ Bit[444] ^ Bit[484] ^ Bit[568] ^ Bit[582] ^ Bit[655] ^ Bit[701] ^ Bit[870] ^ Bit[942] ^ Bit[978] ^ Bit[1008] ^ Bit[1083] ^ Bit[1147] ^ Bit[1250] ^ Bit[1251];
				Check_101 <= Bit[14] ^ Bit[72] ^ Bit[107] ^ Bit[178] ^ Bit[194] ^ Bit[260] ^ Bit[309] ^ Bit[376] ^ Bit[455] ^ Bit[689] ^ Bit[753] ^ Bit[807] ^ Bit[885] ^ Bit[933] ^ Bit[976] ^ Bit[1028] ^ Bit[1077] ^ Bit[1125] ^ Bit[1251] ^ Bit[1252];
				Check_102 <= Bit[45] ^ Bit[69] ^ Bit[109] ^ Bit[177] ^ Bit[211] ^ Bit[242] ^ Bit[295] ^ Bit[447] ^ Bit[544] ^ Bit[577] ^ Bit[781] ^ Bit[857] ^ Bit[890] ^ Bit[952] ^ Bit[987] ^ Bit[1054] ^ Bit[1070] ^ Bit[1120] ^ Bit[1252] ^ Bit[1253];
				Check_103 <= Bit[21] ^ Bit[57] ^ Bit[125] ^ Bit[186] ^ Bit[200] ^ Bit[243] ^ Bit[343] ^ Bit[397] ^ Bit[494] ^ Bit[730] ^ Bit[778] ^ Bit[826] ^ Bit[867] ^ Bit[956] ^ Bit[990] ^ Bit[1029] ^ Bit[1103] ^ Bit[1114] ^ Bit[1253] ^ Bit[1254];
				Check_104 <= Bit[30] ^ Bit[79] ^ Bit[135] ^ Bit[183] ^ Bit[212] ^ Bit[281] ^ Bit[332] ^ Bit[391] ^ Bit[480] ^ Bit[640] ^ Bit[701] ^ Bit[821] ^ Bit[911] ^ Bit[926] ^ Bit[1005] ^ Bit[1037] ^ Bit[1056] ^ Bit[1135] ^ Bit[1254] ^ Bit[1255];
				Check_105 <= Bit[25] ^ Bit[52] ^ Bit[117] ^ Bit[151] ^ Bit[217] ^ Bit[284] ^ Bit[381] ^ Bit[388] ^ Bit[547] ^ Bit[604] ^ Bit[632] ^ Bit[736] ^ Bit[867] ^ Bit[959] ^ Bit[984] ^ Bit[1044] ^ Bit[1074] ^ Bit[1119] ^ Bit[1255] ^ Bit[1256];
				Check_106 <= Bit[44] ^ Bit[55] ^ Bit[142] ^ Bit[150] ^ Bit[215] ^ Bit[269] ^ Bit[445] ^ Bit[485] ^ Bit[569] ^ Bit[583] ^ Bit[656] ^ Bit[702] ^ Bit[871] ^ Bit[943] ^ Bit[979] ^ Bit[1009] ^ Bit[1084] ^ Bit[1148] ^ Bit[1256] ^ Bit[1257];
				Check_107 <= Bit[15] ^ Bit[73] ^ Bit[108] ^ Bit[179] ^ Bit[195] ^ Bit[261] ^ Bit[310] ^ Bit[377] ^ Bit[456] ^ Bit[690] ^ Bit[754] ^ Bit[808] ^ Bit[886] ^ Bit[934] ^ Bit[977] ^ Bit[1029] ^ Bit[1078] ^ Bit[1126] ^ Bit[1257] ^ Bit[1258];
				Check_108 <= Bit[46] ^ Bit[70] ^ Bit[110] ^ Bit[178] ^ Bit[212] ^ Bit[243] ^ Bit[296] ^ Bit[448] ^ Bit[545] ^ Bit[578] ^ Bit[782] ^ Bit[858] ^ Bit[891] ^ Bit[953] ^ Bit[988] ^ Bit[1055] ^ Bit[1071] ^ Bit[1121] ^ Bit[1258] ^ Bit[1259];
				Check_109 <= Bit[22] ^ Bit[58] ^ Bit[126] ^ Bit[187] ^ Bit[201] ^ Bit[244] ^ Bit[344] ^ Bit[398] ^ Bit[495] ^ Bit[731] ^ Bit[779] ^ Bit[827] ^ Bit[868] ^ Bit[957] ^ Bit[991] ^ Bit[1030] ^ Bit[1056] ^ Bit[1115] ^ Bit[1259] ^ Bit[1260];
				Check_110 <= Bit[31] ^ Bit[80] ^ Bit[136] ^ Bit[184] ^ Bit[213] ^ Bit[282] ^ Bit[333] ^ Bit[392] ^ Bit[481] ^ Bit[641] ^ Bit[702] ^ Bit[822] ^ Bit[864] ^ Bit[927] ^ Bit[1006] ^ Bit[1038] ^ Bit[1057] ^ Bit[1136] ^ Bit[1260] ^ Bit[1261];
				Check_111 <= Bit[26] ^ Bit[53] ^ Bit[118] ^ Bit[152] ^ Bit[218] ^ Bit[285] ^ Bit[382] ^ Bit[389] ^ Bit[548] ^ Bit[605] ^ Bit[633] ^ Bit[737] ^ Bit[868] ^ Bit[912] ^ Bit[985] ^ Bit[1045] ^ Bit[1075] ^ Bit[1120] ^ Bit[1261] ^ Bit[1262];
				Check_112 <= Bit[45] ^ Bit[56] ^ Bit[143] ^ Bit[151] ^ Bit[216] ^ Bit[270] ^ Bit[446] ^ Bit[486] ^ Bit[570] ^ Bit[584] ^ Bit[657] ^ Bit[703] ^ Bit[872] ^ Bit[944] ^ Bit[980] ^ Bit[1010] ^ Bit[1085] ^ Bit[1149] ^ Bit[1262] ^ Bit[1263];
				Check_113 <= Bit[16] ^ Bit[74] ^ Bit[109] ^ Bit[180] ^ Bit[196] ^ Bit[262] ^ Bit[311] ^ Bit[378] ^ Bit[457] ^ Bit[691] ^ Bit[755] ^ Bit[809] ^ Bit[887] ^ Bit[935] ^ Bit[978] ^ Bit[1030] ^ Bit[1079] ^ Bit[1127] ^ Bit[1263] ^ Bit[1264];
				Check_114 <= Bit[47] ^ Bit[71] ^ Bit[111] ^ Bit[179] ^ Bit[213] ^ Bit[244] ^ Bit[297] ^ Bit[449] ^ Bit[546] ^ Bit[579] ^ Bit[783] ^ Bit[859] ^ Bit[892] ^ Bit[954] ^ Bit[989] ^ Bit[1008] ^ Bit[1072] ^ Bit[1122] ^ Bit[1264] ^ Bit[1265];
				Check_115 <= Bit[23] ^ Bit[59] ^ Bit[127] ^ Bit[188] ^ Bit[202] ^ Bit[245] ^ Bit[345] ^ Bit[399] ^ Bit[496] ^ Bit[732] ^ Bit[780] ^ Bit[828] ^ Bit[869] ^ Bit[958] ^ Bit[992] ^ Bit[1031] ^ Bit[1057] ^ Bit[1116] ^ Bit[1265] ^ Bit[1266];
				Check_116 <= Bit[32] ^ Bit[81] ^ Bit[137] ^ Bit[185] ^ Bit[214] ^ Bit[283] ^ Bit[334] ^ Bit[393] ^ Bit[482] ^ Bit[642] ^ Bit[703] ^ Bit[823] ^ Bit[865] ^ Bit[928] ^ Bit[1007] ^ Bit[1039] ^ Bit[1058] ^ Bit[1137] ^ Bit[1266] ^ Bit[1267];
				Check_117 <= Bit[27] ^ Bit[54] ^ Bit[119] ^ Bit[153] ^ Bit[219] ^ Bit[286] ^ Bit[383] ^ Bit[390] ^ Bit[549] ^ Bit[606] ^ Bit[634] ^ Bit[738] ^ Bit[869] ^ Bit[913] ^ Bit[986] ^ Bit[1046] ^ Bit[1076] ^ Bit[1121] ^ Bit[1267] ^ Bit[1268];
				Check_118 <= Bit[46] ^ Bit[57] ^ Bit[96] ^ Bit[152] ^ Bit[217] ^ Bit[271] ^ Bit[447] ^ Bit[487] ^ Bit[571] ^ Bit[585] ^ Bit[658] ^ Bit[704] ^ Bit[873] ^ Bit[945] ^ Bit[981] ^ Bit[1011] ^ Bit[1086] ^ Bit[1150] ^ Bit[1268] ^ Bit[1269];
				Check_119 <= Bit[17] ^ Bit[75] ^ Bit[110] ^ Bit[181] ^ Bit[197] ^ Bit[263] ^ Bit[312] ^ Bit[379] ^ Bit[458] ^ Bit[692] ^ Bit[756] ^ Bit[810] ^ Bit[888] ^ Bit[936] ^ Bit[979] ^ Bit[1031] ^ Bit[1080] ^ Bit[1128] ^ Bit[1269] ^ Bit[1270];
				Check_120 <= Bit[0] ^ Bit[72] ^ Bit[112] ^ Bit[180] ^ Bit[214] ^ Bit[245] ^ Bit[298] ^ Bit[450] ^ Bit[547] ^ Bit[580] ^ Bit[784] ^ Bit[860] ^ Bit[893] ^ Bit[955] ^ Bit[990] ^ Bit[1009] ^ Bit[1073] ^ Bit[1123] ^ Bit[1270] ^ Bit[1271];
				Check_121 <= Bit[24] ^ Bit[60] ^ Bit[128] ^ Bit[189] ^ Bit[203] ^ Bit[246] ^ Bit[346] ^ Bit[400] ^ Bit[497] ^ Bit[733] ^ Bit[781] ^ Bit[829] ^ Bit[870] ^ Bit[959] ^ Bit[993] ^ Bit[1032] ^ Bit[1058] ^ Bit[1117] ^ Bit[1271] ^ Bit[1272];
				Check_122 <= Bit[33] ^ Bit[82] ^ Bit[138] ^ Bit[186] ^ Bit[215] ^ Bit[284] ^ Bit[335] ^ Bit[394] ^ Bit[483] ^ Bit[643] ^ Bit[704] ^ Bit[824] ^ Bit[866] ^ Bit[929] ^ Bit[960] ^ Bit[1040] ^ Bit[1059] ^ Bit[1138] ^ Bit[1272] ^ Bit[1273];
				Check_123 <= Bit[28] ^ Bit[55] ^ Bit[120] ^ Bit[154] ^ Bit[220] ^ Bit[287] ^ Bit[336] ^ Bit[391] ^ Bit[550] ^ Bit[607] ^ Bit[635] ^ Bit[739] ^ Bit[870] ^ Bit[914] ^ Bit[987] ^ Bit[1047] ^ Bit[1077] ^ Bit[1122] ^ Bit[1273] ^ Bit[1274];
				Check_124 <= Bit[47] ^ Bit[58] ^ Bit[97] ^ Bit[153] ^ Bit[218] ^ Bit[272] ^ Bit[448] ^ Bit[488] ^ Bit[572] ^ Bit[586] ^ Bit[659] ^ Bit[705] ^ Bit[874] ^ Bit[946] ^ Bit[982] ^ Bit[1012] ^ Bit[1087] ^ Bit[1151] ^ Bit[1274] ^ Bit[1275];
				Check_125 <= Bit[18] ^ Bit[76] ^ Bit[111] ^ Bit[182] ^ Bit[198] ^ Bit[264] ^ Bit[313] ^ Bit[380] ^ Bit[459] ^ Bit[693] ^ Bit[757] ^ Bit[811] ^ Bit[889] ^ Bit[937] ^ Bit[980] ^ Bit[1032] ^ Bit[1081] ^ Bit[1129] ^ Bit[1275] ^ Bit[1276];
				Check_126 <= Bit[1] ^ Bit[73] ^ Bit[113] ^ Bit[181] ^ Bit[215] ^ Bit[246] ^ Bit[299] ^ Bit[451] ^ Bit[548] ^ Bit[581] ^ Bit[785] ^ Bit[861] ^ Bit[894] ^ Bit[956] ^ Bit[991] ^ Bit[1010] ^ Bit[1074] ^ Bit[1124] ^ Bit[1276] ^ Bit[1277];
				Check_127 <= Bit[25] ^ Bit[61] ^ Bit[129] ^ Bit[190] ^ Bit[204] ^ Bit[247] ^ Bit[347] ^ Bit[401] ^ Bit[498] ^ Bit[734] ^ Bit[782] ^ Bit[830] ^ Bit[871] ^ Bit[912] ^ Bit[994] ^ Bit[1033] ^ Bit[1059] ^ Bit[1118] ^ Bit[1277] ^ Bit[1278];
				Check_128 <= Bit[34] ^ Bit[83] ^ Bit[139] ^ Bit[187] ^ Bit[216] ^ Bit[285] ^ Bit[288] ^ Bit[395] ^ Bit[484] ^ Bit[644] ^ Bit[705] ^ Bit[825] ^ Bit[867] ^ Bit[930] ^ Bit[961] ^ Bit[1041] ^ Bit[1060] ^ Bit[1139] ^ Bit[1278] ^ Bit[1279];
				Check_129 <= Bit[29] ^ Bit[56] ^ Bit[121] ^ Bit[155] ^ Bit[221] ^ Bit[240] ^ Bit[337] ^ Bit[392] ^ Bit[551] ^ Bit[608] ^ Bit[636] ^ Bit[740] ^ Bit[871] ^ Bit[915] ^ Bit[988] ^ Bit[1048] ^ Bit[1078] ^ Bit[1123] ^ Bit[1279] ^ Bit[1280];
				Check_130 <= Bit[0] ^ Bit[59] ^ Bit[98] ^ Bit[154] ^ Bit[219] ^ Bit[273] ^ Bit[449] ^ Bit[489] ^ Bit[573] ^ Bit[587] ^ Bit[660] ^ Bit[706] ^ Bit[875] ^ Bit[947] ^ Bit[983] ^ Bit[1013] ^ Bit[1088] ^ Bit[1104] ^ Bit[1280] ^ Bit[1281];
				Check_131 <= Bit[19] ^ Bit[77] ^ Bit[112] ^ Bit[183] ^ Bit[199] ^ Bit[265] ^ Bit[314] ^ Bit[381] ^ Bit[460] ^ Bit[694] ^ Bit[758] ^ Bit[812] ^ Bit[890] ^ Bit[938] ^ Bit[981] ^ Bit[1033] ^ Bit[1082] ^ Bit[1130] ^ Bit[1281] ^ Bit[1282];
				Check_132 <= Bit[2] ^ Bit[74] ^ Bit[114] ^ Bit[182] ^ Bit[216] ^ Bit[247] ^ Bit[300] ^ Bit[452] ^ Bit[549] ^ Bit[582] ^ Bit[786] ^ Bit[862] ^ Bit[895] ^ Bit[957] ^ Bit[992] ^ Bit[1011] ^ Bit[1075] ^ Bit[1125] ^ Bit[1282] ^ Bit[1283];
				Check_133 <= Bit[26] ^ Bit[62] ^ Bit[130] ^ Bit[191] ^ Bit[205] ^ Bit[248] ^ Bit[348] ^ Bit[402] ^ Bit[499] ^ Bit[735] ^ Bit[783] ^ Bit[831] ^ Bit[872] ^ Bit[913] ^ Bit[995] ^ Bit[1034] ^ Bit[1060] ^ Bit[1119] ^ Bit[1283] ^ Bit[1284];
				Check_134 <= Bit[35] ^ Bit[84] ^ Bit[140] ^ Bit[188] ^ Bit[217] ^ Bit[286] ^ Bit[289] ^ Bit[396] ^ Bit[485] ^ Bit[645] ^ Bit[706] ^ Bit[826] ^ Bit[868] ^ Bit[931] ^ Bit[962] ^ Bit[1042] ^ Bit[1061] ^ Bit[1140] ^ Bit[1284] ^ Bit[1285];
				Check_135 <= Bit[30] ^ Bit[57] ^ Bit[122] ^ Bit[156] ^ Bit[222] ^ Bit[241] ^ Bit[338] ^ Bit[393] ^ Bit[552] ^ Bit[609] ^ Bit[637] ^ Bit[741] ^ Bit[872] ^ Bit[916] ^ Bit[989] ^ Bit[1049] ^ Bit[1079] ^ Bit[1124] ^ Bit[1285] ^ Bit[1286];
				Check_136 <= Bit[1] ^ Bit[60] ^ Bit[99] ^ Bit[155] ^ Bit[220] ^ Bit[274] ^ Bit[450] ^ Bit[490] ^ Bit[574] ^ Bit[588] ^ Bit[661] ^ Bit[707] ^ Bit[876] ^ Bit[948] ^ Bit[984] ^ Bit[1014] ^ Bit[1089] ^ Bit[1105] ^ Bit[1286] ^ Bit[1287];
				Check_137 <= Bit[20] ^ Bit[78] ^ Bit[113] ^ Bit[184] ^ Bit[200] ^ Bit[266] ^ Bit[315] ^ Bit[382] ^ Bit[461] ^ Bit[695] ^ Bit[759] ^ Bit[813] ^ Bit[891] ^ Bit[939] ^ Bit[982] ^ Bit[1034] ^ Bit[1083] ^ Bit[1131] ^ Bit[1287] ^ Bit[1288];
				Check_138 <= Bit[3] ^ Bit[75] ^ Bit[115] ^ Bit[183] ^ Bit[217] ^ Bit[248] ^ Bit[301] ^ Bit[453] ^ Bit[550] ^ Bit[583] ^ Bit[787] ^ Bit[863] ^ Bit[896] ^ Bit[958] ^ Bit[993] ^ Bit[1012] ^ Bit[1076] ^ Bit[1126] ^ Bit[1288] ^ Bit[1289];
				Check_139 <= Bit[27] ^ Bit[63] ^ Bit[131] ^ Bit[144] ^ Bit[206] ^ Bit[249] ^ Bit[349] ^ Bit[403] ^ Bit[500] ^ Bit[736] ^ Bit[784] ^ Bit[832] ^ Bit[873] ^ Bit[914] ^ Bit[996] ^ Bit[1035] ^ Bit[1061] ^ Bit[1120] ^ Bit[1289] ^ Bit[1290];
				Check_140 <= Bit[36] ^ Bit[85] ^ Bit[141] ^ Bit[189] ^ Bit[218] ^ Bit[287] ^ Bit[290] ^ Bit[397] ^ Bit[486] ^ Bit[646] ^ Bit[707] ^ Bit[827] ^ Bit[869] ^ Bit[932] ^ Bit[963] ^ Bit[1043] ^ Bit[1062] ^ Bit[1141] ^ Bit[1290] ^ Bit[1291];
				Check_141 <= Bit[31] ^ Bit[58] ^ Bit[123] ^ Bit[157] ^ Bit[223] ^ Bit[242] ^ Bit[339] ^ Bit[394] ^ Bit[553] ^ Bit[610] ^ Bit[638] ^ Bit[742] ^ Bit[873] ^ Bit[917] ^ Bit[990] ^ Bit[1050] ^ Bit[1080] ^ Bit[1125] ^ Bit[1291] ^ Bit[1292];
				Check_142 <= Bit[2] ^ Bit[61] ^ Bit[100] ^ Bit[156] ^ Bit[221] ^ Bit[275] ^ Bit[451] ^ Bit[491] ^ Bit[575] ^ Bit[589] ^ Bit[662] ^ Bit[708] ^ Bit[877] ^ Bit[949] ^ Bit[985] ^ Bit[1015] ^ Bit[1090] ^ Bit[1106] ^ Bit[1292] ^ Bit[1293];
				Check_143 <= Bit[21] ^ Bit[79] ^ Bit[114] ^ Bit[185] ^ Bit[201] ^ Bit[267] ^ Bit[316] ^ Bit[383] ^ Bit[462] ^ Bit[696] ^ Bit[760] ^ Bit[814] ^ Bit[892] ^ Bit[940] ^ Bit[983] ^ Bit[1035] ^ Bit[1084] ^ Bit[1132] ^ Bit[1293] ^ Bit[1294];
				Check_144 <= Bit[4] ^ Bit[76] ^ Bit[116] ^ Bit[184] ^ Bit[218] ^ Bit[249] ^ Bit[302] ^ Bit[454] ^ Bit[551] ^ Bit[584] ^ Bit[788] ^ Bit[816] ^ Bit[897] ^ Bit[959] ^ Bit[994] ^ Bit[1013] ^ Bit[1077] ^ Bit[1127] ^ Bit[1294] ^ Bit[1295];
				Check_145 <= Bit[28] ^ Bit[64] ^ Bit[132] ^ Bit[145] ^ Bit[207] ^ Bit[250] ^ Bit[350] ^ Bit[404] ^ Bit[501] ^ Bit[737] ^ Bit[785] ^ Bit[833] ^ Bit[874] ^ Bit[915] ^ Bit[997] ^ Bit[1036] ^ Bit[1062] ^ Bit[1121] ^ Bit[1295] ^ Bit[1296];
				Check_146 <= Bit[37] ^ Bit[86] ^ Bit[142] ^ Bit[190] ^ Bit[219] ^ Bit[240] ^ Bit[291] ^ Bit[398] ^ Bit[487] ^ Bit[647] ^ Bit[708] ^ Bit[828] ^ Bit[870] ^ Bit[933] ^ Bit[964] ^ Bit[1044] ^ Bit[1063] ^ Bit[1142] ^ Bit[1296] ^ Bit[1297];
				Check_147 <= Bit[32] ^ Bit[59] ^ Bit[124] ^ Bit[158] ^ Bit[224] ^ Bit[243] ^ Bit[340] ^ Bit[395] ^ Bit[554] ^ Bit[611] ^ Bit[639] ^ Bit[743] ^ Bit[874] ^ Bit[918] ^ Bit[991] ^ Bit[1051] ^ Bit[1081] ^ Bit[1126] ^ Bit[1297] ^ Bit[1298];
				Check_148 <= Bit[3] ^ Bit[62] ^ Bit[101] ^ Bit[157] ^ Bit[222] ^ Bit[276] ^ Bit[452] ^ Bit[492] ^ Bit[528] ^ Bit[590] ^ Bit[663] ^ Bit[709] ^ Bit[878] ^ Bit[950] ^ Bit[986] ^ Bit[1016] ^ Bit[1091] ^ Bit[1107] ^ Bit[1298] ^ Bit[1299];
				Check_149 <= Bit[22] ^ Bit[80] ^ Bit[115] ^ Bit[186] ^ Bit[202] ^ Bit[268] ^ Bit[317] ^ Bit[336] ^ Bit[463] ^ Bit[697] ^ Bit[761] ^ Bit[815] ^ Bit[893] ^ Bit[941] ^ Bit[984] ^ Bit[1036] ^ Bit[1085] ^ Bit[1133] ^ Bit[1299] ^ Bit[1300];
				Check_150 <= Bit[5] ^ Bit[77] ^ Bit[117] ^ Bit[185] ^ Bit[219] ^ Bit[250] ^ Bit[303] ^ Bit[455] ^ Bit[552] ^ Bit[585] ^ Bit[789] ^ Bit[817] ^ Bit[898] ^ Bit[912] ^ Bit[995] ^ Bit[1014] ^ Bit[1078] ^ Bit[1128] ^ Bit[1300] ^ Bit[1301];
				Check_151 <= Bit[29] ^ Bit[65] ^ Bit[133] ^ Bit[146] ^ Bit[208] ^ Bit[251] ^ Bit[351] ^ Bit[405] ^ Bit[502] ^ Bit[738] ^ Bit[786] ^ Bit[834] ^ Bit[875] ^ Bit[916] ^ Bit[998] ^ Bit[1037] ^ Bit[1063] ^ Bit[1122] ^ Bit[1301] ^ Bit[1302];
				Check_152 <= Bit[38] ^ Bit[87] ^ Bit[143] ^ Bit[191] ^ Bit[220] ^ Bit[241] ^ Bit[292] ^ Bit[399] ^ Bit[488] ^ Bit[648] ^ Bit[709] ^ Bit[829] ^ Bit[871] ^ Bit[934] ^ Bit[965] ^ Bit[1045] ^ Bit[1064] ^ Bit[1143] ^ Bit[1302] ^ Bit[1303];
				Check_153 <= Bit[33] ^ Bit[60] ^ Bit[125] ^ Bit[159] ^ Bit[225] ^ Bit[244] ^ Bit[341] ^ Bit[396] ^ Bit[555] ^ Bit[612] ^ Bit[640] ^ Bit[744] ^ Bit[875] ^ Bit[919] ^ Bit[992] ^ Bit[1052] ^ Bit[1082] ^ Bit[1127] ^ Bit[1303] ^ Bit[1304];
				Check_154 <= Bit[4] ^ Bit[63] ^ Bit[102] ^ Bit[158] ^ Bit[223] ^ Bit[277] ^ Bit[453] ^ Bit[493] ^ Bit[529] ^ Bit[591] ^ Bit[664] ^ Bit[710] ^ Bit[879] ^ Bit[951] ^ Bit[987] ^ Bit[1017] ^ Bit[1092] ^ Bit[1108] ^ Bit[1304] ^ Bit[1305];
				Check_155 <= Bit[23] ^ Bit[81] ^ Bit[116] ^ Bit[187] ^ Bit[203] ^ Bit[269] ^ Bit[318] ^ Bit[337] ^ Bit[464] ^ Bit[698] ^ Bit[762] ^ Bit[768] ^ Bit[894] ^ Bit[942] ^ Bit[985] ^ Bit[1037] ^ Bit[1086] ^ Bit[1134] ^ Bit[1305] ^ Bit[1306];
				Check_156 <= Bit[6] ^ Bit[78] ^ Bit[118] ^ Bit[186] ^ Bit[220] ^ Bit[251] ^ Bit[304] ^ Bit[456] ^ Bit[553] ^ Bit[586] ^ Bit[790] ^ Bit[818] ^ Bit[899] ^ Bit[913] ^ Bit[996] ^ Bit[1015] ^ Bit[1079] ^ Bit[1129] ^ Bit[1306] ^ Bit[1307];
				Check_157 <= Bit[30] ^ Bit[66] ^ Bit[134] ^ Bit[147] ^ Bit[209] ^ Bit[252] ^ Bit[352] ^ Bit[406] ^ Bit[503] ^ Bit[739] ^ Bit[787] ^ Bit[835] ^ Bit[876] ^ Bit[917] ^ Bit[999] ^ Bit[1038] ^ Bit[1064] ^ Bit[1123] ^ Bit[1307] ^ Bit[1308];
				Check_158 <= Bit[39] ^ Bit[88] ^ Bit[96] ^ Bit[144] ^ Bit[221] ^ Bit[242] ^ Bit[293] ^ Bit[400] ^ Bit[489] ^ Bit[649] ^ Bit[710] ^ Bit[830] ^ Bit[872] ^ Bit[935] ^ Bit[966] ^ Bit[1046] ^ Bit[1065] ^ Bit[1144] ^ Bit[1308] ^ Bit[1309];
				Check_159 <= Bit[34] ^ Bit[61] ^ Bit[126] ^ Bit[160] ^ Bit[226] ^ Bit[245] ^ Bit[342] ^ Bit[397] ^ Bit[556] ^ Bit[613] ^ Bit[641] ^ Bit[745] ^ Bit[876] ^ Bit[920] ^ Bit[993] ^ Bit[1053] ^ Bit[1083] ^ Bit[1128] ^ Bit[1309] ^ Bit[1310];
				Check_160 <= Bit[5] ^ Bit[64] ^ Bit[103] ^ Bit[159] ^ Bit[224] ^ Bit[278] ^ Bit[454] ^ Bit[494] ^ Bit[530] ^ Bit[592] ^ Bit[665] ^ Bit[711] ^ Bit[880] ^ Bit[952] ^ Bit[988] ^ Bit[1018] ^ Bit[1093] ^ Bit[1109] ^ Bit[1310] ^ Bit[1311];
				Check_161 <= Bit[24] ^ Bit[82] ^ Bit[117] ^ Bit[188] ^ Bit[204] ^ Bit[270] ^ Bit[319] ^ Bit[338] ^ Bit[465] ^ Bit[699] ^ Bit[763] ^ Bit[769] ^ Bit[895] ^ Bit[943] ^ Bit[986] ^ Bit[1038] ^ Bit[1087] ^ Bit[1135] ^ Bit[1311] ^ Bit[1312];
				Check_162 <= Bit[7] ^ Bit[79] ^ Bit[119] ^ Bit[187] ^ Bit[221] ^ Bit[252] ^ Bit[305] ^ Bit[457] ^ Bit[554] ^ Bit[587] ^ Bit[791] ^ Bit[819] ^ Bit[900] ^ Bit[914] ^ Bit[997] ^ Bit[1016] ^ Bit[1080] ^ Bit[1130] ^ Bit[1312] ^ Bit[1313];
				Check_163 <= Bit[31] ^ Bit[67] ^ Bit[135] ^ Bit[148] ^ Bit[210] ^ Bit[253] ^ Bit[353] ^ Bit[407] ^ Bit[504] ^ Bit[740] ^ Bit[788] ^ Bit[836] ^ Bit[877] ^ Bit[918] ^ Bit[1000] ^ Bit[1039] ^ Bit[1065] ^ Bit[1124] ^ Bit[1313] ^ Bit[1314];
				Check_164 <= Bit[40] ^ Bit[89] ^ Bit[97] ^ Bit[145] ^ Bit[222] ^ Bit[243] ^ Bit[294] ^ Bit[401] ^ Bit[490] ^ Bit[650] ^ Bit[711] ^ Bit[831] ^ Bit[873] ^ Bit[936] ^ Bit[967] ^ Bit[1047] ^ Bit[1066] ^ Bit[1145] ^ Bit[1314] ^ Bit[1315];
				Check_165 <= Bit[35] ^ Bit[62] ^ Bit[127] ^ Bit[161] ^ Bit[227] ^ Bit[246] ^ Bit[343] ^ Bit[398] ^ Bit[557] ^ Bit[614] ^ Bit[642] ^ Bit[746] ^ Bit[877] ^ Bit[921] ^ Bit[994] ^ Bit[1054] ^ Bit[1084] ^ Bit[1129] ^ Bit[1315] ^ Bit[1316];
				Check_166 <= Bit[6] ^ Bit[65] ^ Bit[104] ^ Bit[160] ^ Bit[225] ^ Bit[279] ^ Bit[455] ^ Bit[495] ^ Bit[531] ^ Bit[593] ^ Bit[666] ^ Bit[712] ^ Bit[881] ^ Bit[953] ^ Bit[989] ^ Bit[1019] ^ Bit[1094] ^ Bit[1110] ^ Bit[1316] ^ Bit[1317];
				Check_167 <= Bit[25] ^ Bit[83] ^ Bit[118] ^ Bit[189] ^ Bit[205] ^ Bit[271] ^ Bit[320] ^ Bit[339] ^ Bit[466] ^ Bit[700] ^ Bit[764] ^ Bit[770] ^ Bit[896] ^ Bit[944] ^ Bit[987] ^ Bit[1039] ^ Bit[1088] ^ Bit[1136] ^ Bit[1317] ^ Bit[1318];
				Check_168 <= Bit[8] ^ Bit[80] ^ Bit[120] ^ Bit[188] ^ Bit[222] ^ Bit[253] ^ Bit[306] ^ Bit[458] ^ Bit[555] ^ Bit[588] ^ Bit[792] ^ Bit[820] ^ Bit[901] ^ Bit[915] ^ Bit[998] ^ Bit[1017] ^ Bit[1081] ^ Bit[1131] ^ Bit[1318] ^ Bit[1319];
				Check_169 <= Bit[32] ^ Bit[68] ^ Bit[136] ^ Bit[149] ^ Bit[211] ^ Bit[254] ^ Bit[354] ^ Bit[408] ^ Bit[505] ^ Bit[741] ^ Bit[789] ^ Bit[837] ^ Bit[878] ^ Bit[919] ^ Bit[1001] ^ Bit[1040] ^ Bit[1066] ^ Bit[1125] ^ Bit[1319] ^ Bit[1320];
				Check_170 <= Bit[41] ^ Bit[90] ^ Bit[98] ^ Bit[146] ^ Bit[223] ^ Bit[244] ^ Bit[295] ^ Bit[402] ^ Bit[491] ^ Bit[651] ^ Bit[712] ^ Bit[832] ^ Bit[874] ^ Bit[937] ^ Bit[968] ^ Bit[1048] ^ Bit[1067] ^ Bit[1146] ^ Bit[1320] ^ Bit[1321];
				Check_171 <= Bit[36] ^ Bit[63] ^ Bit[128] ^ Bit[162] ^ Bit[228] ^ Bit[247] ^ Bit[344] ^ Bit[399] ^ Bit[558] ^ Bit[615] ^ Bit[643] ^ Bit[747] ^ Bit[878] ^ Bit[922] ^ Bit[995] ^ Bit[1055] ^ Bit[1085] ^ Bit[1130] ^ Bit[1321] ^ Bit[1322];
				Check_172 <= Bit[7] ^ Bit[66] ^ Bit[105] ^ Bit[161] ^ Bit[226] ^ Bit[280] ^ Bit[456] ^ Bit[496] ^ Bit[532] ^ Bit[594] ^ Bit[667] ^ Bit[713] ^ Bit[882] ^ Bit[954] ^ Bit[990] ^ Bit[1020] ^ Bit[1095] ^ Bit[1111] ^ Bit[1322] ^ Bit[1323];
				Check_173 <= Bit[26] ^ Bit[84] ^ Bit[119] ^ Bit[190] ^ Bit[206] ^ Bit[272] ^ Bit[321] ^ Bit[340] ^ Bit[467] ^ Bit[701] ^ Bit[765] ^ Bit[771] ^ Bit[897] ^ Bit[945] ^ Bit[988] ^ Bit[1040] ^ Bit[1089] ^ Bit[1137] ^ Bit[1323] ^ Bit[1324];
				Check_174 <= Bit[9] ^ Bit[81] ^ Bit[121] ^ Bit[189] ^ Bit[223] ^ Bit[254] ^ Bit[307] ^ Bit[459] ^ Bit[556] ^ Bit[589] ^ Bit[793] ^ Bit[821] ^ Bit[902] ^ Bit[916] ^ Bit[999] ^ Bit[1018] ^ Bit[1082] ^ Bit[1132] ^ Bit[1324] ^ Bit[1325];
				Check_175 <= Bit[33] ^ Bit[69] ^ Bit[137] ^ Bit[150] ^ Bit[212] ^ Bit[255] ^ Bit[355] ^ Bit[409] ^ Bit[506] ^ Bit[742] ^ Bit[790] ^ Bit[838] ^ Bit[879] ^ Bit[920] ^ Bit[1002] ^ Bit[1041] ^ Bit[1067] ^ Bit[1126] ^ Bit[1325] ^ Bit[1326];
				Check_176 <= Bit[42] ^ Bit[91] ^ Bit[99] ^ Bit[147] ^ Bit[224] ^ Bit[245] ^ Bit[296] ^ Bit[403] ^ Bit[492] ^ Bit[652] ^ Bit[713] ^ Bit[833] ^ Bit[875] ^ Bit[938] ^ Bit[969] ^ Bit[1049] ^ Bit[1068] ^ Bit[1147] ^ Bit[1326] ^ Bit[1327];
				Check_177 <= Bit[37] ^ Bit[64] ^ Bit[129] ^ Bit[163] ^ Bit[229] ^ Bit[248] ^ Bit[345] ^ Bit[400] ^ Bit[559] ^ Bit[616] ^ Bit[644] ^ Bit[748] ^ Bit[879] ^ Bit[923] ^ Bit[996] ^ Bit[1008] ^ Bit[1086] ^ Bit[1131] ^ Bit[1327] ^ Bit[1328];
				Check_178 <= Bit[8] ^ Bit[67] ^ Bit[106] ^ Bit[162] ^ Bit[227] ^ Bit[281] ^ Bit[457] ^ Bit[497] ^ Bit[533] ^ Bit[595] ^ Bit[668] ^ Bit[714] ^ Bit[883] ^ Bit[955] ^ Bit[991] ^ Bit[1021] ^ Bit[1096] ^ Bit[1112] ^ Bit[1328] ^ Bit[1329];
				Check_179 <= Bit[27] ^ Bit[85] ^ Bit[120] ^ Bit[191] ^ Bit[207] ^ Bit[273] ^ Bit[322] ^ Bit[341] ^ Bit[468] ^ Bit[702] ^ Bit[766] ^ Bit[772] ^ Bit[898] ^ Bit[946] ^ Bit[989] ^ Bit[1041] ^ Bit[1090] ^ Bit[1138] ^ Bit[1329] ^ Bit[1330];
				Check_180 <= Bit[10] ^ Bit[82] ^ Bit[122] ^ Bit[190] ^ Bit[224] ^ Bit[255] ^ Bit[308] ^ Bit[460] ^ Bit[557] ^ Bit[590] ^ Bit[794] ^ Bit[822] ^ Bit[903] ^ Bit[917] ^ Bit[1000] ^ Bit[1019] ^ Bit[1083] ^ Bit[1133] ^ Bit[1330] ^ Bit[1331];
				Check_181 <= Bit[34] ^ Bit[70] ^ Bit[138] ^ Bit[151] ^ Bit[213] ^ Bit[256] ^ Bit[356] ^ Bit[410] ^ Bit[507] ^ Bit[743] ^ Bit[791] ^ Bit[839] ^ Bit[880] ^ Bit[921] ^ Bit[1003] ^ Bit[1042] ^ Bit[1068] ^ Bit[1127] ^ Bit[1331] ^ Bit[1332];
				Check_182 <= Bit[43] ^ Bit[92] ^ Bit[100] ^ Bit[148] ^ Bit[225] ^ Bit[246] ^ Bit[297] ^ Bit[404] ^ Bit[493] ^ Bit[653] ^ Bit[714] ^ Bit[834] ^ Bit[876] ^ Bit[939] ^ Bit[970] ^ Bit[1050] ^ Bit[1069] ^ Bit[1148] ^ Bit[1332] ^ Bit[1333];
				Check_183 <= Bit[38] ^ Bit[65] ^ Bit[130] ^ Bit[164] ^ Bit[230] ^ Bit[249] ^ Bit[346] ^ Bit[401] ^ Bit[560] ^ Bit[617] ^ Bit[645] ^ Bit[749] ^ Bit[880] ^ Bit[924] ^ Bit[997] ^ Bit[1009] ^ Bit[1087] ^ Bit[1132] ^ Bit[1333] ^ Bit[1334];
				Check_184 <= Bit[9] ^ Bit[68] ^ Bit[107] ^ Bit[163] ^ Bit[228] ^ Bit[282] ^ Bit[458] ^ Bit[498] ^ Bit[534] ^ Bit[596] ^ Bit[669] ^ Bit[715] ^ Bit[884] ^ Bit[956] ^ Bit[992] ^ Bit[1022] ^ Bit[1097] ^ Bit[1113] ^ Bit[1334] ^ Bit[1335];
				Check_185 <= Bit[28] ^ Bit[86] ^ Bit[121] ^ Bit[144] ^ Bit[208] ^ Bit[274] ^ Bit[323] ^ Bit[342] ^ Bit[469] ^ Bit[703] ^ Bit[767] ^ Bit[773] ^ Bit[899] ^ Bit[947] ^ Bit[990] ^ Bit[1042] ^ Bit[1091] ^ Bit[1139] ^ Bit[1335] ^ Bit[1336];
				Check_186 <= Bit[11] ^ Bit[83] ^ Bit[123] ^ Bit[191] ^ Bit[225] ^ Bit[256] ^ Bit[309] ^ Bit[461] ^ Bit[558] ^ Bit[591] ^ Bit[795] ^ Bit[823] ^ Bit[904] ^ Bit[918] ^ Bit[1001] ^ Bit[1020] ^ Bit[1084] ^ Bit[1134] ^ Bit[1336] ^ Bit[1337];
				Check_187 <= Bit[35] ^ Bit[71] ^ Bit[139] ^ Bit[152] ^ Bit[214] ^ Bit[257] ^ Bit[357] ^ Bit[411] ^ Bit[508] ^ Bit[744] ^ Bit[792] ^ Bit[840] ^ Bit[881] ^ Bit[922] ^ Bit[1004] ^ Bit[1043] ^ Bit[1069] ^ Bit[1128] ^ Bit[1337] ^ Bit[1338];
				Check_188 <= Bit[44] ^ Bit[93] ^ Bit[101] ^ Bit[149] ^ Bit[226] ^ Bit[247] ^ Bit[298] ^ Bit[405] ^ Bit[494] ^ Bit[654] ^ Bit[715] ^ Bit[835] ^ Bit[877] ^ Bit[940] ^ Bit[971] ^ Bit[1051] ^ Bit[1070] ^ Bit[1149] ^ Bit[1338] ^ Bit[1339];
				Check_189 <= Bit[39] ^ Bit[66] ^ Bit[131] ^ Bit[165] ^ Bit[231] ^ Bit[250] ^ Bit[347] ^ Bit[402] ^ Bit[561] ^ Bit[618] ^ Bit[646] ^ Bit[750] ^ Bit[881] ^ Bit[925] ^ Bit[998] ^ Bit[1010] ^ Bit[1088] ^ Bit[1133] ^ Bit[1339] ^ Bit[1340];
				Check_190 <= Bit[10] ^ Bit[69] ^ Bit[108] ^ Bit[164] ^ Bit[229] ^ Bit[283] ^ Bit[459] ^ Bit[499] ^ Bit[535] ^ Bit[597] ^ Bit[670] ^ Bit[716] ^ Bit[885] ^ Bit[957] ^ Bit[993] ^ Bit[1023] ^ Bit[1098] ^ Bit[1114] ^ Bit[1340] ^ Bit[1341];
				Check_191 <= Bit[29] ^ Bit[87] ^ Bit[122] ^ Bit[145] ^ Bit[209] ^ Bit[275] ^ Bit[324] ^ Bit[343] ^ Bit[470] ^ Bit[704] ^ Bit[720] ^ Bit[774] ^ Bit[900] ^ Bit[948] ^ Bit[991] ^ Bit[1043] ^ Bit[1092] ^ Bit[1140] ^ Bit[1341] ^ Bit[1342];
				Check_192 <= Bit[12] ^ Bit[84] ^ Bit[124] ^ Bit[144] ^ Bit[226] ^ Bit[257] ^ Bit[310] ^ Bit[462] ^ Bit[559] ^ Bit[592] ^ Bit[796] ^ Bit[824] ^ Bit[905] ^ Bit[919] ^ Bit[1002] ^ Bit[1021] ^ Bit[1085] ^ Bit[1135] ^ Bit[1342] ^ Bit[1343];
				Check_193 <= Bit[36] ^ Bit[72] ^ Bit[140] ^ Bit[153] ^ Bit[215] ^ Bit[258] ^ Bit[358] ^ Bit[412] ^ Bit[509] ^ Bit[745] ^ Bit[793] ^ Bit[841] ^ Bit[882] ^ Bit[923] ^ Bit[1005] ^ Bit[1044] ^ Bit[1070] ^ Bit[1129] ^ Bit[1343] ^ Bit[1344];
				Check_194 <= Bit[45] ^ Bit[94] ^ Bit[102] ^ Bit[150] ^ Bit[227] ^ Bit[248] ^ Bit[299] ^ Bit[406] ^ Bit[495] ^ Bit[655] ^ Bit[716] ^ Bit[836] ^ Bit[878] ^ Bit[941] ^ Bit[972] ^ Bit[1052] ^ Bit[1071] ^ Bit[1150] ^ Bit[1344] ^ Bit[1345];
				Check_195 <= Bit[40] ^ Bit[67] ^ Bit[132] ^ Bit[166] ^ Bit[232] ^ Bit[251] ^ Bit[348] ^ Bit[403] ^ Bit[562] ^ Bit[619] ^ Bit[647] ^ Bit[751] ^ Bit[882] ^ Bit[926] ^ Bit[999] ^ Bit[1011] ^ Bit[1089] ^ Bit[1134] ^ Bit[1345] ^ Bit[1346];
				Check_196 <= Bit[11] ^ Bit[70] ^ Bit[109] ^ Bit[165] ^ Bit[230] ^ Bit[284] ^ Bit[460] ^ Bit[500] ^ Bit[536] ^ Bit[598] ^ Bit[671] ^ Bit[717] ^ Bit[886] ^ Bit[958] ^ Bit[994] ^ Bit[1024] ^ Bit[1099] ^ Bit[1115] ^ Bit[1346] ^ Bit[1347];
				Check_197 <= Bit[30] ^ Bit[88] ^ Bit[123] ^ Bit[146] ^ Bit[210] ^ Bit[276] ^ Bit[325] ^ Bit[344] ^ Bit[471] ^ Bit[705] ^ Bit[721] ^ Bit[775] ^ Bit[901] ^ Bit[949] ^ Bit[992] ^ Bit[1044] ^ Bit[1093] ^ Bit[1141] ^ Bit[1347] ^ Bit[1348];
				Check_198 <= Bit[13] ^ Bit[85] ^ Bit[125] ^ Bit[145] ^ Bit[227] ^ Bit[258] ^ Bit[311] ^ Bit[463] ^ Bit[560] ^ Bit[593] ^ Bit[797] ^ Bit[825] ^ Bit[906] ^ Bit[920] ^ Bit[1003] ^ Bit[1022] ^ Bit[1086] ^ Bit[1136] ^ Bit[1348] ^ Bit[1349];
				Check_199 <= Bit[37] ^ Bit[73] ^ Bit[141] ^ Bit[154] ^ Bit[216] ^ Bit[259] ^ Bit[359] ^ Bit[413] ^ Bit[510] ^ Bit[746] ^ Bit[794] ^ Bit[842] ^ Bit[883] ^ Bit[924] ^ Bit[1006] ^ Bit[1045] ^ Bit[1071] ^ Bit[1130] ^ Bit[1349] ^ Bit[1350];
				Check_200 <= Bit[46] ^ Bit[95] ^ Bit[103] ^ Bit[151] ^ Bit[228] ^ Bit[249] ^ Bit[300] ^ Bit[407] ^ Bit[496] ^ Bit[656] ^ Bit[717] ^ Bit[837] ^ Bit[879] ^ Bit[942] ^ Bit[973] ^ Bit[1053] ^ Bit[1072] ^ Bit[1151] ^ Bit[1350] ^ Bit[1351];
				Check_201 <= Bit[41] ^ Bit[68] ^ Bit[133] ^ Bit[167] ^ Bit[233] ^ Bit[252] ^ Bit[349] ^ Bit[404] ^ Bit[563] ^ Bit[620] ^ Bit[648] ^ Bit[752] ^ Bit[883] ^ Bit[927] ^ Bit[1000] ^ Bit[1012] ^ Bit[1090] ^ Bit[1135] ^ Bit[1351] ^ Bit[1352];
				Check_202 <= Bit[12] ^ Bit[71] ^ Bit[110] ^ Bit[166] ^ Bit[231] ^ Bit[285] ^ Bit[461] ^ Bit[501] ^ Bit[537] ^ Bit[599] ^ Bit[624] ^ Bit[718] ^ Bit[887] ^ Bit[959] ^ Bit[995] ^ Bit[1025] ^ Bit[1100] ^ Bit[1116] ^ Bit[1352] ^ Bit[1353];
				Check_203 <= Bit[31] ^ Bit[89] ^ Bit[124] ^ Bit[147] ^ Bit[211] ^ Bit[277] ^ Bit[326] ^ Bit[345] ^ Bit[472] ^ Bit[706] ^ Bit[722] ^ Bit[776] ^ Bit[902] ^ Bit[950] ^ Bit[993] ^ Bit[1045] ^ Bit[1094] ^ Bit[1142] ^ Bit[1353] ^ Bit[1354];
				Check_204 <= Bit[14] ^ Bit[86] ^ Bit[126] ^ Bit[146] ^ Bit[228] ^ Bit[259] ^ Bit[312] ^ Bit[464] ^ Bit[561] ^ Bit[594] ^ Bit[798] ^ Bit[826] ^ Bit[907] ^ Bit[921] ^ Bit[1004] ^ Bit[1023] ^ Bit[1087] ^ Bit[1137] ^ Bit[1354] ^ Bit[1355];
				Check_205 <= Bit[38] ^ Bit[74] ^ Bit[142] ^ Bit[155] ^ Bit[217] ^ Bit[260] ^ Bit[360] ^ Bit[414] ^ Bit[511] ^ Bit[747] ^ Bit[795] ^ Bit[843] ^ Bit[884] ^ Bit[925] ^ Bit[1007] ^ Bit[1046] ^ Bit[1072] ^ Bit[1131] ^ Bit[1355] ^ Bit[1356];
				Check_206 <= Bit[47] ^ Bit[48] ^ Bit[104] ^ Bit[152] ^ Bit[229] ^ Bit[250] ^ Bit[301] ^ Bit[408] ^ Bit[497] ^ Bit[657] ^ Bit[718] ^ Bit[838] ^ Bit[880] ^ Bit[943] ^ Bit[974] ^ Bit[1054] ^ Bit[1073] ^ Bit[1104] ^ Bit[1356] ^ Bit[1357];
				Check_207 <= Bit[42] ^ Bit[69] ^ Bit[134] ^ Bit[168] ^ Bit[234] ^ Bit[253] ^ Bit[350] ^ Bit[405] ^ Bit[564] ^ Bit[621] ^ Bit[649] ^ Bit[753] ^ Bit[884] ^ Bit[928] ^ Bit[1001] ^ Bit[1013] ^ Bit[1091] ^ Bit[1136] ^ Bit[1357] ^ Bit[1358];
				Check_208 <= Bit[13] ^ Bit[72] ^ Bit[111] ^ Bit[167] ^ Bit[232] ^ Bit[286] ^ Bit[462] ^ Bit[502] ^ Bit[538] ^ Bit[600] ^ Bit[625] ^ Bit[719] ^ Bit[888] ^ Bit[912] ^ Bit[996] ^ Bit[1026] ^ Bit[1101] ^ Bit[1117] ^ Bit[1358] ^ Bit[1359];
				Check_209 <= Bit[32] ^ Bit[90] ^ Bit[125] ^ Bit[148] ^ Bit[212] ^ Bit[278] ^ Bit[327] ^ Bit[346] ^ Bit[473] ^ Bit[707] ^ Bit[723] ^ Bit[777] ^ Bit[903] ^ Bit[951] ^ Bit[994] ^ Bit[1046] ^ Bit[1095] ^ Bit[1143] ^ Bit[1359] ^ Bit[1360];
				Check_210 <= Bit[15] ^ Bit[87] ^ Bit[127] ^ Bit[147] ^ Bit[229] ^ Bit[260] ^ Bit[313] ^ Bit[465] ^ Bit[562] ^ Bit[595] ^ Bit[799] ^ Bit[827] ^ Bit[908] ^ Bit[922] ^ Bit[1005] ^ Bit[1024] ^ Bit[1088] ^ Bit[1138] ^ Bit[1360] ^ Bit[1361];
				Check_211 <= Bit[39] ^ Bit[75] ^ Bit[143] ^ Bit[156] ^ Bit[218] ^ Bit[261] ^ Bit[361] ^ Bit[415] ^ Bit[512] ^ Bit[748] ^ Bit[796] ^ Bit[844] ^ Bit[885] ^ Bit[926] ^ Bit[960] ^ Bit[1047] ^ Bit[1073] ^ Bit[1132] ^ Bit[1361] ^ Bit[1362];
				Check_212 <= Bit[0] ^ Bit[49] ^ Bit[105] ^ Bit[153] ^ Bit[230] ^ Bit[251] ^ Bit[302] ^ Bit[409] ^ Bit[498] ^ Bit[658] ^ Bit[719] ^ Bit[839] ^ Bit[881] ^ Bit[944] ^ Bit[975] ^ Bit[1055] ^ Bit[1074] ^ Bit[1105] ^ Bit[1362] ^ Bit[1363];
				Check_213 <= Bit[43] ^ Bit[70] ^ Bit[135] ^ Bit[169] ^ Bit[235] ^ Bit[254] ^ Bit[351] ^ Bit[406] ^ Bit[565] ^ Bit[622] ^ Bit[650] ^ Bit[754] ^ Bit[885] ^ Bit[929] ^ Bit[1002] ^ Bit[1014] ^ Bit[1092] ^ Bit[1137] ^ Bit[1363] ^ Bit[1364];
				Check_214 <= Bit[14] ^ Bit[73] ^ Bit[112] ^ Bit[168] ^ Bit[233] ^ Bit[287] ^ Bit[463] ^ Bit[503] ^ Bit[539] ^ Bit[601] ^ Bit[626] ^ Bit[672] ^ Bit[889] ^ Bit[913] ^ Bit[997] ^ Bit[1027] ^ Bit[1102] ^ Bit[1118] ^ Bit[1364] ^ Bit[1365];
				Check_215 <= Bit[33] ^ Bit[91] ^ Bit[126] ^ Bit[149] ^ Bit[213] ^ Bit[279] ^ Bit[328] ^ Bit[347] ^ Bit[474] ^ Bit[708] ^ Bit[724] ^ Bit[778] ^ Bit[904] ^ Bit[952] ^ Bit[995] ^ Bit[1047] ^ Bit[1096] ^ Bit[1144] ^ Bit[1365] ^ Bit[1366];
				Check_216 <= Bit[16] ^ Bit[88] ^ Bit[128] ^ Bit[148] ^ Bit[230] ^ Bit[261] ^ Bit[314] ^ Bit[466] ^ Bit[563] ^ Bit[596] ^ Bit[800] ^ Bit[828] ^ Bit[909] ^ Bit[923] ^ Bit[1006] ^ Bit[1025] ^ Bit[1089] ^ Bit[1139] ^ Bit[1366] ^ Bit[1367];
				Check_217 <= Bit[40] ^ Bit[76] ^ Bit[96] ^ Bit[157] ^ Bit[219] ^ Bit[262] ^ Bit[362] ^ Bit[416] ^ Bit[513] ^ Bit[749] ^ Bit[797] ^ Bit[845] ^ Bit[886] ^ Bit[927] ^ Bit[961] ^ Bit[1048] ^ Bit[1074] ^ Bit[1133] ^ Bit[1367] ^ Bit[1368];
				Check_218 <= Bit[1] ^ Bit[50] ^ Bit[106] ^ Bit[154] ^ Bit[231] ^ Bit[252] ^ Bit[303] ^ Bit[410] ^ Bit[499] ^ Bit[659] ^ Bit[672] ^ Bit[840] ^ Bit[882] ^ Bit[945] ^ Bit[976] ^ Bit[1008] ^ Bit[1075] ^ Bit[1106] ^ Bit[1368] ^ Bit[1369];
				Check_219 <= Bit[44] ^ Bit[71] ^ Bit[136] ^ Bit[170] ^ Bit[236] ^ Bit[255] ^ Bit[352] ^ Bit[407] ^ Bit[566] ^ Bit[623] ^ Bit[651] ^ Bit[755] ^ Bit[886] ^ Bit[930] ^ Bit[1003] ^ Bit[1015] ^ Bit[1093] ^ Bit[1138] ^ Bit[1369] ^ Bit[1370];
				Check_220 <= Bit[15] ^ Bit[74] ^ Bit[113] ^ Bit[169] ^ Bit[234] ^ Bit[240] ^ Bit[464] ^ Bit[504] ^ Bit[540] ^ Bit[602] ^ Bit[627] ^ Bit[673] ^ Bit[890] ^ Bit[914] ^ Bit[998] ^ Bit[1028] ^ Bit[1103] ^ Bit[1119] ^ Bit[1370] ^ Bit[1371];
				Check_221 <= Bit[34] ^ Bit[92] ^ Bit[127] ^ Bit[150] ^ Bit[214] ^ Bit[280] ^ Bit[329] ^ Bit[348] ^ Bit[475] ^ Bit[709] ^ Bit[725] ^ Bit[779] ^ Bit[905] ^ Bit[953] ^ Bit[996] ^ Bit[1048] ^ Bit[1097] ^ Bit[1145] ^ Bit[1371] ^ Bit[1372];
				Check_222 <= Bit[17] ^ Bit[89] ^ Bit[129] ^ Bit[149] ^ Bit[231] ^ Bit[262] ^ Bit[315] ^ Bit[467] ^ Bit[564] ^ Bit[597] ^ Bit[801] ^ Bit[829] ^ Bit[910] ^ Bit[924] ^ Bit[1007] ^ Bit[1026] ^ Bit[1090] ^ Bit[1140] ^ Bit[1372] ^ Bit[1373];
				Check_223 <= Bit[41] ^ Bit[77] ^ Bit[97] ^ Bit[158] ^ Bit[220] ^ Bit[263] ^ Bit[363] ^ Bit[417] ^ Bit[514] ^ Bit[750] ^ Bit[798] ^ Bit[846] ^ Bit[887] ^ Bit[928] ^ Bit[962] ^ Bit[1049] ^ Bit[1075] ^ Bit[1134] ^ Bit[1373] ^ Bit[1374];
				Check_224 <= Bit[2] ^ Bit[51] ^ Bit[107] ^ Bit[155] ^ Bit[232] ^ Bit[253] ^ Bit[304] ^ Bit[411] ^ Bit[500] ^ Bit[660] ^ Bit[673] ^ Bit[841] ^ Bit[883] ^ Bit[946] ^ Bit[977] ^ Bit[1009] ^ Bit[1076] ^ Bit[1107] ^ Bit[1374] ^ Bit[1375];
				Check_225 <= Bit[45] ^ Bit[72] ^ Bit[137] ^ Bit[171] ^ Bit[237] ^ Bit[256] ^ Bit[353] ^ Bit[408] ^ Bit[567] ^ Bit[576] ^ Bit[652] ^ Bit[756] ^ Bit[887] ^ Bit[931] ^ Bit[1004] ^ Bit[1016] ^ Bit[1094] ^ Bit[1139] ^ Bit[1375] ^ Bit[1376];
				Check_226 <= Bit[16] ^ Bit[75] ^ Bit[114] ^ Bit[170] ^ Bit[235] ^ Bit[241] ^ Bit[465] ^ Bit[505] ^ Bit[541] ^ Bit[603] ^ Bit[628] ^ Bit[674] ^ Bit[891] ^ Bit[915] ^ Bit[999] ^ Bit[1029] ^ Bit[1056] ^ Bit[1120] ^ Bit[1376] ^ Bit[1377];
				Check_227 <= Bit[35] ^ Bit[93] ^ Bit[128] ^ Bit[151] ^ Bit[215] ^ Bit[281] ^ Bit[330] ^ Bit[349] ^ Bit[476] ^ Bit[710] ^ Bit[726] ^ Bit[780] ^ Bit[906] ^ Bit[954] ^ Bit[997] ^ Bit[1049] ^ Bit[1098] ^ Bit[1146] ^ Bit[1377] ^ Bit[1378];
				Check_228 <= Bit[18] ^ Bit[90] ^ Bit[130] ^ Bit[150] ^ Bit[232] ^ Bit[263] ^ Bit[316] ^ Bit[468] ^ Bit[565] ^ Bit[598] ^ Bit[802] ^ Bit[830] ^ Bit[911] ^ Bit[925] ^ Bit[960] ^ Bit[1027] ^ Bit[1091] ^ Bit[1141] ^ Bit[1378] ^ Bit[1379];
				Check_229 <= Bit[42] ^ Bit[78] ^ Bit[98] ^ Bit[159] ^ Bit[221] ^ Bit[264] ^ Bit[364] ^ Bit[418] ^ Bit[515] ^ Bit[751] ^ Bit[799] ^ Bit[847] ^ Bit[888] ^ Bit[929] ^ Bit[963] ^ Bit[1050] ^ Bit[1076] ^ Bit[1135] ^ Bit[1379] ^ Bit[1380];
				Check_230 <= Bit[3] ^ Bit[52] ^ Bit[108] ^ Bit[156] ^ Bit[233] ^ Bit[254] ^ Bit[305] ^ Bit[412] ^ Bit[501] ^ Bit[661] ^ Bit[674] ^ Bit[842] ^ Bit[884] ^ Bit[947] ^ Bit[978] ^ Bit[1010] ^ Bit[1077] ^ Bit[1108] ^ Bit[1380] ^ Bit[1381];
				Check_231 <= Bit[46] ^ Bit[73] ^ Bit[138] ^ Bit[172] ^ Bit[238] ^ Bit[257] ^ Bit[354] ^ Bit[409] ^ Bit[568] ^ Bit[577] ^ Bit[653] ^ Bit[757] ^ Bit[888] ^ Bit[932] ^ Bit[1005] ^ Bit[1017] ^ Bit[1095] ^ Bit[1140] ^ Bit[1381] ^ Bit[1382];
				Check_232 <= Bit[17] ^ Bit[76] ^ Bit[115] ^ Bit[171] ^ Bit[236] ^ Bit[242] ^ Bit[466] ^ Bit[506] ^ Bit[542] ^ Bit[604] ^ Bit[629] ^ Bit[675] ^ Bit[892] ^ Bit[916] ^ Bit[1000] ^ Bit[1030] ^ Bit[1057] ^ Bit[1121] ^ Bit[1382] ^ Bit[1383];
				Check_233 <= Bit[36] ^ Bit[94] ^ Bit[129] ^ Bit[152] ^ Bit[216] ^ Bit[282] ^ Bit[331] ^ Bit[350] ^ Bit[477] ^ Bit[711] ^ Bit[727] ^ Bit[781] ^ Bit[907] ^ Bit[955] ^ Bit[998] ^ Bit[1050] ^ Bit[1099] ^ Bit[1147] ^ Bit[1383] ^ Bit[1384];
				Check_234 <= Bit[19] ^ Bit[91] ^ Bit[131] ^ Bit[151] ^ Bit[233] ^ Bit[264] ^ Bit[317] ^ Bit[469] ^ Bit[566] ^ Bit[599] ^ Bit[803] ^ Bit[831] ^ Bit[864] ^ Bit[926] ^ Bit[961] ^ Bit[1028] ^ Bit[1092] ^ Bit[1142] ^ Bit[1384] ^ Bit[1385];
				Check_235 <= Bit[43] ^ Bit[79] ^ Bit[99] ^ Bit[160] ^ Bit[222] ^ Bit[265] ^ Bit[365] ^ Bit[419] ^ Bit[516] ^ Bit[752] ^ Bit[800] ^ Bit[848] ^ Bit[889] ^ Bit[930] ^ Bit[964] ^ Bit[1051] ^ Bit[1077] ^ Bit[1136] ^ Bit[1385] ^ Bit[1386];
				Check_236 <= Bit[4] ^ Bit[53] ^ Bit[109] ^ Bit[157] ^ Bit[234] ^ Bit[255] ^ Bit[306] ^ Bit[413] ^ Bit[502] ^ Bit[662] ^ Bit[675] ^ Bit[843] ^ Bit[885] ^ Bit[948] ^ Bit[979] ^ Bit[1011] ^ Bit[1078] ^ Bit[1109] ^ Bit[1386] ^ Bit[1387];
				Check_237 <= Bit[47] ^ Bit[74] ^ Bit[139] ^ Bit[173] ^ Bit[239] ^ Bit[258] ^ Bit[355] ^ Bit[410] ^ Bit[569] ^ Bit[578] ^ Bit[654] ^ Bit[758] ^ Bit[889] ^ Bit[933] ^ Bit[1006] ^ Bit[1018] ^ Bit[1096] ^ Bit[1141] ^ Bit[1387] ^ Bit[1388];
				Check_238 <= Bit[18] ^ Bit[77] ^ Bit[116] ^ Bit[172] ^ Bit[237] ^ Bit[243] ^ Bit[467] ^ Bit[507] ^ Bit[543] ^ Bit[605] ^ Bit[630] ^ Bit[676] ^ Bit[893] ^ Bit[917] ^ Bit[1001] ^ Bit[1031] ^ Bit[1058] ^ Bit[1122] ^ Bit[1388] ^ Bit[1389];
				Check_239 <= Bit[37] ^ Bit[95] ^ Bit[130] ^ Bit[153] ^ Bit[217] ^ Bit[283] ^ Bit[332] ^ Bit[351] ^ Bit[478] ^ Bit[712] ^ Bit[728] ^ Bit[782] ^ Bit[908] ^ Bit[956] ^ Bit[999] ^ Bit[1051] ^ Bit[1100] ^ Bit[1148] ^ Bit[1389] ^ Bit[1390];
				Check_240 <= Bit[20] ^ Bit[92] ^ Bit[132] ^ Bit[152] ^ Bit[234] ^ Bit[265] ^ Bit[318] ^ Bit[470] ^ Bit[567] ^ Bit[600] ^ Bit[804] ^ Bit[832] ^ Bit[865] ^ Bit[927] ^ Bit[962] ^ Bit[1029] ^ Bit[1093] ^ Bit[1143] ^ Bit[1390] ^ Bit[1391];
				Check_241 <= Bit[44] ^ Bit[80] ^ Bit[100] ^ Bit[161] ^ Bit[223] ^ Bit[266] ^ Bit[366] ^ Bit[420] ^ Bit[517] ^ Bit[753] ^ Bit[801] ^ Bit[849] ^ Bit[890] ^ Bit[931] ^ Bit[965] ^ Bit[1052] ^ Bit[1078] ^ Bit[1137] ^ Bit[1391] ^ Bit[1392];
				Check_242 <= Bit[5] ^ Bit[54] ^ Bit[110] ^ Bit[158] ^ Bit[235] ^ Bit[256] ^ Bit[307] ^ Bit[414] ^ Bit[503] ^ Bit[663] ^ Bit[676] ^ Bit[844] ^ Bit[886] ^ Bit[949] ^ Bit[980] ^ Bit[1012] ^ Bit[1079] ^ Bit[1110] ^ Bit[1392] ^ Bit[1393];
				Check_243 <= Bit[0] ^ Bit[75] ^ Bit[140] ^ Bit[174] ^ Bit[192] ^ Bit[259] ^ Bit[356] ^ Bit[411] ^ Bit[570] ^ Bit[579] ^ Bit[655] ^ Bit[759] ^ Bit[890] ^ Bit[934] ^ Bit[1007] ^ Bit[1019] ^ Bit[1097] ^ Bit[1142] ^ Bit[1393] ^ Bit[1394];
				Check_244 <= Bit[19] ^ Bit[78] ^ Bit[117] ^ Bit[173] ^ Bit[238] ^ Bit[244] ^ Bit[468] ^ Bit[508] ^ Bit[544] ^ Bit[606] ^ Bit[631] ^ Bit[677] ^ Bit[894] ^ Bit[918] ^ Bit[1002] ^ Bit[1032] ^ Bit[1059] ^ Bit[1123] ^ Bit[1394] ^ Bit[1395];
				Check_245 <= Bit[38] ^ Bit[48] ^ Bit[131] ^ Bit[154] ^ Bit[218] ^ Bit[284] ^ Bit[333] ^ Bit[352] ^ Bit[479] ^ Bit[713] ^ Bit[729] ^ Bit[783] ^ Bit[909] ^ Bit[957] ^ Bit[1000] ^ Bit[1052] ^ Bit[1101] ^ Bit[1149] ^ Bit[1395] ^ Bit[1396];
				Check_246 <= Bit[21] ^ Bit[93] ^ Bit[133] ^ Bit[153] ^ Bit[235] ^ Bit[266] ^ Bit[319] ^ Bit[471] ^ Bit[568] ^ Bit[601] ^ Bit[805] ^ Bit[833] ^ Bit[866] ^ Bit[928] ^ Bit[963] ^ Bit[1030] ^ Bit[1094] ^ Bit[1144] ^ Bit[1396] ^ Bit[1397];
				Check_247 <= Bit[45] ^ Bit[81] ^ Bit[101] ^ Bit[162] ^ Bit[224] ^ Bit[267] ^ Bit[367] ^ Bit[421] ^ Bit[518] ^ Bit[754] ^ Bit[802] ^ Bit[850] ^ Bit[891] ^ Bit[932] ^ Bit[966] ^ Bit[1053] ^ Bit[1079] ^ Bit[1138] ^ Bit[1397] ^ Bit[1398];
				Check_248 <= Bit[6] ^ Bit[55] ^ Bit[111] ^ Bit[159] ^ Bit[236] ^ Bit[257] ^ Bit[308] ^ Bit[415] ^ Bit[504] ^ Bit[664] ^ Bit[677] ^ Bit[845] ^ Bit[887] ^ Bit[950] ^ Bit[981] ^ Bit[1013] ^ Bit[1080] ^ Bit[1111] ^ Bit[1398] ^ Bit[1399];
				Check_249 <= Bit[1] ^ Bit[76] ^ Bit[141] ^ Bit[175] ^ Bit[193] ^ Bit[260] ^ Bit[357] ^ Bit[412] ^ Bit[571] ^ Bit[580] ^ Bit[656] ^ Bit[760] ^ Bit[891] ^ Bit[935] ^ Bit[960] ^ Bit[1020] ^ Bit[1098] ^ Bit[1143] ^ Bit[1399] ^ Bit[1400];
				Check_250 <= Bit[20] ^ Bit[79] ^ Bit[118] ^ Bit[174] ^ Bit[239] ^ Bit[245] ^ Bit[469] ^ Bit[509] ^ Bit[545] ^ Bit[607] ^ Bit[632] ^ Bit[678] ^ Bit[895] ^ Bit[919] ^ Bit[1003] ^ Bit[1033] ^ Bit[1060] ^ Bit[1124] ^ Bit[1400] ^ Bit[1401];
				Check_251 <= Bit[39] ^ Bit[49] ^ Bit[132] ^ Bit[155] ^ Bit[219] ^ Bit[285] ^ Bit[334] ^ Bit[353] ^ Bit[432] ^ Bit[714] ^ Bit[730] ^ Bit[784] ^ Bit[910] ^ Bit[958] ^ Bit[1001] ^ Bit[1053] ^ Bit[1102] ^ Bit[1150] ^ Bit[1401] ^ Bit[1402];
				Check_252 <= Bit[22] ^ Bit[94] ^ Bit[134] ^ Bit[154] ^ Bit[236] ^ Bit[267] ^ Bit[320] ^ Bit[472] ^ Bit[569] ^ Bit[602] ^ Bit[806] ^ Bit[834] ^ Bit[867] ^ Bit[929] ^ Bit[964] ^ Bit[1031] ^ Bit[1095] ^ Bit[1145] ^ Bit[1402] ^ Bit[1403];
				Check_253 <= Bit[46] ^ Bit[82] ^ Bit[102] ^ Bit[163] ^ Bit[225] ^ Bit[268] ^ Bit[368] ^ Bit[422] ^ Bit[519] ^ Bit[755] ^ Bit[803] ^ Bit[851] ^ Bit[892] ^ Bit[933] ^ Bit[967] ^ Bit[1054] ^ Bit[1080] ^ Bit[1139] ^ Bit[1403] ^ Bit[1404];
				Check_254 <= Bit[7] ^ Bit[56] ^ Bit[112] ^ Bit[160] ^ Bit[237] ^ Bit[258] ^ Bit[309] ^ Bit[416] ^ Bit[505] ^ Bit[665] ^ Bit[678] ^ Bit[846] ^ Bit[888] ^ Bit[951] ^ Bit[982] ^ Bit[1014] ^ Bit[1081] ^ Bit[1112] ^ Bit[1404] ^ Bit[1405];
				Check_255 <= Bit[2] ^ Bit[77] ^ Bit[142] ^ Bit[176] ^ Bit[194] ^ Bit[261] ^ Bit[358] ^ Bit[413] ^ Bit[572] ^ Bit[581] ^ Bit[657] ^ Bit[761] ^ Bit[892] ^ Bit[936] ^ Bit[961] ^ Bit[1021] ^ Bit[1099] ^ Bit[1144] ^ Bit[1405] ^ Bit[1406];
				Check_256 <= Bit[21] ^ Bit[80] ^ Bit[119] ^ Bit[175] ^ Bit[192] ^ Bit[246] ^ Bit[470] ^ Bit[510] ^ Bit[546] ^ Bit[608] ^ Bit[633] ^ Bit[679] ^ Bit[896] ^ Bit[920] ^ Bit[1004] ^ Bit[1034] ^ Bit[1061] ^ Bit[1125] ^ Bit[1406] ^ Bit[1407];
				Check_257 <= Bit[40] ^ Bit[50] ^ Bit[133] ^ Bit[156] ^ Bit[220] ^ Bit[286] ^ Bit[335] ^ Bit[354] ^ Bit[433] ^ Bit[715] ^ Bit[731] ^ Bit[785] ^ Bit[911] ^ Bit[959] ^ Bit[1002] ^ Bit[1054] ^ Bit[1103] ^ Bit[1151] ^ Bit[1407] ^ Bit[1408];
				Check_258 <= Bit[23] ^ Bit[95] ^ Bit[135] ^ Bit[155] ^ Bit[237] ^ Bit[268] ^ Bit[321] ^ Bit[473] ^ Bit[570] ^ Bit[603] ^ Bit[807] ^ Bit[835] ^ Bit[868] ^ Bit[930] ^ Bit[965] ^ Bit[1032] ^ Bit[1096] ^ Bit[1146] ^ Bit[1408] ^ Bit[1409];
				Check_259 <= Bit[47] ^ Bit[83] ^ Bit[103] ^ Bit[164] ^ Bit[226] ^ Bit[269] ^ Bit[369] ^ Bit[423] ^ Bit[520] ^ Bit[756] ^ Bit[804] ^ Bit[852] ^ Bit[893] ^ Bit[934] ^ Bit[968] ^ Bit[1055] ^ Bit[1081] ^ Bit[1140] ^ Bit[1409] ^ Bit[1410];
				Check_260 <= Bit[8] ^ Bit[57] ^ Bit[113] ^ Bit[161] ^ Bit[238] ^ Bit[259] ^ Bit[310] ^ Bit[417] ^ Bit[506] ^ Bit[666] ^ Bit[679] ^ Bit[847] ^ Bit[889] ^ Bit[952] ^ Bit[983] ^ Bit[1015] ^ Bit[1082] ^ Bit[1113] ^ Bit[1410] ^ Bit[1411];
				Check_261 <= Bit[3] ^ Bit[78] ^ Bit[143] ^ Bit[177] ^ Bit[195] ^ Bit[262] ^ Bit[359] ^ Bit[414] ^ Bit[573] ^ Bit[582] ^ Bit[658] ^ Bit[762] ^ Bit[893] ^ Bit[937] ^ Bit[962] ^ Bit[1022] ^ Bit[1100] ^ Bit[1145] ^ Bit[1411] ^ Bit[1412];
				Check_262 <= Bit[22] ^ Bit[81] ^ Bit[120] ^ Bit[176] ^ Bit[193] ^ Bit[247] ^ Bit[471] ^ Bit[511] ^ Bit[547] ^ Bit[609] ^ Bit[634] ^ Bit[680] ^ Bit[897] ^ Bit[921] ^ Bit[1005] ^ Bit[1035] ^ Bit[1062] ^ Bit[1126] ^ Bit[1412] ^ Bit[1413];
				Check_263 <= Bit[41] ^ Bit[51] ^ Bit[134] ^ Bit[157] ^ Bit[221] ^ Bit[287] ^ Bit[288] ^ Bit[355] ^ Bit[434] ^ Bit[716] ^ Bit[732] ^ Bit[786] ^ Bit[864] ^ Bit[912] ^ Bit[1003] ^ Bit[1055] ^ Bit[1056] ^ Bit[1104] ^ Bit[1413] ^ Bit[1414];
				Check_264 <= Bit[24] ^ Bit[48] ^ Bit[136] ^ Bit[156] ^ Bit[238] ^ Bit[269] ^ Bit[322] ^ Bit[474] ^ Bit[571] ^ Bit[604] ^ Bit[808] ^ Bit[836] ^ Bit[869] ^ Bit[931] ^ Bit[966] ^ Bit[1033] ^ Bit[1097] ^ Bit[1147] ^ Bit[1414] ^ Bit[1415];
				Check_265 <= Bit[0] ^ Bit[84] ^ Bit[104] ^ Bit[165] ^ Bit[227] ^ Bit[270] ^ Bit[370] ^ Bit[424] ^ Bit[521] ^ Bit[757] ^ Bit[805] ^ Bit[853] ^ Bit[894] ^ Bit[935] ^ Bit[969] ^ Bit[1008] ^ Bit[1082] ^ Bit[1141] ^ Bit[1415] ^ Bit[1416];
				Check_266 <= Bit[9] ^ Bit[58] ^ Bit[114] ^ Bit[162] ^ Bit[239] ^ Bit[260] ^ Bit[311] ^ Bit[418] ^ Bit[507] ^ Bit[667] ^ Bit[680] ^ Bit[848] ^ Bit[890] ^ Bit[953] ^ Bit[984] ^ Bit[1016] ^ Bit[1083] ^ Bit[1114] ^ Bit[1416] ^ Bit[1417];
				Check_267 <= Bit[4] ^ Bit[79] ^ Bit[96] ^ Bit[178] ^ Bit[196] ^ Bit[263] ^ Bit[360] ^ Bit[415] ^ Bit[574] ^ Bit[583] ^ Bit[659] ^ Bit[763] ^ Bit[894] ^ Bit[938] ^ Bit[963] ^ Bit[1023] ^ Bit[1101] ^ Bit[1146] ^ Bit[1417] ^ Bit[1418];
				Check_268 <= Bit[23] ^ Bit[82] ^ Bit[121] ^ Bit[177] ^ Bit[194] ^ Bit[248] ^ Bit[472] ^ Bit[512] ^ Bit[548] ^ Bit[610] ^ Bit[635] ^ Bit[681] ^ Bit[898] ^ Bit[922] ^ Bit[1006] ^ Bit[1036] ^ Bit[1063] ^ Bit[1127] ^ Bit[1418] ^ Bit[1419];
				Check_269 <= Bit[42] ^ Bit[52] ^ Bit[135] ^ Bit[158] ^ Bit[222] ^ Bit[240] ^ Bit[289] ^ Bit[356] ^ Bit[435] ^ Bit[717] ^ Bit[733] ^ Bit[787] ^ Bit[865] ^ Bit[913] ^ Bit[1004] ^ Bit[1008] ^ Bit[1057] ^ Bit[1105] ^ Bit[1419] ^ Bit[1420];
				Check_270 <= Bit[25] ^ Bit[49] ^ Bit[137] ^ Bit[157] ^ Bit[239] ^ Bit[270] ^ Bit[323] ^ Bit[475] ^ Bit[572] ^ Bit[605] ^ Bit[809] ^ Bit[837] ^ Bit[870] ^ Bit[932] ^ Bit[967] ^ Bit[1034] ^ Bit[1098] ^ Bit[1148] ^ Bit[1420] ^ Bit[1421];
				Check_271 <= Bit[1] ^ Bit[85] ^ Bit[105] ^ Bit[166] ^ Bit[228] ^ Bit[271] ^ Bit[371] ^ Bit[425] ^ Bit[522] ^ Bit[758] ^ Bit[806] ^ Bit[854] ^ Bit[895] ^ Bit[936] ^ Bit[970] ^ Bit[1009] ^ Bit[1083] ^ Bit[1142] ^ Bit[1421] ^ Bit[1422];
				Check_272 <= Bit[10] ^ Bit[59] ^ Bit[115] ^ Bit[163] ^ Bit[192] ^ Bit[261] ^ Bit[312] ^ Bit[419] ^ Bit[508] ^ Bit[668] ^ Bit[681] ^ Bit[849] ^ Bit[891] ^ Bit[954] ^ Bit[985] ^ Bit[1017] ^ Bit[1084] ^ Bit[1115] ^ Bit[1422] ^ Bit[1423];
				Check_273 <= Bit[5] ^ Bit[80] ^ Bit[97] ^ Bit[179] ^ Bit[197] ^ Bit[264] ^ Bit[361] ^ Bit[416] ^ Bit[575] ^ Bit[584] ^ Bit[660] ^ Bit[764] ^ Bit[895] ^ Bit[939] ^ Bit[964] ^ Bit[1024] ^ Bit[1102] ^ Bit[1147] ^ Bit[1423] ^ Bit[1424];
				Check_274 <= Bit[24] ^ Bit[83] ^ Bit[122] ^ Bit[178] ^ Bit[195] ^ Bit[249] ^ Bit[473] ^ Bit[513] ^ Bit[549] ^ Bit[611] ^ Bit[636] ^ Bit[682] ^ Bit[899] ^ Bit[923] ^ Bit[1007] ^ Bit[1037] ^ Bit[1064] ^ Bit[1128] ^ Bit[1424] ^ Bit[1425];
				Check_275 <= Bit[43] ^ Bit[53] ^ Bit[136] ^ Bit[159] ^ Bit[223] ^ Bit[241] ^ Bit[290] ^ Bit[357] ^ Bit[436] ^ Bit[718] ^ Bit[734] ^ Bit[788] ^ Bit[866] ^ Bit[914] ^ Bit[1005] ^ Bit[1009] ^ Bit[1058] ^ Bit[1106] ^ Bit[1425] ^ Bit[1426];
				Check_276 <= Bit[26] ^ Bit[50] ^ Bit[138] ^ Bit[158] ^ Bit[192] ^ Bit[271] ^ Bit[324] ^ Bit[476] ^ Bit[573] ^ Bit[606] ^ Bit[810] ^ Bit[838] ^ Bit[871] ^ Bit[933] ^ Bit[968] ^ Bit[1035] ^ Bit[1099] ^ Bit[1149] ^ Bit[1426] ^ Bit[1427];
				Check_277 <= Bit[2] ^ Bit[86] ^ Bit[106] ^ Bit[167] ^ Bit[229] ^ Bit[272] ^ Bit[372] ^ Bit[426] ^ Bit[523] ^ Bit[759] ^ Bit[807] ^ Bit[855] ^ Bit[896] ^ Bit[937] ^ Bit[971] ^ Bit[1010] ^ Bit[1084] ^ Bit[1143] ^ Bit[1427] ^ Bit[1428];
				Check_278 <= Bit[11] ^ Bit[60] ^ Bit[116] ^ Bit[164] ^ Bit[193] ^ Bit[262] ^ Bit[313] ^ Bit[420] ^ Bit[509] ^ Bit[669] ^ Bit[682] ^ Bit[850] ^ Bit[892] ^ Bit[955] ^ Bit[986] ^ Bit[1018] ^ Bit[1085] ^ Bit[1116] ^ Bit[1428] ^ Bit[1429];
				Check_279 <= Bit[6] ^ Bit[81] ^ Bit[98] ^ Bit[180] ^ Bit[198] ^ Bit[265] ^ Bit[362] ^ Bit[417] ^ Bit[528] ^ Bit[585] ^ Bit[661] ^ Bit[765] ^ Bit[896] ^ Bit[940] ^ Bit[965] ^ Bit[1025] ^ Bit[1103] ^ Bit[1148] ^ Bit[1429] ^ Bit[1430];
				Check_280 <= Bit[25] ^ Bit[84] ^ Bit[123] ^ Bit[179] ^ Bit[196] ^ Bit[250] ^ Bit[474] ^ Bit[514] ^ Bit[550] ^ Bit[612] ^ Bit[637] ^ Bit[683] ^ Bit[900] ^ Bit[924] ^ Bit[960] ^ Bit[1038] ^ Bit[1065] ^ Bit[1129] ^ Bit[1430] ^ Bit[1431];
				Check_281 <= Bit[44] ^ Bit[54] ^ Bit[137] ^ Bit[160] ^ Bit[224] ^ Bit[242] ^ Bit[291] ^ Bit[358] ^ Bit[437] ^ Bit[719] ^ Bit[735] ^ Bit[789] ^ Bit[867] ^ Bit[915] ^ Bit[1006] ^ Bit[1010] ^ Bit[1059] ^ Bit[1107] ^ Bit[1431] ^ Bit[1432];
				Check_282 <= Bit[27] ^ Bit[51] ^ Bit[139] ^ Bit[159] ^ Bit[193] ^ Bit[272] ^ Bit[325] ^ Bit[477] ^ Bit[574] ^ Bit[607] ^ Bit[811] ^ Bit[839] ^ Bit[872] ^ Bit[934] ^ Bit[969] ^ Bit[1036] ^ Bit[1100] ^ Bit[1150] ^ Bit[1432] ^ Bit[1433];
				Check_283 <= Bit[3] ^ Bit[87] ^ Bit[107] ^ Bit[168] ^ Bit[230] ^ Bit[273] ^ Bit[373] ^ Bit[427] ^ Bit[524] ^ Bit[760] ^ Bit[808] ^ Bit[856] ^ Bit[897] ^ Bit[938] ^ Bit[972] ^ Bit[1011] ^ Bit[1085] ^ Bit[1144] ^ Bit[1433] ^ Bit[1434];
				Check_284 <= Bit[12] ^ Bit[61] ^ Bit[117] ^ Bit[165] ^ Bit[194] ^ Bit[263] ^ Bit[314] ^ Bit[421] ^ Bit[510] ^ Bit[670] ^ Bit[683] ^ Bit[851] ^ Bit[893] ^ Bit[956] ^ Bit[987] ^ Bit[1019] ^ Bit[1086] ^ Bit[1117] ^ Bit[1434] ^ Bit[1435];
				Check_285 <= Bit[7] ^ Bit[82] ^ Bit[99] ^ Bit[181] ^ Bit[199] ^ Bit[266] ^ Bit[363] ^ Bit[418] ^ Bit[529] ^ Bit[586] ^ Bit[662] ^ Bit[766] ^ Bit[897] ^ Bit[941] ^ Bit[966] ^ Bit[1026] ^ Bit[1056] ^ Bit[1149] ^ Bit[1435] ^ Bit[1436];
				Check_286 <= Bit[26] ^ Bit[85] ^ Bit[124] ^ Bit[180] ^ Bit[197] ^ Bit[251] ^ Bit[475] ^ Bit[515] ^ Bit[551] ^ Bit[613] ^ Bit[638] ^ Bit[684] ^ Bit[901] ^ Bit[925] ^ Bit[961] ^ Bit[1039] ^ Bit[1066] ^ Bit[1130] ^ Bit[1436] ^ Bit[1437];
				Check_287 <= Bit[45] ^ Bit[55] ^ Bit[138] ^ Bit[161] ^ Bit[225] ^ Bit[243] ^ Bit[292] ^ Bit[359] ^ Bit[438] ^ Bit[672] ^ Bit[736] ^ Bit[790] ^ Bit[868] ^ Bit[916] ^ Bit[1007] ^ Bit[1011] ^ Bit[1060] ^ Bit[1108] ^ Bit[1437] ^ Bit[1438];
				Check_288 <= Bit[28] ^ Bit[52] ^ Bit[140] ^ Bit[160] ^ Bit[194] ^ Bit[273] ^ Bit[326] ^ Bit[478] ^ Bit[575] ^ Bit[608] ^ Bit[812] ^ Bit[840] ^ Bit[873] ^ Bit[935] ^ Bit[970] ^ Bit[1037] ^ Bit[1101] ^ Bit[1151] ^ Bit[1438] ^ Bit[1439];
				cnt <= cnt + 1;
			end
			else if (cnt == 8'd16) begin
				Check_Sum <= Check_1 | Check_2 | Check_3 | Check_4 | Check_5 | Check_6 | Check_7 | Check_8 | Check_9 | Check_10 | Check_11 | Check_12 | Check_13 | Check_14 | Check_15 | Check_16 | Check_17 | Check_18 | Check_19 | Check_20 | Check_21 | Check_22 | Check_23 | Check_24 | Check_25 | Check_26 | Check_27 | Check_28 | Check_29 | Check_30 | Check_31 | Check_32 | Check_33 | Check_34 | Check_35 | Check_36 | Check_37 | Check_38 | Check_39 | Check_40 | Check_41 | Check_42 | Check_43 | Check_44 | Check_45 | Check_46 | Check_47 | Check_48 | Check_49 | Check_50 | Check_51 | Check_52 | Check_53 | Check_54 | Check_55 | Check_56 | Check_57 | Check_58 | Check_59 | Check_60 | Check_61 | Check_62 | Check_63 | Check_64 | Check_65 | Check_66 | Check_67 | Check_68 | Check_69 | Check_70 | Check_71 | Check_72 | Check_73 | Check_74 | Check_75 | Check_76 | Check_77 | Check_78 | Check_79 | Check_80 | Check_81 | Check_82 | Check_83 | Check_84 | Check_85 | Check_86 | Check_87 | Check_88 | Check_89 | Check_90 | Check_91 | Check_92 | Check_93 | Check_94 | Check_95 | Check_96 | Check_97 | Check_98 | Check_99 | Check_100 | Check_101 | Check_102 | Check_103 | Check_104 | Check_105 | Check_106 | Check_107 | Check_108 | Check_109 | Check_110 | Check_111 | Check_112 | Check_113 | Check_114 | Check_115 | Check_116 | Check_117 | Check_118 | Check_119 | Check_120 | Check_121 | Check_122 | Check_123 | Check_124 | Check_125 | Check_126 | Check_127 | Check_128 | Check_129 | Check_130 | Check_131 | Check_132 | Check_133 | Check_134 | Check_135 | Check_136 | Check_137 | Check_138 | Check_139 | Check_140 | Check_141 | Check_142 | Check_143 | Check_144 | Check_145 | Check_146 | Check_147 | Check_148 | Check_149 | Check_150 | Check_151 | Check_152 | Check_153 | Check_154 | Check_155 | Check_156 | Check_157 | Check_158 | Check_159 | Check_160 | Check_161 | Check_162 | Check_163 | Check_164 | Check_165 | Check_166 | Check_167 | Check_168 | Check_169 | Check_170 | Check_171 | Check_172 | Check_173 | Check_174 | Check_175 | Check_176 | Check_177 | Check_178 | Check_179 | Check_180 | Check_181 | Check_182 | Check_183 | Check_184 | Check_185 | Check_186 | Check_187 | Check_188 | Check_189 | Check_190 | Check_191 | Check_192 | Check_193 | Check_194 | Check_195 | Check_196 | Check_197 | Check_198 | Check_199 | Check_200 | Check_201 | Check_202 | Check_203 | Check_204 | Check_205 | Check_206 | Check_207 | Check_208 | Check_209 | Check_210 | Check_211 | Check_212 | Check_213 | Check_214 | Check_215 | Check_216 | Check_217 | Check_218 | Check_219 | Check_220 | Check_221 | Check_222 | Check_223 | Check_224 | Check_225 | Check_226 | Check_227 | Check_228 | Check_229 | Check_230 | Check_231 | Check_232 | Check_233 | Check_234 | Check_235 | Check_236 | Check_237 | Check_238 | Check_239 | Check_240 | Check_241 | Check_242 | Check_243 | Check_244 | Check_245 | Check_246 | Check_247 | Check_248 | Check_249 | Check_250 | Check_251 | Check_252 | Check_253 | Check_254 | Check_255 | Check_256 | Check_257 | Check_258 | Check_259 | Check_260 | Check_261 | Check_262 | Check_263 | Check_264 | Check_265 | Check_266 | Check_267 | Check_268 | Check_269 | Check_270 | Check_271 | Check_272 | Check_273 | Check_274 | Check_275 | Check_276 | Check_277 | Check_278 | Check_279 | Check_280 | Check_281 | Check_282 | Check_283 | Check_284 | Check_285 | Check_286 | Check_287 | Check_288;
				cnt <= cnt + 1;
			end
			else if (cnt == 8'd17) begin
				if (Check_Sum == 0 || iter == 5'd30) begin
					cnt <= cnt + 1;
					out_valid <= 1;
				end
				else begin
					out_valid <= 0;
					cnt <= 2;
					iter <= iter + 1;
				end
			end
		end
	end
end
assign Bit[0] = V_1[quan_width-1];
assign Bit[1] = V_2[quan_width-1];
assign Bit[2] = V_3[quan_width-1];
assign Bit[3] = V_4[quan_width-1];
assign Bit[4] = V_5[quan_width-1];
assign Bit[5] = V_6[quan_width-1];
assign Bit[6] = V_7[quan_width-1];
assign Bit[7] = V_8[quan_width-1];
assign Bit[8] = V_9[quan_width-1];
assign Bit[9] = V_10[quan_width-1];
assign Bit[10] = V_11[quan_width-1];
assign Bit[11] = V_12[quan_width-1];
assign Bit[12] = V_13[quan_width-1];
assign Bit[13] = V_14[quan_width-1];
assign Bit[14] = V_15[quan_width-1];
assign Bit[15] = V_16[quan_width-1];
assign Bit[16] = V_17[quan_width-1];
assign Bit[17] = V_18[quan_width-1];
assign Bit[18] = V_19[quan_width-1];
assign Bit[19] = V_20[quan_width-1];
assign Bit[20] = V_21[quan_width-1];
assign Bit[21] = V_22[quan_width-1];
assign Bit[22] = V_23[quan_width-1];
assign Bit[23] = V_24[quan_width-1];
assign Bit[24] = V_25[quan_width-1];
assign Bit[25] = V_26[quan_width-1];
assign Bit[26] = V_27[quan_width-1];
assign Bit[27] = V_28[quan_width-1];
assign Bit[28] = V_29[quan_width-1];
assign Bit[29] = V_30[quan_width-1];
assign Bit[30] = V_31[quan_width-1];
assign Bit[31] = V_32[quan_width-1];
assign Bit[32] = V_33[quan_width-1];
assign Bit[33] = V_34[quan_width-1];
assign Bit[34] = V_35[quan_width-1];
assign Bit[35] = V_36[quan_width-1];
assign Bit[36] = V_37[quan_width-1];
assign Bit[37] = V_38[quan_width-1];
assign Bit[38] = V_39[quan_width-1];
assign Bit[39] = V_40[quan_width-1];
assign Bit[40] = V_41[quan_width-1];
assign Bit[41] = V_42[quan_width-1];
assign Bit[42] = V_43[quan_width-1];
assign Bit[43] = V_44[quan_width-1];
assign Bit[44] = V_45[quan_width-1];
assign Bit[45] = V_46[quan_width-1];
assign Bit[46] = V_47[quan_width-1];
assign Bit[47] = V_48[quan_width-1];
assign Bit[48] = V_49[quan_width-1];
assign Bit[49] = V_50[quan_width-1];
assign Bit[50] = V_51[quan_width-1];
assign Bit[51] = V_52[quan_width-1];
assign Bit[52] = V_53[quan_width-1];
assign Bit[53] = V_54[quan_width-1];
assign Bit[54] = V_55[quan_width-1];
assign Bit[55] = V_56[quan_width-1];
assign Bit[56] = V_57[quan_width-1];
assign Bit[57] = V_58[quan_width-1];
assign Bit[58] = V_59[quan_width-1];
assign Bit[59] = V_60[quan_width-1];
assign Bit[60] = V_61[quan_width-1];
assign Bit[61] = V_62[quan_width-1];
assign Bit[62] = V_63[quan_width-1];
assign Bit[63] = V_64[quan_width-1];
assign Bit[64] = V_65[quan_width-1];
assign Bit[65] = V_66[quan_width-1];
assign Bit[66] = V_67[quan_width-1];
assign Bit[67] = V_68[quan_width-1];
assign Bit[68] = V_69[quan_width-1];
assign Bit[69] = V_70[quan_width-1];
assign Bit[70] = V_71[quan_width-1];
assign Bit[71] = V_72[quan_width-1];
assign Bit[72] = V_73[quan_width-1];
assign Bit[73] = V_74[quan_width-1];
assign Bit[74] = V_75[quan_width-1];
assign Bit[75] = V_76[quan_width-1];
assign Bit[76] = V_77[quan_width-1];
assign Bit[77] = V_78[quan_width-1];
assign Bit[78] = V_79[quan_width-1];
assign Bit[79] = V_80[quan_width-1];
assign Bit[80] = V_81[quan_width-1];
assign Bit[81] = V_82[quan_width-1];
assign Bit[82] = V_83[quan_width-1];
assign Bit[83] = V_84[quan_width-1];
assign Bit[84] = V_85[quan_width-1];
assign Bit[85] = V_86[quan_width-1];
assign Bit[86] = V_87[quan_width-1];
assign Bit[87] = V_88[quan_width-1];
assign Bit[88] = V_89[quan_width-1];
assign Bit[89] = V_90[quan_width-1];
assign Bit[90] = V_91[quan_width-1];
assign Bit[91] = V_92[quan_width-1];
assign Bit[92] = V_93[quan_width-1];
assign Bit[93] = V_94[quan_width-1];
assign Bit[94] = V_95[quan_width-1];
assign Bit[95] = V_96[quan_width-1];
assign Bit[96] = V_97[quan_width-1];
assign Bit[97] = V_98[quan_width-1];
assign Bit[98] = V_99[quan_width-1];
assign Bit[99] = V_100[quan_width-1];
assign Bit[100] = V_101[quan_width-1];
assign Bit[101] = V_102[quan_width-1];
assign Bit[102] = V_103[quan_width-1];
assign Bit[103] = V_104[quan_width-1];
assign Bit[104] = V_105[quan_width-1];
assign Bit[105] = V_106[quan_width-1];
assign Bit[106] = V_107[quan_width-1];
assign Bit[107] = V_108[quan_width-1];
assign Bit[108] = V_109[quan_width-1];
assign Bit[109] = V_110[quan_width-1];
assign Bit[110] = V_111[quan_width-1];
assign Bit[111] = V_112[quan_width-1];
assign Bit[112] = V_113[quan_width-1];
assign Bit[113] = V_114[quan_width-1];
assign Bit[114] = V_115[quan_width-1];
assign Bit[115] = V_116[quan_width-1];
assign Bit[116] = V_117[quan_width-1];
assign Bit[117] = V_118[quan_width-1];
assign Bit[118] = V_119[quan_width-1];
assign Bit[119] = V_120[quan_width-1];
assign Bit[120] = V_121[quan_width-1];
assign Bit[121] = V_122[quan_width-1];
assign Bit[122] = V_123[quan_width-1];
assign Bit[123] = V_124[quan_width-1];
assign Bit[124] = V_125[quan_width-1];
assign Bit[125] = V_126[quan_width-1];
assign Bit[126] = V_127[quan_width-1];
assign Bit[127] = V_128[quan_width-1];
assign Bit[128] = V_129[quan_width-1];
assign Bit[129] = V_130[quan_width-1];
assign Bit[130] = V_131[quan_width-1];
assign Bit[131] = V_132[quan_width-1];
assign Bit[132] = V_133[quan_width-1];
assign Bit[133] = V_134[quan_width-1];
assign Bit[134] = V_135[quan_width-1];
assign Bit[135] = V_136[quan_width-1];
assign Bit[136] = V_137[quan_width-1];
assign Bit[137] = V_138[quan_width-1];
assign Bit[138] = V_139[quan_width-1];
assign Bit[139] = V_140[quan_width-1];
assign Bit[140] = V_141[quan_width-1];
assign Bit[141] = V_142[quan_width-1];
assign Bit[142] = V_143[quan_width-1];
assign Bit[143] = V_144[quan_width-1];
assign Bit[144] = V_145[quan_width-1];
assign Bit[145] = V_146[quan_width-1];
assign Bit[146] = V_147[quan_width-1];
assign Bit[147] = V_148[quan_width-1];
assign Bit[148] = V_149[quan_width-1];
assign Bit[149] = V_150[quan_width-1];
assign Bit[150] = V_151[quan_width-1];
assign Bit[151] = V_152[quan_width-1];
assign Bit[152] = V_153[quan_width-1];
assign Bit[153] = V_154[quan_width-1];
assign Bit[154] = V_155[quan_width-1];
assign Bit[155] = V_156[quan_width-1];
assign Bit[156] = V_157[quan_width-1];
assign Bit[157] = V_158[quan_width-1];
assign Bit[158] = V_159[quan_width-1];
assign Bit[159] = V_160[quan_width-1];
assign Bit[160] = V_161[quan_width-1];
assign Bit[161] = V_162[quan_width-1];
assign Bit[162] = V_163[quan_width-1];
assign Bit[163] = V_164[quan_width-1];
assign Bit[164] = V_165[quan_width-1];
assign Bit[165] = V_166[quan_width-1];
assign Bit[166] = V_167[quan_width-1];
assign Bit[167] = V_168[quan_width-1];
assign Bit[168] = V_169[quan_width-1];
assign Bit[169] = V_170[quan_width-1];
assign Bit[170] = V_171[quan_width-1];
assign Bit[171] = V_172[quan_width-1];
assign Bit[172] = V_173[quan_width-1];
assign Bit[173] = V_174[quan_width-1];
assign Bit[174] = V_175[quan_width-1];
assign Bit[175] = V_176[quan_width-1];
assign Bit[176] = V_177[quan_width-1];
assign Bit[177] = V_178[quan_width-1];
assign Bit[178] = V_179[quan_width-1];
assign Bit[179] = V_180[quan_width-1];
assign Bit[180] = V_181[quan_width-1];
assign Bit[181] = V_182[quan_width-1];
assign Bit[182] = V_183[quan_width-1];
assign Bit[183] = V_184[quan_width-1];
assign Bit[184] = V_185[quan_width-1];
assign Bit[185] = V_186[quan_width-1];
assign Bit[186] = V_187[quan_width-1];
assign Bit[187] = V_188[quan_width-1];
assign Bit[188] = V_189[quan_width-1];
assign Bit[189] = V_190[quan_width-1];
assign Bit[190] = V_191[quan_width-1];
assign Bit[191] = V_192[quan_width-1];
assign Bit[192] = V_193[quan_width-1];
assign Bit[193] = V_194[quan_width-1];
assign Bit[194] = V_195[quan_width-1];
assign Bit[195] = V_196[quan_width-1];
assign Bit[196] = V_197[quan_width-1];
assign Bit[197] = V_198[quan_width-1];
assign Bit[198] = V_199[quan_width-1];
assign Bit[199] = V_200[quan_width-1];
assign Bit[200] = V_201[quan_width-1];
assign Bit[201] = V_202[quan_width-1];
assign Bit[202] = V_203[quan_width-1];
assign Bit[203] = V_204[quan_width-1];
assign Bit[204] = V_205[quan_width-1];
assign Bit[205] = V_206[quan_width-1];
assign Bit[206] = V_207[quan_width-1];
assign Bit[207] = V_208[quan_width-1];
assign Bit[208] = V_209[quan_width-1];
assign Bit[209] = V_210[quan_width-1];
assign Bit[210] = V_211[quan_width-1];
assign Bit[211] = V_212[quan_width-1];
assign Bit[212] = V_213[quan_width-1];
assign Bit[213] = V_214[quan_width-1];
assign Bit[214] = V_215[quan_width-1];
assign Bit[215] = V_216[quan_width-1];
assign Bit[216] = V_217[quan_width-1];
assign Bit[217] = V_218[quan_width-1];
assign Bit[218] = V_219[quan_width-1];
assign Bit[219] = V_220[quan_width-1];
assign Bit[220] = V_221[quan_width-1];
assign Bit[221] = V_222[quan_width-1];
assign Bit[222] = V_223[quan_width-1];
assign Bit[223] = V_224[quan_width-1];
assign Bit[224] = V_225[quan_width-1];
assign Bit[225] = V_226[quan_width-1];
assign Bit[226] = V_227[quan_width-1];
assign Bit[227] = V_228[quan_width-1];
assign Bit[228] = V_229[quan_width-1];
assign Bit[229] = V_230[quan_width-1];
assign Bit[230] = V_231[quan_width-1];
assign Bit[231] = V_232[quan_width-1];
assign Bit[232] = V_233[quan_width-1];
assign Bit[233] = V_234[quan_width-1];
assign Bit[234] = V_235[quan_width-1];
assign Bit[235] = V_236[quan_width-1];
assign Bit[236] = V_237[quan_width-1];
assign Bit[237] = V_238[quan_width-1];
assign Bit[238] = V_239[quan_width-1];
assign Bit[239] = V_240[quan_width-1];
assign Bit[240] = V_241[quan_width-1];
assign Bit[241] = V_242[quan_width-1];
assign Bit[242] = V_243[quan_width-1];
assign Bit[243] = V_244[quan_width-1];
assign Bit[244] = V_245[quan_width-1];
assign Bit[245] = V_246[quan_width-1];
assign Bit[246] = V_247[quan_width-1];
assign Bit[247] = V_248[quan_width-1];
assign Bit[248] = V_249[quan_width-1];
assign Bit[249] = V_250[quan_width-1];
assign Bit[250] = V_251[quan_width-1];
assign Bit[251] = V_252[quan_width-1];
assign Bit[252] = V_253[quan_width-1];
assign Bit[253] = V_254[quan_width-1];
assign Bit[254] = V_255[quan_width-1];
assign Bit[255] = V_256[quan_width-1];
assign Bit[256] = V_257[quan_width-1];
assign Bit[257] = V_258[quan_width-1];
assign Bit[258] = V_259[quan_width-1];
assign Bit[259] = V_260[quan_width-1];
assign Bit[260] = V_261[quan_width-1];
assign Bit[261] = V_262[quan_width-1];
assign Bit[262] = V_263[quan_width-1];
assign Bit[263] = V_264[quan_width-1];
assign Bit[264] = V_265[quan_width-1];
assign Bit[265] = V_266[quan_width-1];
assign Bit[266] = V_267[quan_width-1];
assign Bit[267] = V_268[quan_width-1];
assign Bit[268] = V_269[quan_width-1];
assign Bit[269] = V_270[quan_width-1];
assign Bit[270] = V_271[quan_width-1];
assign Bit[271] = V_272[quan_width-1];
assign Bit[272] = V_273[quan_width-1];
assign Bit[273] = V_274[quan_width-1];
assign Bit[274] = V_275[quan_width-1];
assign Bit[275] = V_276[quan_width-1];
assign Bit[276] = V_277[quan_width-1];
assign Bit[277] = V_278[quan_width-1];
assign Bit[278] = V_279[quan_width-1];
assign Bit[279] = V_280[quan_width-1];
assign Bit[280] = V_281[quan_width-1];
assign Bit[281] = V_282[quan_width-1];
assign Bit[282] = V_283[quan_width-1];
assign Bit[283] = V_284[quan_width-1];
assign Bit[284] = V_285[quan_width-1];
assign Bit[285] = V_286[quan_width-1];
assign Bit[286] = V_287[quan_width-1];
assign Bit[287] = V_288[quan_width-1];
assign Bit[288] = V_289[quan_width-1];
assign Bit[289] = V_290[quan_width-1];
assign Bit[290] = V_291[quan_width-1];
assign Bit[291] = V_292[quan_width-1];
assign Bit[292] = V_293[quan_width-1];
assign Bit[293] = V_294[quan_width-1];
assign Bit[294] = V_295[quan_width-1];
assign Bit[295] = V_296[quan_width-1];
assign Bit[296] = V_297[quan_width-1];
assign Bit[297] = V_298[quan_width-1];
assign Bit[298] = V_299[quan_width-1];
assign Bit[299] = V_300[quan_width-1];
assign Bit[300] = V_301[quan_width-1];
assign Bit[301] = V_302[quan_width-1];
assign Bit[302] = V_303[quan_width-1];
assign Bit[303] = V_304[quan_width-1];
assign Bit[304] = V_305[quan_width-1];
assign Bit[305] = V_306[quan_width-1];
assign Bit[306] = V_307[quan_width-1];
assign Bit[307] = V_308[quan_width-1];
assign Bit[308] = V_309[quan_width-1];
assign Bit[309] = V_310[quan_width-1];
assign Bit[310] = V_311[quan_width-1];
assign Bit[311] = V_312[quan_width-1];
assign Bit[312] = V_313[quan_width-1];
assign Bit[313] = V_314[quan_width-1];
assign Bit[314] = V_315[quan_width-1];
assign Bit[315] = V_316[quan_width-1];
assign Bit[316] = V_317[quan_width-1];
assign Bit[317] = V_318[quan_width-1];
assign Bit[318] = V_319[quan_width-1];
assign Bit[319] = V_320[quan_width-1];
assign Bit[320] = V_321[quan_width-1];
assign Bit[321] = V_322[quan_width-1];
assign Bit[322] = V_323[quan_width-1];
assign Bit[323] = V_324[quan_width-1];
assign Bit[324] = V_325[quan_width-1];
assign Bit[325] = V_326[quan_width-1];
assign Bit[326] = V_327[quan_width-1];
assign Bit[327] = V_328[quan_width-1];
assign Bit[328] = V_329[quan_width-1];
assign Bit[329] = V_330[quan_width-1];
assign Bit[330] = V_331[quan_width-1];
assign Bit[331] = V_332[quan_width-1];
assign Bit[332] = V_333[quan_width-1];
assign Bit[333] = V_334[quan_width-1];
assign Bit[334] = V_335[quan_width-1];
assign Bit[335] = V_336[quan_width-1];
assign Bit[336] = V_337[quan_width-1];
assign Bit[337] = V_338[quan_width-1];
assign Bit[338] = V_339[quan_width-1];
assign Bit[339] = V_340[quan_width-1];
assign Bit[340] = V_341[quan_width-1];
assign Bit[341] = V_342[quan_width-1];
assign Bit[342] = V_343[quan_width-1];
assign Bit[343] = V_344[quan_width-1];
assign Bit[344] = V_345[quan_width-1];
assign Bit[345] = V_346[quan_width-1];
assign Bit[346] = V_347[quan_width-1];
assign Bit[347] = V_348[quan_width-1];
assign Bit[348] = V_349[quan_width-1];
assign Bit[349] = V_350[quan_width-1];
assign Bit[350] = V_351[quan_width-1];
assign Bit[351] = V_352[quan_width-1];
assign Bit[352] = V_353[quan_width-1];
assign Bit[353] = V_354[quan_width-1];
assign Bit[354] = V_355[quan_width-1];
assign Bit[355] = V_356[quan_width-1];
assign Bit[356] = V_357[quan_width-1];
assign Bit[357] = V_358[quan_width-1];
assign Bit[358] = V_359[quan_width-1];
assign Bit[359] = V_360[quan_width-1];
assign Bit[360] = V_361[quan_width-1];
assign Bit[361] = V_362[quan_width-1];
assign Bit[362] = V_363[quan_width-1];
assign Bit[363] = V_364[quan_width-1];
assign Bit[364] = V_365[quan_width-1];
assign Bit[365] = V_366[quan_width-1];
assign Bit[366] = V_367[quan_width-1];
assign Bit[367] = V_368[quan_width-1];
assign Bit[368] = V_369[quan_width-1];
assign Bit[369] = V_370[quan_width-1];
assign Bit[370] = V_371[quan_width-1];
assign Bit[371] = V_372[quan_width-1];
assign Bit[372] = V_373[quan_width-1];
assign Bit[373] = V_374[quan_width-1];
assign Bit[374] = V_375[quan_width-1];
assign Bit[375] = V_376[quan_width-1];
assign Bit[376] = V_377[quan_width-1];
assign Bit[377] = V_378[quan_width-1];
assign Bit[378] = V_379[quan_width-1];
assign Bit[379] = V_380[quan_width-1];
assign Bit[380] = V_381[quan_width-1];
assign Bit[381] = V_382[quan_width-1];
assign Bit[382] = V_383[quan_width-1];
assign Bit[383] = V_384[quan_width-1];
assign Bit[384] = V_385[quan_width-1];
assign Bit[385] = V_386[quan_width-1];
assign Bit[386] = V_387[quan_width-1];
assign Bit[387] = V_388[quan_width-1];
assign Bit[388] = V_389[quan_width-1];
assign Bit[389] = V_390[quan_width-1];
assign Bit[390] = V_391[quan_width-1];
assign Bit[391] = V_392[quan_width-1];
assign Bit[392] = V_393[quan_width-1];
assign Bit[393] = V_394[quan_width-1];
assign Bit[394] = V_395[quan_width-1];
assign Bit[395] = V_396[quan_width-1];
assign Bit[396] = V_397[quan_width-1];
assign Bit[397] = V_398[quan_width-1];
assign Bit[398] = V_399[quan_width-1];
assign Bit[399] = V_400[quan_width-1];
assign Bit[400] = V_401[quan_width-1];
assign Bit[401] = V_402[quan_width-1];
assign Bit[402] = V_403[quan_width-1];
assign Bit[403] = V_404[quan_width-1];
assign Bit[404] = V_405[quan_width-1];
assign Bit[405] = V_406[quan_width-1];
assign Bit[406] = V_407[quan_width-1];
assign Bit[407] = V_408[quan_width-1];
assign Bit[408] = V_409[quan_width-1];
assign Bit[409] = V_410[quan_width-1];
assign Bit[410] = V_411[quan_width-1];
assign Bit[411] = V_412[quan_width-1];
assign Bit[412] = V_413[quan_width-1];
assign Bit[413] = V_414[quan_width-1];
assign Bit[414] = V_415[quan_width-1];
assign Bit[415] = V_416[quan_width-1];
assign Bit[416] = V_417[quan_width-1];
assign Bit[417] = V_418[quan_width-1];
assign Bit[418] = V_419[quan_width-1];
assign Bit[419] = V_420[quan_width-1];
assign Bit[420] = V_421[quan_width-1];
assign Bit[421] = V_422[quan_width-1];
assign Bit[422] = V_423[quan_width-1];
assign Bit[423] = V_424[quan_width-1];
assign Bit[424] = V_425[quan_width-1];
assign Bit[425] = V_426[quan_width-1];
assign Bit[426] = V_427[quan_width-1];
assign Bit[427] = V_428[quan_width-1];
assign Bit[428] = V_429[quan_width-1];
assign Bit[429] = V_430[quan_width-1];
assign Bit[430] = V_431[quan_width-1];
assign Bit[431] = V_432[quan_width-1];
assign Bit[432] = V_433[quan_width-1];
assign Bit[433] = V_434[quan_width-1];
assign Bit[434] = V_435[quan_width-1];
assign Bit[435] = V_436[quan_width-1];
assign Bit[436] = V_437[quan_width-1];
assign Bit[437] = V_438[quan_width-1];
assign Bit[438] = V_439[quan_width-1];
assign Bit[439] = V_440[quan_width-1];
assign Bit[440] = V_441[quan_width-1];
assign Bit[441] = V_442[quan_width-1];
assign Bit[442] = V_443[quan_width-1];
assign Bit[443] = V_444[quan_width-1];
assign Bit[444] = V_445[quan_width-1];
assign Bit[445] = V_446[quan_width-1];
assign Bit[446] = V_447[quan_width-1];
assign Bit[447] = V_448[quan_width-1];
assign Bit[448] = V_449[quan_width-1];
assign Bit[449] = V_450[quan_width-1];
assign Bit[450] = V_451[quan_width-1];
assign Bit[451] = V_452[quan_width-1];
assign Bit[452] = V_453[quan_width-1];
assign Bit[453] = V_454[quan_width-1];
assign Bit[454] = V_455[quan_width-1];
assign Bit[455] = V_456[quan_width-1];
assign Bit[456] = V_457[quan_width-1];
assign Bit[457] = V_458[quan_width-1];
assign Bit[458] = V_459[quan_width-1];
assign Bit[459] = V_460[quan_width-1];
assign Bit[460] = V_461[quan_width-1];
assign Bit[461] = V_462[quan_width-1];
assign Bit[462] = V_463[quan_width-1];
assign Bit[463] = V_464[quan_width-1];
assign Bit[464] = V_465[quan_width-1];
assign Bit[465] = V_466[quan_width-1];
assign Bit[466] = V_467[quan_width-1];
assign Bit[467] = V_468[quan_width-1];
assign Bit[468] = V_469[quan_width-1];
assign Bit[469] = V_470[quan_width-1];
assign Bit[470] = V_471[quan_width-1];
assign Bit[471] = V_472[quan_width-1];
assign Bit[472] = V_473[quan_width-1];
assign Bit[473] = V_474[quan_width-1];
assign Bit[474] = V_475[quan_width-1];
assign Bit[475] = V_476[quan_width-1];
assign Bit[476] = V_477[quan_width-1];
assign Bit[477] = V_478[quan_width-1];
assign Bit[478] = V_479[quan_width-1];
assign Bit[479] = V_480[quan_width-1];
assign Bit[480] = V_481[quan_width-1];
assign Bit[481] = V_482[quan_width-1];
assign Bit[482] = V_483[quan_width-1];
assign Bit[483] = V_484[quan_width-1];
assign Bit[484] = V_485[quan_width-1];
assign Bit[485] = V_486[quan_width-1];
assign Bit[486] = V_487[quan_width-1];
assign Bit[487] = V_488[quan_width-1];
assign Bit[488] = V_489[quan_width-1];
assign Bit[489] = V_490[quan_width-1];
assign Bit[490] = V_491[quan_width-1];
assign Bit[491] = V_492[quan_width-1];
assign Bit[492] = V_493[quan_width-1];
assign Bit[493] = V_494[quan_width-1];
assign Bit[494] = V_495[quan_width-1];
assign Bit[495] = V_496[quan_width-1];
assign Bit[496] = V_497[quan_width-1];
assign Bit[497] = V_498[quan_width-1];
assign Bit[498] = V_499[quan_width-1];
assign Bit[499] = V_500[quan_width-1];
assign Bit[500] = V_501[quan_width-1];
assign Bit[501] = V_502[quan_width-1];
assign Bit[502] = V_503[quan_width-1];
assign Bit[503] = V_504[quan_width-1];
assign Bit[504] = V_505[quan_width-1];
assign Bit[505] = V_506[quan_width-1];
assign Bit[506] = V_507[quan_width-1];
assign Bit[507] = V_508[quan_width-1];
assign Bit[508] = V_509[quan_width-1];
assign Bit[509] = V_510[quan_width-1];
assign Bit[510] = V_511[quan_width-1];
assign Bit[511] = V_512[quan_width-1];
assign Bit[512] = V_513[quan_width-1];
assign Bit[513] = V_514[quan_width-1];
assign Bit[514] = V_515[quan_width-1];
assign Bit[515] = V_516[quan_width-1];
assign Bit[516] = V_517[quan_width-1];
assign Bit[517] = V_518[quan_width-1];
assign Bit[518] = V_519[quan_width-1];
assign Bit[519] = V_520[quan_width-1];
assign Bit[520] = V_521[quan_width-1];
assign Bit[521] = V_522[quan_width-1];
assign Bit[522] = V_523[quan_width-1];
assign Bit[523] = V_524[quan_width-1];
assign Bit[524] = V_525[quan_width-1];
assign Bit[525] = V_526[quan_width-1];
assign Bit[526] = V_527[quan_width-1];
assign Bit[527] = V_528[quan_width-1];
assign Bit[528] = V_529[quan_width-1];
assign Bit[529] = V_530[quan_width-1];
assign Bit[530] = V_531[quan_width-1];
assign Bit[531] = V_532[quan_width-1];
assign Bit[532] = V_533[quan_width-1];
assign Bit[533] = V_534[quan_width-1];
assign Bit[534] = V_535[quan_width-1];
assign Bit[535] = V_536[quan_width-1];
assign Bit[536] = V_537[quan_width-1];
assign Bit[537] = V_538[quan_width-1];
assign Bit[538] = V_539[quan_width-1];
assign Bit[539] = V_540[quan_width-1];
assign Bit[540] = V_541[quan_width-1];
assign Bit[541] = V_542[quan_width-1];
assign Bit[542] = V_543[quan_width-1];
assign Bit[543] = V_544[quan_width-1];
assign Bit[544] = V_545[quan_width-1];
assign Bit[545] = V_546[quan_width-1];
assign Bit[546] = V_547[quan_width-1];
assign Bit[547] = V_548[quan_width-1];
assign Bit[548] = V_549[quan_width-1];
assign Bit[549] = V_550[quan_width-1];
assign Bit[550] = V_551[quan_width-1];
assign Bit[551] = V_552[quan_width-1];
assign Bit[552] = V_553[quan_width-1];
assign Bit[553] = V_554[quan_width-1];
assign Bit[554] = V_555[quan_width-1];
assign Bit[555] = V_556[quan_width-1];
assign Bit[556] = V_557[quan_width-1];
assign Bit[557] = V_558[quan_width-1];
assign Bit[558] = V_559[quan_width-1];
assign Bit[559] = V_560[quan_width-1];
assign Bit[560] = V_561[quan_width-1];
assign Bit[561] = V_562[quan_width-1];
assign Bit[562] = V_563[quan_width-1];
assign Bit[563] = V_564[quan_width-1];
assign Bit[564] = V_565[quan_width-1];
assign Bit[565] = V_566[quan_width-1];
assign Bit[566] = V_567[quan_width-1];
assign Bit[567] = V_568[quan_width-1];
assign Bit[568] = V_569[quan_width-1];
assign Bit[569] = V_570[quan_width-1];
assign Bit[570] = V_571[quan_width-1];
assign Bit[571] = V_572[quan_width-1];
assign Bit[572] = V_573[quan_width-1];
assign Bit[573] = V_574[quan_width-1];
assign Bit[574] = V_575[quan_width-1];
assign Bit[575] = V_576[quan_width-1];
assign Bit[576] = V_577[quan_width-1];
assign Bit[577] = V_578[quan_width-1];
assign Bit[578] = V_579[quan_width-1];
assign Bit[579] = V_580[quan_width-1];
assign Bit[580] = V_581[quan_width-1];
assign Bit[581] = V_582[quan_width-1];
assign Bit[582] = V_583[quan_width-1];
assign Bit[583] = V_584[quan_width-1];
assign Bit[584] = V_585[quan_width-1];
assign Bit[585] = V_586[quan_width-1];
assign Bit[586] = V_587[quan_width-1];
assign Bit[587] = V_588[quan_width-1];
assign Bit[588] = V_589[quan_width-1];
assign Bit[589] = V_590[quan_width-1];
assign Bit[590] = V_591[quan_width-1];
assign Bit[591] = V_592[quan_width-1];
assign Bit[592] = V_593[quan_width-1];
assign Bit[593] = V_594[quan_width-1];
assign Bit[594] = V_595[quan_width-1];
assign Bit[595] = V_596[quan_width-1];
assign Bit[596] = V_597[quan_width-1];
assign Bit[597] = V_598[quan_width-1];
assign Bit[598] = V_599[quan_width-1];
assign Bit[599] = V_600[quan_width-1];
assign Bit[600] = V_601[quan_width-1];
assign Bit[601] = V_602[quan_width-1];
assign Bit[602] = V_603[quan_width-1];
assign Bit[603] = V_604[quan_width-1];
assign Bit[604] = V_605[quan_width-1];
assign Bit[605] = V_606[quan_width-1];
assign Bit[606] = V_607[quan_width-1];
assign Bit[607] = V_608[quan_width-1];
assign Bit[608] = V_609[quan_width-1];
assign Bit[609] = V_610[quan_width-1];
assign Bit[610] = V_611[quan_width-1];
assign Bit[611] = V_612[quan_width-1];
assign Bit[612] = V_613[quan_width-1];
assign Bit[613] = V_614[quan_width-1];
assign Bit[614] = V_615[quan_width-1];
assign Bit[615] = V_616[quan_width-1];
assign Bit[616] = V_617[quan_width-1];
assign Bit[617] = V_618[quan_width-1];
assign Bit[618] = V_619[quan_width-1];
assign Bit[619] = V_620[quan_width-1];
assign Bit[620] = V_621[quan_width-1];
assign Bit[621] = V_622[quan_width-1];
assign Bit[622] = V_623[quan_width-1];
assign Bit[623] = V_624[quan_width-1];
assign Bit[624] = V_625[quan_width-1];
assign Bit[625] = V_626[quan_width-1];
assign Bit[626] = V_627[quan_width-1];
assign Bit[627] = V_628[quan_width-1];
assign Bit[628] = V_629[quan_width-1];
assign Bit[629] = V_630[quan_width-1];
assign Bit[630] = V_631[quan_width-1];
assign Bit[631] = V_632[quan_width-1];
assign Bit[632] = V_633[quan_width-1];
assign Bit[633] = V_634[quan_width-1];
assign Bit[634] = V_635[quan_width-1];
assign Bit[635] = V_636[quan_width-1];
assign Bit[636] = V_637[quan_width-1];
assign Bit[637] = V_638[quan_width-1];
assign Bit[638] = V_639[quan_width-1];
assign Bit[639] = V_640[quan_width-1];
assign Bit[640] = V_641[quan_width-1];
assign Bit[641] = V_642[quan_width-1];
assign Bit[642] = V_643[quan_width-1];
assign Bit[643] = V_644[quan_width-1];
assign Bit[644] = V_645[quan_width-1];
assign Bit[645] = V_646[quan_width-1];
assign Bit[646] = V_647[quan_width-1];
assign Bit[647] = V_648[quan_width-1];
assign Bit[648] = V_649[quan_width-1];
assign Bit[649] = V_650[quan_width-1];
assign Bit[650] = V_651[quan_width-1];
assign Bit[651] = V_652[quan_width-1];
assign Bit[652] = V_653[quan_width-1];
assign Bit[653] = V_654[quan_width-1];
assign Bit[654] = V_655[quan_width-1];
assign Bit[655] = V_656[quan_width-1];
assign Bit[656] = V_657[quan_width-1];
assign Bit[657] = V_658[quan_width-1];
assign Bit[658] = V_659[quan_width-1];
assign Bit[659] = V_660[quan_width-1];
assign Bit[660] = V_661[quan_width-1];
assign Bit[661] = V_662[quan_width-1];
assign Bit[662] = V_663[quan_width-1];
assign Bit[663] = V_664[quan_width-1];
assign Bit[664] = V_665[quan_width-1];
assign Bit[665] = V_666[quan_width-1];
assign Bit[666] = V_667[quan_width-1];
assign Bit[667] = V_668[quan_width-1];
assign Bit[668] = V_669[quan_width-1];
assign Bit[669] = V_670[quan_width-1];
assign Bit[670] = V_671[quan_width-1];
assign Bit[671] = V_672[quan_width-1];
assign Bit[672] = V_673[quan_width-1];
assign Bit[673] = V_674[quan_width-1];
assign Bit[674] = V_675[quan_width-1];
assign Bit[675] = V_676[quan_width-1];
assign Bit[676] = V_677[quan_width-1];
assign Bit[677] = V_678[quan_width-1];
assign Bit[678] = V_679[quan_width-1];
assign Bit[679] = V_680[quan_width-1];
assign Bit[680] = V_681[quan_width-1];
assign Bit[681] = V_682[quan_width-1];
assign Bit[682] = V_683[quan_width-1];
assign Bit[683] = V_684[quan_width-1];
assign Bit[684] = V_685[quan_width-1];
assign Bit[685] = V_686[quan_width-1];
assign Bit[686] = V_687[quan_width-1];
assign Bit[687] = V_688[quan_width-1];
assign Bit[688] = V_689[quan_width-1];
assign Bit[689] = V_690[quan_width-1];
assign Bit[690] = V_691[quan_width-1];
assign Bit[691] = V_692[quan_width-1];
assign Bit[692] = V_693[quan_width-1];
assign Bit[693] = V_694[quan_width-1];
assign Bit[694] = V_695[quan_width-1];
assign Bit[695] = V_696[quan_width-1];
assign Bit[696] = V_697[quan_width-1];
assign Bit[697] = V_698[quan_width-1];
assign Bit[698] = V_699[quan_width-1];
assign Bit[699] = V_700[quan_width-1];
assign Bit[700] = V_701[quan_width-1];
assign Bit[701] = V_702[quan_width-1];
assign Bit[702] = V_703[quan_width-1];
assign Bit[703] = V_704[quan_width-1];
assign Bit[704] = V_705[quan_width-1];
assign Bit[705] = V_706[quan_width-1];
assign Bit[706] = V_707[quan_width-1];
assign Bit[707] = V_708[quan_width-1];
assign Bit[708] = V_709[quan_width-1];
assign Bit[709] = V_710[quan_width-1];
assign Bit[710] = V_711[quan_width-1];
assign Bit[711] = V_712[quan_width-1];
assign Bit[712] = V_713[quan_width-1];
assign Bit[713] = V_714[quan_width-1];
assign Bit[714] = V_715[quan_width-1];
assign Bit[715] = V_716[quan_width-1];
assign Bit[716] = V_717[quan_width-1];
assign Bit[717] = V_718[quan_width-1];
assign Bit[718] = V_719[quan_width-1];
assign Bit[719] = V_720[quan_width-1];
assign Bit[720] = V_721[quan_width-1];
assign Bit[721] = V_722[quan_width-1];
assign Bit[722] = V_723[quan_width-1];
assign Bit[723] = V_724[quan_width-1];
assign Bit[724] = V_725[quan_width-1];
assign Bit[725] = V_726[quan_width-1];
assign Bit[726] = V_727[quan_width-1];
assign Bit[727] = V_728[quan_width-1];
assign Bit[728] = V_729[quan_width-1];
assign Bit[729] = V_730[quan_width-1];
assign Bit[730] = V_731[quan_width-1];
assign Bit[731] = V_732[quan_width-1];
assign Bit[732] = V_733[quan_width-1];
assign Bit[733] = V_734[quan_width-1];
assign Bit[734] = V_735[quan_width-1];
assign Bit[735] = V_736[quan_width-1];
assign Bit[736] = V_737[quan_width-1];
assign Bit[737] = V_738[quan_width-1];
assign Bit[738] = V_739[quan_width-1];
assign Bit[739] = V_740[quan_width-1];
assign Bit[740] = V_741[quan_width-1];
assign Bit[741] = V_742[quan_width-1];
assign Bit[742] = V_743[quan_width-1];
assign Bit[743] = V_744[quan_width-1];
assign Bit[744] = V_745[quan_width-1];
assign Bit[745] = V_746[quan_width-1];
assign Bit[746] = V_747[quan_width-1];
assign Bit[747] = V_748[quan_width-1];
assign Bit[748] = V_749[quan_width-1];
assign Bit[749] = V_750[quan_width-1];
assign Bit[750] = V_751[quan_width-1];
assign Bit[751] = V_752[quan_width-1];
assign Bit[752] = V_753[quan_width-1];
assign Bit[753] = V_754[quan_width-1];
assign Bit[754] = V_755[quan_width-1];
assign Bit[755] = V_756[quan_width-1];
assign Bit[756] = V_757[quan_width-1];
assign Bit[757] = V_758[quan_width-1];
assign Bit[758] = V_759[quan_width-1];
assign Bit[759] = V_760[quan_width-1];
assign Bit[760] = V_761[quan_width-1];
assign Bit[761] = V_762[quan_width-1];
assign Bit[762] = V_763[quan_width-1];
assign Bit[763] = V_764[quan_width-1];
assign Bit[764] = V_765[quan_width-1];
assign Bit[765] = V_766[quan_width-1];
assign Bit[766] = V_767[quan_width-1];
assign Bit[767] = V_768[quan_width-1];
assign Bit[768] = V_769[quan_width-1];
assign Bit[769] = V_770[quan_width-1];
assign Bit[770] = V_771[quan_width-1];
assign Bit[771] = V_772[quan_width-1];
assign Bit[772] = V_773[quan_width-1];
assign Bit[773] = V_774[quan_width-1];
assign Bit[774] = V_775[quan_width-1];
assign Bit[775] = V_776[quan_width-1];
assign Bit[776] = V_777[quan_width-1];
assign Bit[777] = V_778[quan_width-1];
assign Bit[778] = V_779[quan_width-1];
assign Bit[779] = V_780[quan_width-1];
assign Bit[780] = V_781[quan_width-1];
assign Bit[781] = V_782[quan_width-1];
assign Bit[782] = V_783[quan_width-1];
assign Bit[783] = V_784[quan_width-1];
assign Bit[784] = V_785[quan_width-1];
assign Bit[785] = V_786[quan_width-1];
assign Bit[786] = V_787[quan_width-1];
assign Bit[787] = V_788[quan_width-1];
assign Bit[788] = V_789[quan_width-1];
assign Bit[789] = V_790[quan_width-1];
assign Bit[790] = V_791[quan_width-1];
assign Bit[791] = V_792[quan_width-1];
assign Bit[792] = V_793[quan_width-1];
assign Bit[793] = V_794[quan_width-1];
assign Bit[794] = V_795[quan_width-1];
assign Bit[795] = V_796[quan_width-1];
assign Bit[796] = V_797[quan_width-1];
assign Bit[797] = V_798[quan_width-1];
assign Bit[798] = V_799[quan_width-1];
assign Bit[799] = V_800[quan_width-1];
assign Bit[800] = V_801[quan_width-1];
assign Bit[801] = V_802[quan_width-1];
assign Bit[802] = V_803[quan_width-1];
assign Bit[803] = V_804[quan_width-1];
assign Bit[804] = V_805[quan_width-1];
assign Bit[805] = V_806[quan_width-1];
assign Bit[806] = V_807[quan_width-1];
assign Bit[807] = V_808[quan_width-1];
assign Bit[808] = V_809[quan_width-1];
assign Bit[809] = V_810[quan_width-1];
assign Bit[810] = V_811[quan_width-1];
assign Bit[811] = V_812[quan_width-1];
assign Bit[812] = V_813[quan_width-1];
assign Bit[813] = V_814[quan_width-1];
assign Bit[814] = V_815[quan_width-1];
assign Bit[815] = V_816[quan_width-1];
assign Bit[816] = V_817[quan_width-1];
assign Bit[817] = V_818[quan_width-1];
assign Bit[818] = V_819[quan_width-1];
assign Bit[819] = V_820[quan_width-1];
assign Bit[820] = V_821[quan_width-1];
assign Bit[821] = V_822[quan_width-1];
assign Bit[822] = V_823[quan_width-1];
assign Bit[823] = V_824[quan_width-1];
assign Bit[824] = V_825[quan_width-1];
assign Bit[825] = V_826[quan_width-1];
assign Bit[826] = V_827[quan_width-1];
assign Bit[827] = V_828[quan_width-1];
assign Bit[828] = V_829[quan_width-1];
assign Bit[829] = V_830[quan_width-1];
assign Bit[830] = V_831[quan_width-1];
assign Bit[831] = V_832[quan_width-1];
assign Bit[832] = V_833[quan_width-1];
assign Bit[833] = V_834[quan_width-1];
assign Bit[834] = V_835[quan_width-1];
assign Bit[835] = V_836[quan_width-1];
assign Bit[836] = V_837[quan_width-1];
assign Bit[837] = V_838[quan_width-1];
assign Bit[838] = V_839[quan_width-1];
assign Bit[839] = V_840[quan_width-1];
assign Bit[840] = V_841[quan_width-1];
assign Bit[841] = V_842[quan_width-1];
assign Bit[842] = V_843[quan_width-1];
assign Bit[843] = V_844[quan_width-1];
assign Bit[844] = V_845[quan_width-1];
assign Bit[845] = V_846[quan_width-1];
assign Bit[846] = V_847[quan_width-1];
assign Bit[847] = V_848[quan_width-1];
assign Bit[848] = V_849[quan_width-1];
assign Bit[849] = V_850[quan_width-1];
assign Bit[850] = V_851[quan_width-1];
assign Bit[851] = V_852[quan_width-1];
assign Bit[852] = V_853[quan_width-1];
assign Bit[853] = V_854[quan_width-1];
assign Bit[854] = V_855[quan_width-1];
assign Bit[855] = V_856[quan_width-1];
assign Bit[856] = V_857[quan_width-1];
assign Bit[857] = V_858[quan_width-1];
assign Bit[858] = V_859[quan_width-1];
assign Bit[859] = V_860[quan_width-1];
assign Bit[860] = V_861[quan_width-1];
assign Bit[861] = V_862[quan_width-1];
assign Bit[862] = V_863[quan_width-1];
assign Bit[863] = V_864[quan_width-1];
assign Bit[864] = V_865[quan_width-1];
assign Bit[865] = V_866[quan_width-1];
assign Bit[866] = V_867[quan_width-1];
assign Bit[867] = V_868[quan_width-1];
assign Bit[868] = V_869[quan_width-1];
assign Bit[869] = V_870[quan_width-1];
assign Bit[870] = V_871[quan_width-1];
assign Bit[871] = V_872[quan_width-1];
assign Bit[872] = V_873[quan_width-1];
assign Bit[873] = V_874[quan_width-1];
assign Bit[874] = V_875[quan_width-1];
assign Bit[875] = V_876[quan_width-1];
assign Bit[876] = V_877[quan_width-1];
assign Bit[877] = V_878[quan_width-1];
assign Bit[878] = V_879[quan_width-1];
assign Bit[879] = V_880[quan_width-1];
assign Bit[880] = V_881[quan_width-1];
assign Bit[881] = V_882[quan_width-1];
assign Bit[882] = V_883[quan_width-1];
assign Bit[883] = V_884[quan_width-1];
assign Bit[884] = V_885[quan_width-1];
assign Bit[885] = V_886[quan_width-1];
assign Bit[886] = V_887[quan_width-1];
assign Bit[887] = V_888[quan_width-1];
assign Bit[888] = V_889[quan_width-1];
assign Bit[889] = V_890[quan_width-1];
assign Bit[890] = V_891[quan_width-1];
assign Bit[891] = V_892[quan_width-1];
assign Bit[892] = V_893[quan_width-1];
assign Bit[893] = V_894[quan_width-1];
assign Bit[894] = V_895[quan_width-1];
assign Bit[895] = V_896[quan_width-1];
assign Bit[896] = V_897[quan_width-1];
assign Bit[897] = V_898[quan_width-1];
assign Bit[898] = V_899[quan_width-1];
assign Bit[899] = V_900[quan_width-1];
assign Bit[900] = V_901[quan_width-1];
assign Bit[901] = V_902[quan_width-1];
assign Bit[902] = V_903[quan_width-1];
assign Bit[903] = V_904[quan_width-1];
assign Bit[904] = V_905[quan_width-1];
assign Bit[905] = V_906[quan_width-1];
assign Bit[906] = V_907[quan_width-1];
assign Bit[907] = V_908[quan_width-1];
assign Bit[908] = V_909[quan_width-1];
assign Bit[909] = V_910[quan_width-1];
assign Bit[910] = V_911[quan_width-1];
assign Bit[911] = V_912[quan_width-1];
assign Bit[912] = V_913[quan_width-1];
assign Bit[913] = V_914[quan_width-1];
assign Bit[914] = V_915[quan_width-1];
assign Bit[915] = V_916[quan_width-1];
assign Bit[916] = V_917[quan_width-1];
assign Bit[917] = V_918[quan_width-1];
assign Bit[918] = V_919[quan_width-1];
assign Bit[919] = V_920[quan_width-1];
assign Bit[920] = V_921[quan_width-1];
assign Bit[921] = V_922[quan_width-1];
assign Bit[922] = V_923[quan_width-1];
assign Bit[923] = V_924[quan_width-1];
assign Bit[924] = V_925[quan_width-1];
assign Bit[925] = V_926[quan_width-1];
assign Bit[926] = V_927[quan_width-1];
assign Bit[927] = V_928[quan_width-1];
assign Bit[928] = V_929[quan_width-1];
assign Bit[929] = V_930[quan_width-1];
assign Bit[930] = V_931[quan_width-1];
assign Bit[931] = V_932[quan_width-1];
assign Bit[932] = V_933[quan_width-1];
assign Bit[933] = V_934[quan_width-1];
assign Bit[934] = V_935[quan_width-1];
assign Bit[935] = V_936[quan_width-1];
assign Bit[936] = V_937[quan_width-1];
assign Bit[937] = V_938[quan_width-1];
assign Bit[938] = V_939[quan_width-1];
assign Bit[939] = V_940[quan_width-1];
assign Bit[940] = V_941[quan_width-1];
assign Bit[941] = V_942[quan_width-1];
assign Bit[942] = V_943[quan_width-1];
assign Bit[943] = V_944[quan_width-1];
assign Bit[944] = V_945[quan_width-1];
assign Bit[945] = V_946[quan_width-1];
assign Bit[946] = V_947[quan_width-1];
assign Bit[947] = V_948[quan_width-1];
assign Bit[948] = V_949[quan_width-1];
assign Bit[949] = V_950[quan_width-1];
assign Bit[950] = V_951[quan_width-1];
assign Bit[951] = V_952[quan_width-1];
assign Bit[952] = V_953[quan_width-1];
assign Bit[953] = V_954[quan_width-1];
assign Bit[954] = V_955[quan_width-1];
assign Bit[955] = V_956[quan_width-1];
assign Bit[956] = V_957[quan_width-1];
assign Bit[957] = V_958[quan_width-1];
assign Bit[958] = V_959[quan_width-1];
assign Bit[959] = V_960[quan_width-1];
assign Bit[960] = V_961[quan_width-1];
assign Bit[961] = V_962[quan_width-1];
assign Bit[962] = V_963[quan_width-1];
assign Bit[963] = V_964[quan_width-1];
assign Bit[964] = V_965[quan_width-1];
assign Bit[965] = V_966[quan_width-1];
assign Bit[966] = V_967[quan_width-1];
assign Bit[967] = V_968[quan_width-1];
assign Bit[968] = V_969[quan_width-1];
assign Bit[969] = V_970[quan_width-1];
assign Bit[970] = V_971[quan_width-1];
assign Bit[971] = V_972[quan_width-1];
assign Bit[972] = V_973[quan_width-1];
assign Bit[973] = V_974[quan_width-1];
assign Bit[974] = V_975[quan_width-1];
assign Bit[975] = V_976[quan_width-1];
assign Bit[976] = V_977[quan_width-1];
assign Bit[977] = V_978[quan_width-1];
assign Bit[978] = V_979[quan_width-1];
assign Bit[979] = V_980[quan_width-1];
assign Bit[980] = V_981[quan_width-1];
assign Bit[981] = V_982[quan_width-1];
assign Bit[982] = V_983[quan_width-1];
assign Bit[983] = V_984[quan_width-1];
assign Bit[984] = V_985[quan_width-1];
assign Bit[985] = V_986[quan_width-1];
assign Bit[986] = V_987[quan_width-1];
assign Bit[987] = V_988[quan_width-1];
assign Bit[988] = V_989[quan_width-1];
assign Bit[989] = V_990[quan_width-1];
assign Bit[990] = V_991[quan_width-1];
assign Bit[991] = V_992[quan_width-1];
assign Bit[992] = V_993[quan_width-1];
assign Bit[993] = V_994[quan_width-1];
assign Bit[994] = V_995[quan_width-1];
assign Bit[995] = V_996[quan_width-1];
assign Bit[996] = V_997[quan_width-1];
assign Bit[997] = V_998[quan_width-1];
assign Bit[998] = V_999[quan_width-1];
assign Bit[999] = V_1000[quan_width-1];
assign Bit[1000] = V_1001[quan_width-1];
assign Bit[1001] = V_1002[quan_width-1];
assign Bit[1002] = V_1003[quan_width-1];
assign Bit[1003] = V_1004[quan_width-1];
assign Bit[1004] = V_1005[quan_width-1];
assign Bit[1005] = V_1006[quan_width-1];
assign Bit[1006] = V_1007[quan_width-1];
assign Bit[1007] = V_1008[quan_width-1];
assign Bit[1008] = V_1009[quan_width-1];
assign Bit[1009] = V_1010[quan_width-1];
assign Bit[1010] = V_1011[quan_width-1];
assign Bit[1011] = V_1012[quan_width-1];
assign Bit[1012] = V_1013[quan_width-1];
assign Bit[1013] = V_1014[quan_width-1];
assign Bit[1014] = V_1015[quan_width-1];
assign Bit[1015] = V_1016[quan_width-1];
assign Bit[1016] = V_1017[quan_width-1];
assign Bit[1017] = V_1018[quan_width-1];
assign Bit[1018] = V_1019[quan_width-1];
assign Bit[1019] = V_1020[quan_width-1];
assign Bit[1020] = V_1021[quan_width-1];
assign Bit[1021] = V_1022[quan_width-1];
assign Bit[1022] = V_1023[quan_width-1];
assign Bit[1023] = V_1024[quan_width-1];
assign Bit[1024] = V_1025[quan_width-1];
assign Bit[1025] = V_1026[quan_width-1];
assign Bit[1026] = V_1027[quan_width-1];
assign Bit[1027] = V_1028[quan_width-1];
assign Bit[1028] = V_1029[quan_width-1];
assign Bit[1029] = V_1030[quan_width-1];
assign Bit[1030] = V_1031[quan_width-1];
assign Bit[1031] = V_1032[quan_width-1];
assign Bit[1032] = V_1033[quan_width-1];
assign Bit[1033] = V_1034[quan_width-1];
assign Bit[1034] = V_1035[quan_width-1];
assign Bit[1035] = V_1036[quan_width-1];
assign Bit[1036] = V_1037[quan_width-1];
assign Bit[1037] = V_1038[quan_width-1];
assign Bit[1038] = V_1039[quan_width-1];
assign Bit[1039] = V_1040[quan_width-1];
assign Bit[1040] = V_1041[quan_width-1];
assign Bit[1041] = V_1042[quan_width-1];
assign Bit[1042] = V_1043[quan_width-1];
assign Bit[1043] = V_1044[quan_width-1];
assign Bit[1044] = V_1045[quan_width-1];
assign Bit[1045] = V_1046[quan_width-1];
assign Bit[1046] = V_1047[quan_width-1];
assign Bit[1047] = V_1048[quan_width-1];
assign Bit[1048] = V_1049[quan_width-1];
assign Bit[1049] = V_1050[quan_width-1];
assign Bit[1050] = V_1051[quan_width-1];
assign Bit[1051] = V_1052[quan_width-1];
assign Bit[1052] = V_1053[quan_width-1];
assign Bit[1053] = V_1054[quan_width-1];
assign Bit[1054] = V_1055[quan_width-1];
assign Bit[1055] = V_1056[quan_width-1];
assign Bit[1056] = V_1057[quan_width-1];
assign Bit[1057] = V_1058[quan_width-1];
assign Bit[1058] = V_1059[quan_width-1];
assign Bit[1059] = V_1060[quan_width-1];
assign Bit[1060] = V_1061[quan_width-1];
assign Bit[1061] = V_1062[quan_width-1];
assign Bit[1062] = V_1063[quan_width-1];
assign Bit[1063] = V_1064[quan_width-1];
assign Bit[1064] = V_1065[quan_width-1];
assign Bit[1065] = V_1066[quan_width-1];
assign Bit[1066] = V_1067[quan_width-1];
assign Bit[1067] = V_1068[quan_width-1];
assign Bit[1068] = V_1069[quan_width-1];
assign Bit[1069] = V_1070[quan_width-1];
assign Bit[1070] = V_1071[quan_width-1];
assign Bit[1071] = V_1072[quan_width-1];
assign Bit[1072] = V_1073[quan_width-1];
assign Bit[1073] = V_1074[quan_width-1];
assign Bit[1074] = V_1075[quan_width-1];
assign Bit[1075] = V_1076[quan_width-1];
assign Bit[1076] = V_1077[quan_width-1];
assign Bit[1077] = V_1078[quan_width-1];
assign Bit[1078] = V_1079[quan_width-1];
assign Bit[1079] = V_1080[quan_width-1];
assign Bit[1080] = V_1081[quan_width-1];
assign Bit[1081] = V_1082[quan_width-1];
assign Bit[1082] = V_1083[quan_width-1];
assign Bit[1083] = V_1084[quan_width-1];
assign Bit[1084] = V_1085[quan_width-1];
assign Bit[1085] = V_1086[quan_width-1];
assign Bit[1086] = V_1087[quan_width-1];
assign Bit[1087] = V_1088[quan_width-1];
assign Bit[1088] = V_1089[quan_width-1];
assign Bit[1089] = V_1090[quan_width-1];
assign Bit[1090] = V_1091[quan_width-1];
assign Bit[1091] = V_1092[quan_width-1];
assign Bit[1092] = V_1093[quan_width-1];
assign Bit[1093] = V_1094[quan_width-1];
assign Bit[1094] = V_1095[quan_width-1];
assign Bit[1095] = V_1096[quan_width-1];
assign Bit[1096] = V_1097[quan_width-1];
assign Bit[1097] = V_1098[quan_width-1];
assign Bit[1098] = V_1099[quan_width-1];
assign Bit[1099] = V_1100[quan_width-1];
assign Bit[1100] = V_1101[quan_width-1];
assign Bit[1101] = V_1102[quan_width-1];
assign Bit[1102] = V_1103[quan_width-1];
assign Bit[1103] = V_1104[quan_width-1];
assign Bit[1104] = V_1105[quan_width-1];
assign Bit[1105] = V_1106[quan_width-1];
assign Bit[1106] = V_1107[quan_width-1];
assign Bit[1107] = V_1108[quan_width-1];
assign Bit[1108] = V_1109[quan_width-1];
assign Bit[1109] = V_1110[quan_width-1];
assign Bit[1110] = V_1111[quan_width-1];
assign Bit[1111] = V_1112[quan_width-1];
assign Bit[1112] = V_1113[quan_width-1];
assign Bit[1113] = V_1114[quan_width-1];
assign Bit[1114] = V_1115[quan_width-1];
assign Bit[1115] = V_1116[quan_width-1];
assign Bit[1116] = V_1117[quan_width-1];
assign Bit[1117] = V_1118[quan_width-1];
assign Bit[1118] = V_1119[quan_width-1];
assign Bit[1119] = V_1120[quan_width-1];
assign Bit[1120] = V_1121[quan_width-1];
assign Bit[1121] = V_1122[quan_width-1];
assign Bit[1122] = V_1123[quan_width-1];
assign Bit[1123] = V_1124[quan_width-1];
assign Bit[1124] = V_1125[quan_width-1];
assign Bit[1125] = V_1126[quan_width-1];
assign Bit[1126] = V_1127[quan_width-1];
assign Bit[1127] = V_1128[quan_width-1];
assign Bit[1128] = V_1129[quan_width-1];
assign Bit[1129] = V_1130[quan_width-1];
assign Bit[1130] = V_1131[quan_width-1];
assign Bit[1131] = V_1132[quan_width-1];
assign Bit[1132] = V_1133[quan_width-1];
assign Bit[1133] = V_1134[quan_width-1];
assign Bit[1134] = V_1135[quan_width-1];
assign Bit[1135] = V_1136[quan_width-1];
assign Bit[1136] = V_1137[quan_width-1];
assign Bit[1137] = V_1138[quan_width-1];
assign Bit[1138] = V_1139[quan_width-1];
assign Bit[1139] = V_1140[quan_width-1];
assign Bit[1140] = V_1141[quan_width-1];
assign Bit[1141] = V_1142[quan_width-1];
assign Bit[1142] = V_1143[quan_width-1];
assign Bit[1143] = V_1144[quan_width-1];
assign Bit[1144] = V_1145[quan_width-1];
assign Bit[1145] = V_1146[quan_width-1];
assign Bit[1146] = V_1147[quan_width-1];
assign Bit[1147] = V_1148[quan_width-1];
assign Bit[1148] = V_1149[quan_width-1];
assign Bit[1149] = V_1150[quan_width-1];
assign Bit[1150] = V_1151[quan_width-1];
assign Bit[1151] = V_1152[quan_width-1];
assign Bit[1152] = V_1153[quan_width-1];
assign Bit[1153] = V_1154[quan_width-1];
assign Bit[1154] = V_1155[quan_width-1];
assign Bit[1155] = V_1156[quan_width-1];
assign Bit[1156] = V_1157[quan_width-1];
assign Bit[1157] = V_1158[quan_width-1];
assign Bit[1158] = V_1159[quan_width-1];
assign Bit[1159] = V_1160[quan_width-1];
assign Bit[1160] = V_1161[quan_width-1];
assign Bit[1161] = V_1162[quan_width-1];
assign Bit[1162] = V_1163[quan_width-1];
assign Bit[1163] = V_1164[quan_width-1];
assign Bit[1164] = V_1165[quan_width-1];
assign Bit[1165] = V_1166[quan_width-1];
assign Bit[1166] = V_1167[quan_width-1];
assign Bit[1167] = V_1168[quan_width-1];
assign Bit[1168] = V_1169[quan_width-1];
assign Bit[1169] = V_1170[quan_width-1];
assign Bit[1170] = V_1171[quan_width-1];
assign Bit[1171] = V_1172[quan_width-1];
assign Bit[1172] = V_1173[quan_width-1];
assign Bit[1173] = V_1174[quan_width-1];
assign Bit[1174] = V_1175[quan_width-1];
assign Bit[1175] = V_1176[quan_width-1];
assign Bit[1176] = V_1177[quan_width-1];
assign Bit[1177] = V_1178[quan_width-1];
assign Bit[1178] = V_1179[quan_width-1];
assign Bit[1179] = V_1180[quan_width-1];
assign Bit[1180] = V_1181[quan_width-1];
assign Bit[1181] = V_1182[quan_width-1];
assign Bit[1182] = V_1183[quan_width-1];
assign Bit[1183] = V_1184[quan_width-1];
assign Bit[1184] = V_1185[quan_width-1];
assign Bit[1185] = V_1186[quan_width-1];
assign Bit[1186] = V_1187[quan_width-1];
assign Bit[1187] = V_1188[quan_width-1];
assign Bit[1188] = V_1189[quan_width-1];
assign Bit[1189] = V_1190[quan_width-1];
assign Bit[1190] = V_1191[quan_width-1];
assign Bit[1191] = V_1192[quan_width-1];
assign Bit[1192] = V_1193[quan_width-1];
assign Bit[1193] = V_1194[quan_width-1];
assign Bit[1194] = V_1195[quan_width-1];
assign Bit[1195] = V_1196[quan_width-1];
assign Bit[1196] = V_1197[quan_width-1];
assign Bit[1197] = V_1198[quan_width-1];
assign Bit[1198] = V_1199[quan_width-1];
assign Bit[1199] = V_1200[quan_width-1];
assign Bit[1200] = V_1201[quan_width-1];
assign Bit[1201] = V_1202[quan_width-1];
assign Bit[1202] = V_1203[quan_width-1];
assign Bit[1203] = V_1204[quan_width-1];
assign Bit[1204] = V_1205[quan_width-1];
assign Bit[1205] = V_1206[quan_width-1];
assign Bit[1206] = V_1207[quan_width-1];
assign Bit[1207] = V_1208[quan_width-1];
assign Bit[1208] = V_1209[quan_width-1];
assign Bit[1209] = V_1210[quan_width-1];
assign Bit[1210] = V_1211[quan_width-1];
assign Bit[1211] = V_1212[quan_width-1];
assign Bit[1212] = V_1213[quan_width-1];
assign Bit[1213] = V_1214[quan_width-1];
assign Bit[1214] = V_1215[quan_width-1];
assign Bit[1215] = V_1216[quan_width-1];
assign Bit[1216] = V_1217[quan_width-1];
assign Bit[1217] = V_1218[quan_width-1];
assign Bit[1218] = V_1219[quan_width-1];
assign Bit[1219] = V_1220[quan_width-1];
assign Bit[1220] = V_1221[quan_width-1];
assign Bit[1221] = V_1222[quan_width-1];
assign Bit[1222] = V_1223[quan_width-1];
assign Bit[1223] = V_1224[quan_width-1];
assign Bit[1224] = V_1225[quan_width-1];
assign Bit[1225] = V_1226[quan_width-1];
assign Bit[1226] = V_1227[quan_width-1];
assign Bit[1227] = V_1228[quan_width-1];
assign Bit[1228] = V_1229[quan_width-1];
assign Bit[1229] = V_1230[quan_width-1];
assign Bit[1230] = V_1231[quan_width-1];
assign Bit[1231] = V_1232[quan_width-1];
assign Bit[1232] = V_1233[quan_width-1];
assign Bit[1233] = V_1234[quan_width-1];
assign Bit[1234] = V_1235[quan_width-1];
assign Bit[1235] = V_1236[quan_width-1];
assign Bit[1236] = V_1237[quan_width-1];
assign Bit[1237] = V_1238[quan_width-1];
assign Bit[1238] = V_1239[quan_width-1];
assign Bit[1239] = V_1240[quan_width-1];
assign Bit[1240] = V_1241[quan_width-1];
assign Bit[1241] = V_1242[quan_width-1];
assign Bit[1242] = V_1243[quan_width-1];
assign Bit[1243] = V_1244[quan_width-1];
assign Bit[1244] = V_1245[quan_width-1];
assign Bit[1245] = V_1246[quan_width-1];
assign Bit[1246] = V_1247[quan_width-1];
assign Bit[1247] = V_1248[quan_width-1];
assign Bit[1248] = V_1249[quan_width-1];
assign Bit[1249] = V_1250[quan_width-1];
assign Bit[1250] = V_1251[quan_width-1];
assign Bit[1251] = V_1252[quan_width-1];
assign Bit[1252] = V_1253[quan_width-1];
assign Bit[1253] = V_1254[quan_width-1];
assign Bit[1254] = V_1255[quan_width-1];
assign Bit[1255] = V_1256[quan_width-1];
assign Bit[1256] = V_1257[quan_width-1];
assign Bit[1257] = V_1258[quan_width-1];
assign Bit[1258] = V_1259[quan_width-1];
assign Bit[1259] = V_1260[quan_width-1];
assign Bit[1260] = V_1261[quan_width-1];
assign Bit[1261] = V_1262[quan_width-1];
assign Bit[1262] = V_1263[quan_width-1];
assign Bit[1263] = V_1264[quan_width-1];
assign Bit[1264] = V_1265[quan_width-1];
assign Bit[1265] = V_1266[quan_width-1];
assign Bit[1266] = V_1267[quan_width-1];
assign Bit[1267] = V_1268[quan_width-1];
assign Bit[1268] = V_1269[quan_width-1];
assign Bit[1269] = V_1270[quan_width-1];
assign Bit[1270] = V_1271[quan_width-1];
assign Bit[1271] = V_1272[quan_width-1];
assign Bit[1272] = V_1273[quan_width-1];
assign Bit[1273] = V_1274[quan_width-1];
assign Bit[1274] = V_1275[quan_width-1];
assign Bit[1275] = V_1276[quan_width-1];
assign Bit[1276] = V_1277[quan_width-1];
assign Bit[1277] = V_1278[quan_width-1];
assign Bit[1278] = V_1279[quan_width-1];
assign Bit[1279] = V_1280[quan_width-1];
assign Bit[1280] = V_1281[quan_width-1];
assign Bit[1281] = V_1282[quan_width-1];
assign Bit[1282] = V_1283[quan_width-1];
assign Bit[1283] = V_1284[quan_width-1];
assign Bit[1284] = V_1285[quan_width-1];
assign Bit[1285] = V_1286[quan_width-1];
assign Bit[1286] = V_1287[quan_width-1];
assign Bit[1287] = V_1288[quan_width-1];
assign Bit[1288] = V_1289[quan_width-1];
assign Bit[1289] = V_1290[quan_width-1];
assign Bit[1290] = V_1291[quan_width-1];
assign Bit[1291] = V_1292[quan_width-1];
assign Bit[1292] = V_1293[quan_width-1];
assign Bit[1293] = V_1294[quan_width-1];
assign Bit[1294] = V_1295[quan_width-1];
assign Bit[1295] = V_1296[quan_width-1];
assign Bit[1296] = V_1297[quan_width-1];
assign Bit[1297] = V_1298[quan_width-1];
assign Bit[1298] = V_1299[quan_width-1];
assign Bit[1299] = V_1300[quan_width-1];
assign Bit[1300] = V_1301[quan_width-1];
assign Bit[1301] = V_1302[quan_width-1];
assign Bit[1302] = V_1303[quan_width-1];
assign Bit[1303] = V_1304[quan_width-1];
assign Bit[1304] = V_1305[quan_width-1];
assign Bit[1305] = V_1306[quan_width-1];
assign Bit[1306] = V_1307[quan_width-1];
assign Bit[1307] = V_1308[quan_width-1];
assign Bit[1308] = V_1309[quan_width-1];
assign Bit[1309] = V_1310[quan_width-1];
assign Bit[1310] = V_1311[quan_width-1];
assign Bit[1311] = V_1312[quan_width-1];
assign Bit[1312] = V_1313[quan_width-1];
assign Bit[1313] = V_1314[quan_width-1];
assign Bit[1314] = V_1315[quan_width-1];
assign Bit[1315] = V_1316[quan_width-1];
assign Bit[1316] = V_1317[quan_width-1];
assign Bit[1317] = V_1318[quan_width-1];
assign Bit[1318] = V_1319[quan_width-1];
assign Bit[1319] = V_1320[quan_width-1];
assign Bit[1320] = V_1321[quan_width-1];
assign Bit[1321] = V_1322[quan_width-1];
assign Bit[1322] = V_1323[quan_width-1];
assign Bit[1323] = V_1324[quan_width-1];
assign Bit[1324] = V_1325[quan_width-1];
assign Bit[1325] = V_1326[quan_width-1];
assign Bit[1326] = V_1327[quan_width-1];
assign Bit[1327] = V_1328[quan_width-1];
assign Bit[1328] = V_1329[quan_width-1];
assign Bit[1329] = V_1330[quan_width-1];
assign Bit[1330] = V_1331[quan_width-1];
assign Bit[1331] = V_1332[quan_width-1];
assign Bit[1332] = V_1333[quan_width-1];
assign Bit[1333] = V_1334[quan_width-1];
assign Bit[1334] = V_1335[quan_width-1];
assign Bit[1335] = V_1336[quan_width-1];
assign Bit[1336] = V_1337[quan_width-1];
assign Bit[1337] = V_1338[quan_width-1];
assign Bit[1338] = V_1339[quan_width-1];
assign Bit[1339] = V_1340[quan_width-1];
assign Bit[1340] = V_1341[quan_width-1];
assign Bit[1341] = V_1342[quan_width-1];
assign Bit[1342] = V_1343[quan_width-1];
assign Bit[1343] = V_1344[quan_width-1];
assign Bit[1344] = V_1345[quan_width-1];
assign Bit[1345] = V_1346[quan_width-1];
assign Bit[1346] = V_1347[quan_width-1];
assign Bit[1347] = V_1348[quan_width-1];
assign Bit[1348] = V_1349[quan_width-1];
assign Bit[1349] = V_1350[quan_width-1];
assign Bit[1350] = V_1351[quan_width-1];
assign Bit[1351] = V_1352[quan_width-1];
assign Bit[1352] = V_1353[quan_width-1];
assign Bit[1353] = V_1354[quan_width-1];
assign Bit[1354] = V_1355[quan_width-1];
assign Bit[1355] = V_1356[quan_width-1];
assign Bit[1356] = V_1357[quan_width-1];
assign Bit[1357] = V_1358[quan_width-1];
assign Bit[1358] = V_1359[quan_width-1];
assign Bit[1359] = V_1360[quan_width-1];
assign Bit[1360] = V_1361[quan_width-1];
assign Bit[1361] = V_1362[quan_width-1];
assign Bit[1362] = V_1363[quan_width-1];
assign Bit[1363] = V_1364[quan_width-1];
assign Bit[1364] = V_1365[quan_width-1];
assign Bit[1365] = V_1366[quan_width-1];
assign Bit[1366] = V_1367[quan_width-1];
assign Bit[1367] = V_1368[quan_width-1];
assign Bit[1368] = V_1369[quan_width-1];
assign Bit[1369] = V_1370[quan_width-1];
assign Bit[1370] = V_1371[quan_width-1];
assign Bit[1371] = V_1372[quan_width-1];
assign Bit[1372] = V_1373[quan_width-1];
assign Bit[1373] = V_1374[quan_width-1];
assign Bit[1374] = V_1375[quan_width-1];
assign Bit[1375] = V_1376[quan_width-1];
assign Bit[1376] = V_1377[quan_width-1];
assign Bit[1377] = V_1378[quan_width-1];
assign Bit[1378] = V_1379[quan_width-1];
assign Bit[1379] = V_1380[quan_width-1];
assign Bit[1380] = V_1381[quan_width-1];
assign Bit[1381] = V_1382[quan_width-1];
assign Bit[1382] = V_1383[quan_width-1];
assign Bit[1383] = V_1384[quan_width-1];
assign Bit[1384] = V_1385[quan_width-1];
assign Bit[1385] = V_1386[quan_width-1];
assign Bit[1386] = V_1387[quan_width-1];
assign Bit[1387] = V_1388[quan_width-1];
assign Bit[1388] = V_1389[quan_width-1];
assign Bit[1389] = V_1390[quan_width-1];
assign Bit[1390] = V_1391[quan_width-1];
assign Bit[1391] = V_1392[quan_width-1];
assign Bit[1392] = V_1393[quan_width-1];
assign Bit[1393] = V_1394[quan_width-1];
assign Bit[1394] = V_1395[quan_width-1];
assign Bit[1395] = V_1396[quan_width-1];
assign Bit[1396] = V_1397[quan_width-1];
assign Bit[1397] = V_1398[quan_width-1];
assign Bit[1398] = V_1399[quan_width-1];
assign Bit[1399] = V_1400[quan_width-1];
assign Bit[1400] = V_1401[quan_width-1];
assign Bit[1401] = V_1402[quan_width-1];
assign Bit[1402] = V_1403[quan_width-1];
assign Bit[1403] = V_1404[quan_width-1];
assign Bit[1404] = V_1405[quan_width-1];
assign Bit[1405] = V_1406[quan_width-1];
assign Bit[1406] = V_1407[quan_width-1];
assign Bit[1407] = V_1408[quan_width-1];
assign Bit[1408] = V_1409[quan_width-1];
assign Bit[1409] = V_1410[quan_width-1];
assign Bit[1410] = V_1411[quan_width-1];
assign Bit[1411] = V_1412[quan_width-1];
assign Bit[1412] = V_1413[quan_width-1];
assign Bit[1413] = V_1414[quan_width-1];
assign Bit[1414] = V_1415[quan_width-1];
assign Bit[1415] = V_1416[quan_width-1];
assign Bit[1416] = V_1417[quan_width-1];
assign Bit[1417] = V_1418[quan_width-1];
assign Bit[1418] = V_1419[quan_width-1];
assign Bit[1419] = V_1420[quan_width-1];
assign Bit[1420] = V_1421[quan_width-1];
assign Bit[1421] = V_1422[quan_width-1];
assign Bit[1422] = V_1423[quan_width-1];
assign Bit[1423] = V_1424[quan_width-1];
assign Bit[1424] = V_1425[quan_width-1];
assign Bit[1425] = V_1426[quan_width-1];
assign Bit[1426] = V_1427[quan_width-1];
assign Bit[1427] = V_1428[quan_width-1];
assign Bit[1428] = V_1429[quan_width-1];
assign Bit[1429] = V_1430[quan_width-1];
assign Bit[1430] = V_1431[quan_width-1];
assign Bit[1431] = V_1432[quan_width-1];
assign Bit[1432] = V_1433[quan_width-1];
assign Bit[1433] = V_1434[quan_width-1];
assign Bit[1434] = V_1435[quan_width-1];
assign Bit[1435] = V_1436[quan_width-1];
assign Bit[1436] = V_1437[quan_width-1];
assign Bit[1437] = V_1438[quan_width-1];
assign Bit[1438] = V_1439[quan_width-1];
assign Bit[1439] = V_1440[quan_width-1];

CNU_19 #(quan_width) CNU1 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_5_1),
	.V2C_2 (V2C_89_1),
	.V2C_3 (V2C_109_1),
	.V2C_4 (V2C_170_1),
	.V2C_5 (V2C_232_1),
	.V2C_6 (V2C_275_1),
	.V2C_7 (V2C_375_1),
	.V2C_8 (V2C_429_1),
	.V2C_9 (V2C_526_1),
	.V2C_10 (V2C_762_1),
	.V2C_11 (V2C_810_1),
	.V2C_12 (V2C_858_1),
	.V2C_13 (V2C_899_1),
	.V2C_14 (V2C_940_1),
	.V2C_15 (V2C_974_1),
	.V2C_16 (V2C_1013_1),
	.V2C_17 (V2C_1087_1),
	.V2C_18 (V2C_1146_1),
	.V2C_19 (V2C_1153_1),
	.C2V_1 (C2V_1_5),
	.C2V_2 (C2V_1_89),
	.C2V_3 (C2V_1_109),
	.C2V_4 (C2V_1_170),
	.C2V_5 (C2V_1_232),
	.C2V_6 (C2V_1_275),
	.C2V_7 (C2V_1_375),
	.C2V_8 (C2V_1_429),
	.C2V_9 (C2V_1_526),
	.C2V_10 (C2V_1_762),
	.C2V_11 (C2V_1_810),
	.C2V_12 (C2V_1_858),
	.C2V_13 (C2V_1_899),
	.C2V_14 (C2V_1_940),
	.C2V_15 (C2V_1_974),
	.C2V_16 (C2V_1_1013),
	.C2V_17 (C2V_1_1087),
	.C2V_18 (C2V_1_1146),
	.C2V_19 (C2V_1_1153),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU2 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_14_2),
	.V2C_2 (V2C_63_2),
	.V2C_3 (V2C_119_2),
	.V2C_4 (V2C_167_2),
	.V2C_5 (V2C_196_2),
	.V2C_6 (V2C_265_2),
	.V2C_7 (V2C_316_2),
	.V2C_8 (V2C_423_2),
	.V2C_9 (V2C_512_2),
	.V2C_10 (V2C_672_2),
	.V2C_11 (V2C_685_2),
	.V2C_12 (V2C_853_2),
	.V2C_13 (V2C_895_2),
	.V2C_14 (V2C_958_2),
	.V2C_15 (V2C_989_2),
	.V2C_16 (V2C_1021_2),
	.V2C_17 (V2C_1088_2),
	.V2C_18 (V2C_1119_2),
	.V2C_19 (V2C_1153_2),
	.V2C_20 (V2C_1154_2),
	.C2V_1 (C2V_2_14),
	.C2V_2 (C2V_2_63),
	.C2V_3 (C2V_2_119),
	.C2V_4 (C2V_2_167),
	.C2V_5 (C2V_2_196),
	.C2V_6 (C2V_2_265),
	.C2V_7 (C2V_2_316),
	.C2V_8 (C2V_2_423),
	.C2V_9 (C2V_2_512),
	.C2V_10 (C2V_2_672),
	.C2V_11 (C2V_2_685),
	.C2V_12 (C2V_2_853),
	.C2V_13 (C2V_2_895),
	.C2V_14 (C2V_2_958),
	.C2V_15 (C2V_2_989),
	.C2V_16 (C2V_2_1021),
	.C2V_17 (C2V_2_1088),
	.C2V_18 (C2V_2_1119),
	.C2V_19 (C2V_2_1153),
	.C2V_20 (C2V_2_1154),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU3 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_9_3),
	.V2C_2 (V2C_84_3),
	.V2C_3 (V2C_101_3),
	.V2C_4 (V2C_183_3),
	.V2C_5 (V2C_201_3),
	.V2C_6 (V2C_268_3),
	.V2C_7 (V2C_365_3),
	.V2C_8 (V2C_420_3),
	.V2C_9 (V2C_531_3),
	.V2C_10 (V2C_588_3),
	.V2C_11 (V2C_664_3),
	.V2C_12 (V2C_768_3),
	.V2C_13 (V2C_899_3),
	.V2C_14 (V2C_943_3),
	.V2C_15 (V2C_968_3),
	.V2C_16 (V2C_1028_3),
	.V2C_17 (V2C_1058_3),
	.V2C_18 (V2C_1151_3),
	.V2C_19 (V2C_1154_3),
	.V2C_20 (V2C_1155_3),
	.C2V_1 (C2V_3_9),
	.C2V_2 (C2V_3_84),
	.C2V_3 (C2V_3_101),
	.C2V_4 (C2V_3_183),
	.C2V_5 (C2V_3_201),
	.C2V_6 (C2V_3_268),
	.C2V_7 (C2V_3_365),
	.C2V_8 (C2V_3_420),
	.C2V_9 (C2V_3_531),
	.C2V_10 (C2V_3_588),
	.C2V_11 (C2V_3_664),
	.C2V_12 (C2V_3_768),
	.C2V_13 (C2V_3_899),
	.C2V_14 (C2V_3_943),
	.C2V_15 (C2V_3_968),
	.C2V_16 (C2V_3_1028),
	.C2V_17 (C2V_3_1058),
	.C2V_18 (C2V_3_1151),
	.C2V_19 (C2V_3_1154),
	.C2V_20 (C2V_3_1155),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU4 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_28_4),
	.V2C_2 (V2C_87_4),
	.V2C_3 (V2C_126_4),
	.V2C_4 (V2C_182_4),
	.V2C_5 (V2C_199_4),
	.V2C_6 (V2C_253_4),
	.V2C_7 (V2C_477_4),
	.V2C_8 (V2C_517_4),
	.V2C_9 (V2C_553_4),
	.V2C_10 (V2C_615_4),
	.V2C_11 (V2C_640_4),
	.V2C_12 (V2C_686_4),
	.V2C_13 (V2C_903_4),
	.V2C_14 (V2C_927_4),
	.V2C_15 (V2C_963_4),
	.V2C_16 (V2C_1041_4),
	.V2C_17 (V2C_1068_4),
	.V2C_18 (V2C_1132_4),
	.V2C_19 (V2C_1155_4),
	.V2C_20 (V2C_1156_4),
	.C2V_1 (C2V_4_28),
	.C2V_2 (C2V_4_87),
	.C2V_3 (C2V_4_126),
	.C2V_4 (C2V_4_182),
	.C2V_5 (C2V_4_199),
	.C2V_6 (C2V_4_253),
	.C2V_7 (C2V_4_477),
	.C2V_8 (C2V_4_517),
	.C2V_9 (C2V_4_553),
	.C2V_10 (C2V_4_615),
	.C2V_11 (C2V_4_640),
	.C2V_12 (C2V_4_686),
	.C2V_13 (C2V_4_903),
	.C2V_14 (C2V_4_927),
	.C2V_15 (C2V_4_963),
	.C2V_16 (C2V_4_1041),
	.C2V_17 (C2V_4_1068),
	.C2V_18 (C2V_4_1132),
	.C2V_19 (C2V_4_1155),
	.C2V_20 (C2V_4_1156),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU5 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_47_5),
	.V2C_2 (V2C_57_5),
	.V2C_3 (V2C_140_5),
	.V2C_4 (V2C_163_5),
	.V2C_5 (V2C_227_5),
	.V2C_6 (V2C_245_5),
	.V2C_7 (V2C_294_5),
	.V2C_8 (V2C_361_5),
	.V2C_9 (V2C_440_5),
	.V2C_10 (V2C_674_5),
	.V2C_11 (V2C_738_5),
	.V2C_12 (V2C_792_5),
	.V2C_13 (V2C_870_5),
	.V2C_14 (V2C_918_5),
	.V2C_15 (V2C_961_5),
	.V2C_16 (V2C_1013_5),
	.V2C_17 (V2C_1062_5),
	.V2C_18 (V2C_1110_5),
	.V2C_19 (V2C_1156_5),
	.V2C_20 (V2C_1157_5),
	.C2V_1 (C2V_5_47),
	.C2V_2 (C2V_5_57),
	.C2V_3 (C2V_5_140),
	.C2V_4 (C2V_5_163),
	.C2V_5 (C2V_5_227),
	.C2V_6 (C2V_5_245),
	.C2V_7 (C2V_5_294),
	.C2V_8 (C2V_5_361),
	.C2V_9 (C2V_5_440),
	.C2V_10 (C2V_5_674),
	.C2V_11 (C2V_5_738),
	.C2V_12 (C2V_5_792),
	.C2V_13 (C2V_5_870),
	.C2V_14 (C2V_5_918),
	.C2V_15 (C2V_5_961),
	.C2V_16 (C2V_5_1013),
	.C2V_17 (C2V_5_1062),
	.C2V_18 (C2V_5_1110),
	.C2V_19 (C2V_5_1156),
	.C2V_20 (C2V_5_1157),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU6 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_30_6),
	.V2C_2 (V2C_54_6),
	.V2C_3 (V2C_142_6),
	.V2C_4 (V2C_162_6),
	.V2C_5 (V2C_196_6),
	.V2C_6 (V2C_275_6),
	.V2C_7 (V2C_328_6),
	.V2C_8 (V2C_480_6),
	.V2C_9 (V2C_529_6),
	.V2C_10 (V2C_610_6),
	.V2C_11 (V2C_814_6),
	.V2C_12 (V2C_842_6),
	.V2C_13 (V2C_875_6),
	.V2C_14 (V2C_937_6),
	.V2C_15 (V2C_972_6),
	.V2C_16 (V2C_1039_6),
	.V2C_17 (V2C_1103_6),
	.V2C_18 (V2C_1105_6),
	.V2C_19 (V2C_1157_6),
	.V2C_20 (V2C_1158_6),
	.C2V_1 (C2V_6_30),
	.C2V_2 (C2V_6_54),
	.C2V_3 (C2V_6_142),
	.C2V_4 (C2V_6_162),
	.C2V_5 (C2V_6_196),
	.C2V_6 (C2V_6_275),
	.C2V_7 (C2V_6_328),
	.C2V_8 (C2V_6_480),
	.C2V_9 (C2V_6_529),
	.C2V_10 (C2V_6_610),
	.C2V_11 (C2V_6_814),
	.C2V_12 (C2V_6_842),
	.C2V_13 (C2V_6_875),
	.C2V_14 (C2V_6_937),
	.C2V_15 (C2V_6_972),
	.C2V_16 (C2V_6_1039),
	.C2V_17 (C2V_6_1103),
	.C2V_18 (C2V_6_1105),
	.C2V_19 (C2V_6_1157),
	.C2V_20 (C2V_6_1158),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU7 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_6_7),
	.V2C_2 (V2C_90_7),
	.V2C_3 (V2C_110_7),
	.V2C_4 (V2C_171_7),
	.V2C_5 (V2C_233_7),
	.V2C_6 (V2C_276_7),
	.V2C_7 (V2C_376_7),
	.V2C_8 (V2C_430_7),
	.V2C_9 (V2C_527_7),
	.V2C_10 (V2C_763_7),
	.V2C_11 (V2C_811_7),
	.V2C_12 (V2C_859_7),
	.V2C_13 (V2C_900_7),
	.V2C_14 (V2C_941_7),
	.V2C_15 (V2C_975_7),
	.V2C_16 (V2C_1014_7),
	.V2C_17 (V2C_1088_7),
	.V2C_18 (V2C_1147_7),
	.V2C_19 (V2C_1158_7),
	.V2C_20 (V2C_1159_7),
	.C2V_1 (C2V_7_6),
	.C2V_2 (C2V_7_90),
	.C2V_3 (C2V_7_110),
	.C2V_4 (C2V_7_171),
	.C2V_5 (C2V_7_233),
	.C2V_6 (C2V_7_276),
	.C2V_7 (C2V_7_376),
	.C2V_8 (C2V_7_430),
	.C2V_9 (C2V_7_527),
	.C2V_10 (C2V_7_763),
	.C2V_11 (C2V_7_811),
	.C2V_12 (C2V_7_859),
	.C2V_13 (C2V_7_900),
	.C2V_14 (C2V_7_941),
	.C2V_15 (C2V_7_975),
	.C2V_16 (C2V_7_1014),
	.C2V_17 (C2V_7_1088),
	.C2V_18 (C2V_7_1147),
	.C2V_19 (C2V_7_1158),
	.C2V_20 (C2V_7_1159),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU8 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_15_8),
	.V2C_2 (V2C_64_8),
	.V2C_3 (V2C_120_8),
	.V2C_4 (V2C_168_8),
	.V2C_5 (V2C_197_8),
	.V2C_6 (V2C_266_8),
	.V2C_7 (V2C_317_8),
	.V2C_8 (V2C_424_8),
	.V2C_9 (V2C_513_8),
	.V2C_10 (V2C_625_8),
	.V2C_11 (V2C_686_8),
	.V2C_12 (V2C_854_8),
	.V2C_13 (V2C_896_8),
	.V2C_14 (V2C_959_8),
	.V2C_15 (V2C_990_8),
	.V2C_16 (V2C_1022_8),
	.V2C_17 (V2C_1089_8),
	.V2C_18 (V2C_1120_8),
	.V2C_19 (V2C_1159_8),
	.V2C_20 (V2C_1160_8),
	.C2V_1 (C2V_8_15),
	.C2V_2 (C2V_8_64),
	.C2V_3 (C2V_8_120),
	.C2V_4 (C2V_8_168),
	.C2V_5 (C2V_8_197),
	.C2V_6 (C2V_8_266),
	.C2V_7 (C2V_8_317),
	.C2V_8 (C2V_8_424),
	.C2V_9 (C2V_8_513),
	.C2V_10 (C2V_8_625),
	.C2V_11 (C2V_8_686),
	.C2V_12 (C2V_8_854),
	.C2V_13 (C2V_8_896),
	.C2V_14 (C2V_8_959),
	.C2V_15 (C2V_8_990),
	.C2V_16 (C2V_8_1022),
	.C2V_17 (C2V_8_1089),
	.C2V_18 (C2V_8_1120),
	.C2V_19 (C2V_8_1159),
	.C2V_20 (C2V_8_1160),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU9 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_10_9),
	.V2C_2 (V2C_85_9),
	.V2C_3 (V2C_102_9),
	.V2C_4 (V2C_184_9),
	.V2C_5 (V2C_202_9),
	.V2C_6 (V2C_269_9),
	.V2C_7 (V2C_366_9),
	.V2C_8 (V2C_421_9),
	.V2C_9 (V2C_532_9),
	.V2C_10 (V2C_589_9),
	.V2C_11 (V2C_665_9),
	.V2C_12 (V2C_721_9),
	.V2C_13 (V2C_900_9),
	.V2C_14 (V2C_944_9),
	.V2C_15 (V2C_969_9),
	.V2C_16 (V2C_1029_9),
	.V2C_17 (V2C_1059_9),
	.V2C_18 (V2C_1152_9),
	.V2C_19 (V2C_1160_9),
	.V2C_20 (V2C_1161_9),
	.C2V_1 (C2V_9_10),
	.C2V_2 (C2V_9_85),
	.C2V_3 (C2V_9_102),
	.C2V_4 (C2V_9_184),
	.C2V_5 (C2V_9_202),
	.C2V_6 (C2V_9_269),
	.C2V_7 (C2V_9_366),
	.C2V_8 (C2V_9_421),
	.C2V_9 (C2V_9_532),
	.C2V_10 (C2V_9_589),
	.C2V_11 (C2V_9_665),
	.C2V_12 (C2V_9_721),
	.C2V_13 (C2V_9_900),
	.C2V_14 (C2V_9_944),
	.C2V_15 (C2V_9_969),
	.C2V_16 (C2V_9_1029),
	.C2V_17 (C2V_9_1059),
	.C2V_18 (C2V_9_1152),
	.C2V_19 (C2V_9_1160),
	.C2V_20 (C2V_9_1161),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU10 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_29_10),
	.V2C_2 (V2C_88_10),
	.V2C_3 (V2C_127_10),
	.V2C_4 (V2C_183_10),
	.V2C_5 (V2C_200_10),
	.V2C_6 (V2C_254_10),
	.V2C_7 (V2C_478_10),
	.V2C_8 (V2C_518_10),
	.V2C_9 (V2C_554_10),
	.V2C_10 (V2C_616_10),
	.V2C_11 (V2C_641_10),
	.V2C_12 (V2C_687_10),
	.V2C_13 (V2C_904_10),
	.V2C_14 (V2C_928_10),
	.V2C_15 (V2C_964_10),
	.V2C_16 (V2C_1042_10),
	.V2C_17 (V2C_1069_10),
	.V2C_18 (V2C_1133_10),
	.V2C_19 (V2C_1161_10),
	.V2C_20 (V2C_1162_10),
	.C2V_1 (C2V_10_29),
	.C2V_2 (C2V_10_88),
	.C2V_3 (C2V_10_127),
	.C2V_4 (C2V_10_183),
	.C2V_5 (C2V_10_200),
	.C2V_6 (C2V_10_254),
	.C2V_7 (C2V_10_478),
	.C2V_8 (C2V_10_518),
	.C2V_9 (C2V_10_554),
	.C2V_10 (C2V_10_616),
	.C2V_11 (C2V_10_641),
	.C2V_12 (C2V_10_687),
	.C2V_13 (C2V_10_904),
	.C2V_14 (C2V_10_928),
	.C2V_15 (C2V_10_964),
	.C2V_16 (C2V_10_1042),
	.C2V_17 (C2V_10_1069),
	.C2V_18 (C2V_10_1133),
	.C2V_19 (C2V_10_1161),
	.C2V_20 (C2V_10_1162),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU11 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_48_11),
	.V2C_2 (V2C_58_11),
	.V2C_3 (V2C_141_11),
	.V2C_4 (V2C_164_11),
	.V2C_5 (V2C_228_11),
	.V2C_6 (V2C_246_11),
	.V2C_7 (V2C_295_11),
	.V2C_8 (V2C_362_11),
	.V2C_9 (V2C_441_11),
	.V2C_10 (V2C_675_11),
	.V2C_11 (V2C_739_11),
	.V2C_12 (V2C_793_11),
	.V2C_13 (V2C_871_11),
	.V2C_14 (V2C_919_11),
	.V2C_15 (V2C_962_11),
	.V2C_16 (V2C_1014_11),
	.V2C_17 (V2C_1063_11),
	.V2C_18 (V2C_1111_11),
	.V2C_19 (V2C_1162_11),
	.V2C_20 (V2C_1163_11),
	.C2V_1 (C2V_11_48),
	.C2V_2 (C2V_11_58),
	.C2V_3 (C2V_11_141),
	.C2V_4 (C2V_11_164),
	.C2V_5 (C2V_11_228),
	.C2V_6 (C2V_11_246),
	.C2V_7 (C2V_11_295),
	.C2V_8 (C2V_11_362),
	.C2V_9 (C2V_11_441),
	.C2V_10 (C2V_11_675),
	.C2V_11 (C2V_11_739),
	.C2V_12 (C2V_11_793),
	.C2V_13 (C2V_11_871),
	.C2V_14 (C2V_11_919),
	.C2V_15 (C2V_11_962),
	.C2V_16 (C2V_11_1014),
	.C2V_17 (C2V_11_1063),
	.C2V_18 (C2V_11_1111),
	.C2V_19 (C2V_11_1162),
	.C2V_20 (C2V_11_1163),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU12 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_31_12),
	.V2C_2 (V2C_55_12),
	.V2C_3 (V2C_143_12),
	.V2C_4 (V2C_163_12),
	.V2C_5 (V2C_197_12),
	.V2C_6 (V2C_276_12),
	.V2C_7 (V2C_329_12),
	.V2C_8 (V2C_433_12),
	.V2C_9 (V2C_530_12),
	.V2C_10 (V2C_611_12),
	.V2C_11 (V2C_815_12),
	.V2C_12 (V2C_843_12),
	.V2C_13 (V2C_876_12),
	.V2C_14 (V2C_938_12),
	.V2C_15 (V2C_973_12),
	.V2C_16 (V2C_1040_12),
	.V2C_17 (V2C_1104_12),
	.V2C_18 (V2C_1106_12),
	.V2C_19 (V2C_1163_12),
	.V2C_20 (V2C_1164_12),
	.C2V_1 (C2V_12_31),
	.C2V_2 (C2V_12_55),
	.C2V_3 (C2V_12_143),
	.C2V_4 (C2V_12_163),
	.C2V_5 (C2V_12_197),
	.C2V_6 (C2V_12_276),
	.C2V_7 (C2V_12_329),
	.C2V_8 (C2V_12_433),
	.C2V_9 (C2V_12_530),
	.C2V_10 (C2V_12_611),
	.C2V_11 (C2V_12_815),
	.C2V_12 (C2V_12_843),
	.C2V_13 (C2V_12_876),
	.C2V_14 (C2V_12_938),
	.C2V_15 (C2V_12_973),
	.C2V_16 (C2V_12_1040),
	.C2V_17 (C2V_12_1104),
	.C2V_18 (C2V_12_1106),
	.C2V_19 (C2V_12_1163),
	.C2V_20 (C2V_12_1164),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU13 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_7_13),
	.V2C_2 (V2C_91_13),
	.V2C_3 (V2C_111_13),
	.V2C_4 (V2C_172_13),
	.V2C_5 (V2C_234_13),
	.V2C_6 (V2C_277_13),
	.V2C_7 (V2C_377_13),
	.V2C_8 (V2C_431_13),
	.V2C_9 (V2C_528_13),
	.V2C_10 (V2C_764_13),
	.V2C_11 (V2C_812_13),
	.V2C_12 (V2C_860_13),
	.V2C_13 (V2C_901_13),
	.V2C_14 (V2C_942_13),
	.V2C_15 (V2C_976_13),
	.V2C_16 (V2C_1015_13),
	.V2C_17 (V2C_1089_13),
	.V2C_18 (V2C_1148_13),
	.V2C_19 (V2C_1164_13),
	.V2C_20 (V2C_1165_13),
	.C2V_1 (C2V_13_7),
	.C2V_2 (C2V_13_91),
	.C2V_3 (C2V_13_111),
	.C2V_4 (C2V_13_172),
	.C2V_5 (C2V_13_234),
	.C2V_6 (C2V_13_277),
	.C2V_7 (C2V_13_377),
	.C2V_8 (C2V_13_431),
	.C2V_9 (C2V_13_528),
	.C2V_10 (C2V_13_764),
	.C2V_11 (C2V_13_812),
	.C2V_12 (C2V_13_860),
	.C2V_13 (C2V_13_901),
	.C2V_14 (C2V_13_942),
	.C2V_15 (C2V_13_976),
	.C2V_16 (C2V_13_1015),
	.C2V_17 (C2V_13_1089),
	.C2V_18 (C2V_13_1148),
	.C2V_19 (C2V_13_1164),
	.C2V_20 (C2V_13_1165),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU14 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_16_14),
	.V2C_2 (V2C_65_14),
	.V2C_3 (V2C_121_14),
	.V2C_4 (V2C_169_14),
	.V2C_5 (V2C_198_14),
	.V2C_6 (V2C_267_14),
	.V2C_7 (V2C_318_14),
	.V2C_8 (V2C_425_14),
	.V2C_9 (V2C_514_14),
	.V2C_10 (V2C_626_14),
	.V2C_11 (V2C_687_14),
	.V2C_12 (V2C_855_14),
	.V2C_13 (V2C_897_14),
	.V2C_14 (V2C_960_14),
	.V2C_15 (V2C_991_14),
	.V2C_16 (V2C_1023_14),
	.V2C_17 (V2C_1090_14),
	.V2C_18 (V2C_1121_14),
	.V2C_19 (V2C_1165_14),
	.V2C_20 (V2C_1166_14),
	.C2V_1 (C2V_14_16),
	.C2V_2 (C2V_14_65),
	.C2V_3 (C2V_14_121),
	.C2V_4 (C2V_14_169),
	.C2V_5 (C2V_14_198),
	.C2V_6 (C2V_14_267),
	.C2V_7 (C2V_14_318),
	.C2V_8 (C2V_14_425),
	.C2V_9 (C2V_14_514),
	.C2V_10 (C2V_14_626),
	.C2V_11 (C2V_14_687),
	.C2V_12 (C2V_14_855),
	.C2V_13 (C2V_14_897),
	.C2V_14 (C2V_14_960),
	.C2V_15 (C2V_14_991),
	.C2V_16 (C2V_14_1023),
	.C2V_17 (C2V_14_1090),
	.C2V_18 (C2V_14_1121),
	.C2V_19 (C2V_14_1165),
	.C2V_20 (C2V_14_1166),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU15 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_11_15),
	.V2C_2 (V2C_86_15),
	.V2C_3 (V2C_103_15),
	.V2C_4 (V2C_185_15),
	.V2C_5 (V2C_203_15),
	.V2C_6 (V2C_270_15),
	.V2C_7 (V2C_367_15),
	.V2C_8 (V2C_422_15),
	.V2C_9 (V2C_533_15),
	.V2C_10 (V2C_590_15),
	.V2C_11 (V2C_666_15),
	.V2C_12 (V2C_722_15),
	.V2C_13 (V2C_901_15),
	.V2C_14 (V2C_945_15),
	.V2C_15 (V2C_970_15),
	.V2C_16 (V2C_1030_15),
	.V2C_17 (V2C_1060_15),
	.V2C_18 (V2C_1105_15),
	.V2C_19 (V2C_1166_15),
	.V2C_20 (V2C_1167_15),
	.C2V_1 (C2V_15_11),
	.C2V_2 (C2V_15_86),
	.C2V_3 (C2V_15_103),
	.C2V_4 (C2V_15_185),
	.C2V_5 (C2V_15_203),
	.C2V_6 (C2V_15_270),
	.C2V_7 (C2V_15_367),
	.C2V_8 (C2V_15_422),
	.C2V_9 (C2V_15_533),
	.C2V_10 (C2V_15_590),
	.C2V_11 (C2V_15_666),
	.C2V_12 (C2V_15_722),
	.C2V_13 (C2V_15_901),
	.C2V_14 (C2V_15_945),
	.C2V_15 (C2V_15_970),
	.C2V_16 (C2V_15_1030),
	.C2V_17 (C2V_15_1060),
	.C2V_18 (C2V_15_1105),
	.C2V_19 (C2V_15_1166),
	.C2V_20 (C2V_15_1167),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU16 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_30_16),
	.V2C_2 (V2C_89_16),
	.V2C_3 (V2C_128_16),
	.V2C_4 (V2C_184_16),
	.V2C_5 (V2C_201_16),
	.V2C_6 (V2C_255_16),
	.V2C_7 (V2C_479_16),
	.V2C_8 (V2C_519_16),
	.V2C_9 (V2C_555_16),
	.V2C_10 (V2C_617_16),
	.V2C_11 (V2C_642_16),
	.V2C_12 (V2C_688_16),
	.V2C_13 (V2C_905_16),
	.V2C_14 (V2C_929_16),
	.V2C_15 (V2C_965_16),
	.V2C_16 (V2C_1043_16),
	.V2C_17 (V2C_1070_16),
	.V2C_18 (V2C_1134_16),
	.V2C_19 (V2C_1167_16),
	.V2C_20 (V2C_1168_16),
	.C2V_1 (C2V_16_30),
	.C2V_2 (C2V_16_89),
	.C2V_3 (C2V_16_128),
	.C2V_4 (C2V_16_184),
	.C2V_5 (C2V_16_201),
	.C2V_6 (C2V_16_255),
	.C2V_7 (C2V_16_479),
	.C2V_8 (C2V_16_519),
	.C2V_9 (C2V_16_555),
	.C2V_10 (C2V_16_617),
	.C2V_11 (C2V_16_642),
	.C2V_12 (C2V_16_688),
	.C2V_13 (C2V_16_905),
	.C2V_14 (C2V_16_929),
	.C2V_15 (C2V_16_965),
	.C2V_16 (C2V_16_1043),
	.C2V_17 (C2V_16_1070),
	.C2V_18 (C2V_16_1134),
	.C2V_19 (C2V_16_1167),
	.C2V_20 (C2V_16_1168),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU17 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_1_17),
	.V2C_2 (V2C_59_17),
	.V2C_3 (V2C_142_17),
	.V2C_4 (V2C_165_17),
	.V2C_5 (V2C_229_17),
	.V2C_6 (V2C_247_17),
	.V2C_7 (V2C_296_17),
	.V2C_8 (V2C_363_17),
	.V2C_9 (V2C_442_17),
	.V2C_10 (V2C_676_17),
	.V2C_11 (V2C_740_17),
	.V2C_12 (V2C_794_17),
	.V2C_13 (V2C_872_17),
	.V2C_14 (V2C_920_17),
	.V2C_15 (V2C_963_17),
	.V2C_16 (V2C_1015_17),
	.V2C_17 (V2C_1064_17),
	.V2C_18 (V2C_1112_17),
	.V2C_19 (V2C_1168_17),
	.V2C_20 (V2C_1169_17),
	.C2V_1 (C2V_17_1),
	.C2V_2 (C2V_17_59),
	.C2V_3 (C2V_17_142),
	.C2V_4 (C2V_17_165),
	.C2V_5 (C2V_17_229),
	.C2V_6 (C2V_17_247),
	.C2V_7 (C2V_17_296),
	.C2V_8 (C2V_17_363),
	.C2V_9 (C2V_17_442),
	.C2V_10 (C2V_17_676),
	.C2V_11 (C2V_17_740),
	.C2V_12 (C2V_17_794),
	.C2V_13 (C2V_17_872),
	.C2V_14 (C2V_17_920),
	.C2V_15 (C2V_17_963),
	.C2V_16 (C2V_17_1015),
	.C2V_17 (C2V_17_1064),
	.C2V_18 (C2V_17_1112),
	.C2V_19 (C2V_17_1168),
	.C2V_20 (C2V_17_1169),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU18 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_32_18),
	.V2C_2 (V2C_56_18),
	.V2C_3 (V2C_144_18),
	.V2C_4 (V2C_164_18),
	.V2C_5 (V2C_198_18),
	.V2C_6 (V2C_277_18),
	.V2C_7 (V2C_330_18),
	.V2C_8 (V2C_434_18),
	.V2C_9 (V2C_531_18),
	.V2C_10 (V2C_612_18),
	.V2C_11 (V2C_816_18),
	.V2C_12 (V2C_844_18),
	.V2C_13 (V2C_877_18),
	.V2C_14 (V2C_939_18),
	.V2C_15 (V2C_974_18),
	.V2C_16 (V2C_1041_18),
	.V2C_17 (V2C_1057_18),
	.V2C_18 (V2C_1107_18),
	.V2C_19 (V2C_1169_18),
	.V2C_20 (V2C_1170_18),
	.C2V_1 (C2V_18_32),
	.C2V_2 (C2V_18_56),
	.C2V_3 (C2V_18_144),
	.C2V_4 (C2V_18_164),
	.C2V_5 (C2V_18_198),
	.C2V_6 (C2V_18_277),
	.C2V_7 (C2V_18_330),
	.C2V_8 (C2V_18_434),
	.C2V_9 (C2V_18_531),
	.C2V_10 (C2V_18_612),
	.C2V_11 (C2V_18_816),
	.C2V_12 (C2V_18_844),
	.C2V_13 (C2V_18_877),
	.C2V_14 (C2V_18_939),
	.C2V_15 (C2V_18_974),
	.C2V_16 (C2V_18_1041),
	.C2V_17 (C2V_18_1057),
	.C2V_18 (C2V_18_1107),
	.C2V_19 (C2V_18_1169),
	.C2V_20 (C2V_18_1170),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU19 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_8_19),
	.V2C_2 (V2C_92_19),
	.V2C_3 (V2C_112_19),
	.V2C_4 (V2C_173_19),
	.V2C_5 (V2C_235_19),
	.V2C_6 (V2C_278_19),
	.V2C_7 (V2C_378_19),
	.V2C_8 (V2C_432_19),
	.V2C_9 (V2C_481_19),
	.V2C_10 (V2C_765_19),
	.V2C_11 (V2C_813_19),
	.V2C_12 (V2C_861_19),
	.V2C_13 (V2C_902_19),
	.V2C_14 (V2C_943_19),
	.V2C_15 (V2C_977_19),
	.V2C_16 (V2C_1016_19),
	.V2C_17 (V2C_1090_19),
	.V2C_18 (V2C_1149_19),
	.V2C_19 (V2C_1170_19),
	.V2C_20 (V2C_1171_19),
	.C2V_1 (C2V_19_8),
	.C2V_2 (C2V_19_92),
	.C2V_3 (C2V_19_112),
	.C2V_4 (C2V_19_173),
	.C2V_5 (C2V_19_235),
	.C2V_6 (C2V_19_278),
	.C2V_7 (C2V_19_378),
	.C2V_8 (C2V_19_432),
	.C2V_9 (C2V_19_481),
	.C2V_10 (C2V_19_765),
	.C2V_11 (C2V_19_813),
	.C2V_12 (C2V_19_861),
	.C2V_13 (C2V_19_902),
	.C2V_14 (C2V_19_943),
	.C2V_15 (C2V_19_977),
	.C2V_16 (C2V_19_1016),
	.C2V_17 (C2V_19_1090),
	.C2V_18 (C2V_19_1149),
	.C2V_19 (C2V_19_1170),
	.C2V_20 (C2V_19_1171),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU20 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_17_20),
	.V2C_2 (V2C_66_20),
	.V2C_3 (V2C_122_20),
	.V2C_4 (V2C_170_20),
	.V2C_5 (V2C_199_20),
	.V2C_6 (V2C_268_20),
	.V2C_7 (V2C_319_20),
	.V2C_8 (V2C_426_20),
	.V2C_9 (V2C_515_20),
	.V2C_10 (V2C_627_20),
	.V2C_11 (V2C_688_20),
	.V2C_12 (V2C_856_20),
	.V2C_13 (V2C_898_20),
	.V2C_14 (V2C_913_20),
	.V2C_15 (V2C_992_20),
	.V2C_16 (V2C_1024_20),
	.V2C_17 (V2C_1091_20),
	.V2C_18 (V2C_1122_20),
	.V2C_19 (V2C_1171_20),
	.V2C_20 (V2C_1172_20),
	.C2V_1 (C2V_20_17),
	.C2V_2 (C2V_20_66),
	.C2V_3 (C2V_20_122),
	.C2V_4 (C2V_20_170),
	.C2V_5 (C2V_20_199),
	.C2V_6 (C2V_20_268),
	.C2V_7 (C2V_20_319),
	.C2V_8 (C2V_20_426),
	.C2V_9 (C2V_20_515),
	.C2V_10 (C2V_20_627),
	.C2V_11 (C2V_20_688),
	.C2V_12 (C2V_20_856),
	.C2V_13 (C2V_20_898),
	.C2V_14 (C2V_20_913),
	.C2V_15 (C2V_20_992),
	.C2V_16 (C2V_20_1024),
	.C2V_17 (C2V_20_1091),
	.C2V_18 (C2V_20_1122),
	.C2V_19 (C2V_20_1171),
	.C2V_20 (C2V_20_1172),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU21 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_12_21),
	.V2C_2 (V2C_87_21),
	.V2C_3 (V2C_104_21),
	.V2C_4 (V2C_186_21),
	.V2C_5 (V2C_204_21),
	.V2C_6 (V2C_271_21),
	.V2C_7 (V2C_368_21),
	.V2C_8 (V2C_423_21),
	.V2C_9 (V2C_534_21),
	.V2C_10 (V2C_591_21),
	.V2C_11 (V2C_667_21),
	.V2C_12 (V2C_723_21),
	.V2C_13 (V2C_902_21),
	.V2C_14 (V2C_946_21),
	.V2C_15 (V2C_971_21),
	.V2C_16 (V2C_1031_21),
	.V2C_17 (V2C_1061_21),
	.V2C_18 (V2C_1106_21),
	.V2C_19 (V2C_1172_21),
	.V2C_20 (V2C_1173_21),
	.C2V_1 (C2V_21_12),
	.C2V_2 (C2V_21_87),
	.C2V_3 (C2V_21_104),
	.C2V_4 (C2V_21_186),
	.C2V_5 (C2V_21_204),
	.C2V_6 (C2V_21_271),
	.C2V_7 (C2V_21_368),
	.C2V_8 (C2V_21_423),
	.C2V_9 (C2V_21_534),
	.C2V_10 (C2V_21_591),
	.C2V_11 (C2V_21_667),
	.C2V_12 (C2V_21_723),
	.C2V_13 (C2V_21_902),
	.C2V_14 (C2V_21_946),
	.C2V_15 (C2V_21_971),
	.C2V_16 (C2V_21_1031),
	.C2V_17 (C2V_21_1061),
	.C2V_18 (C2V_21_1106),
	.C2V_19 (C2V_21_1172),
	.C2V_20 (C2V_21_1173),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU22 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_31_22),
	.V2C_2 (V2C_90_22),
	.V2C_3 (V2C_129_22),
	.V2C_4 (V2C_185_22),
	.V2C_5 (V2C_202_22),
	.V2C_6 (V2C_256_22),
	.V2C_7 (V2C_480_22),
	.V2C_8 (V2C_520_22),
	.V2C_9 (V2C_556_22),
	.V2C_10 (V2C_618_22),
	.V2C_11 (V2C_643_22),
	.V2C_12 (V2C_689_22),
	.V2C_13 (V2C_906_22),
	.V2C_14 (V2C_930_22),
	.V2C_15 (V2C_966_22),
	.V2C_16 (V2C_1044_22),
	.V2C_17 (V2C_1071_22),
	.V2C_18 (V2C_1135_22),
	.V2C_19 (V2C_1173_22),
	.V2C_20 (V2C_1174_22),
	.C2V_1 (C2V_22_31),
	.C2V_2 (C2V_22_90),
	.C2V_3 (C2V_22_129),
	.C2V_4 (C2V_22_185),
	.C2V_5 (C2V_22_202),
	.C2V_6 (C2V_22_256),
	.C2V_7 (C2V_22_480),
	.C2V_8 (C2V_22_520),
	.C2V_9 (C2V_22_556),
	.C2V_10 (C2V_22_618),
	.C2V_11 (C2V_22_643),
	.C2V_12 (C2V_22_689),
	.C2V_13 (C2V_22_906),
	.C2V_14 (C2V_22_930),
	.C2V_15 (C2V_22_966),
	.C2V_16 (C2V_22_1044),
	.C2V_17 (C2V_22_1071),
	.C2V_18 (C2V_22_1135),
	.C2V_19 (C2V_22_1173),
	.C2V_20 (C2V_22_1174),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU23 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_2_23),
	.V2C_2 (V2C_60_23),
	.V2C_3 (V2C_143_23),
	.V2C_4 (V2C_166_23),
	.V2C_5 (V2C_230_23),
	.V2C_6 (V2C_248_23),
	.V2C_7 (V2C_297_23),
	.V2C_8 (V2C_364_23),
	.V2C_9 (V2C_443_23),
	.V2C_10 (V2C_677_23),
	.V2C_11 (V2C_741_23),
	.V2C_12 (V2C_795_23),
	.V2C_13 (V2C_873_23),
	.V2C_14 (V2C_921_23),
	.V2C_15 (V2C_964_23),
	.V2C_16 (V2C_1016_23),
	.V2C_17 (V2C_1065_23),
	.V2C_18 (V2C_1113_23),
	.V2C_19 (V2C_1174_23),
	.V2C_20 (V2C_1175_23),
	.C2V_1 (C2V_23_2),
	.C2V_2 (C2V_23_60),
	.C2V_3 (C2V_23_143),
	.C2V_4 (C2V_23_166),
	.C2V_5 (C2V_23_230),
	.C2V_6 (C2V_23_248),
	.C2V_7 (C2V_23_297),
	.C2V_8 (C2V_23_364),
	.C2V_9 (C2V_23_443),
	.C2V_10 (C2V_23_677),
	.C2V_11 (C2V_23_741),
	.C2V_12 (C2V_23_795),
	.C2V_13 (C2V_23_873),
	.C2V_14 (C2V_23_921),
	.C2V_15 (C2V_23_964),
	.C2V_16 (C2V_23_1016),
	.C2V_17 (C2V_23_1065),
	.C2V_18 (C2V_23_1113),
	.C2V_19 (C2V_23_1174),
	.C2V_20 (C2V_23_1175),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU24 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_33_24),
	.V2C_2 (V2C_57_24),
	.V2C_3 (V2C_97_24),
	.V2C_4 (V2C_165_24),
	.V2C_5 (V2C_199_24),
	.V2C_6 (V2C_278_24),
	.V2C_7 (V2C_331_24),
	.V2C_8 (V2C_435_24),
	.V2C_9 (V2C_532_24),
	.V2C_10 (V2C_613_24),
	.V2C_11 (V2C_769_24),
	.V2C_12 (V2C_845_24),
	.V2C_13 (V2C_878_24),
	.V2C_14 (V2C_940_24),
	.V2C_15 (V2C_975_24),
	.V2C_16 (V2C_1042_24),
	.V2C_17 (V2C_1058_24),
	.V2C_18 (V2C_1108_24),
	.V2C_19 (V2C_1175_24),
	.V2C_20 (V2C_1176_24),
	.C2V_1 (C2V_24_33),
	.C2V_2 (C2V_24_57),
	.C2V_3 (C2V_24_97),
	.C2V_4 (C2V_24_165),
	.C2V_5 (C2V_24_199),
	.C2V_6 (C2V_24_278),
	.C2V_7 (C2V_24_331),
	.C2V_8 (C2V_24_435),
	.C2V_9 (C2V_24_532),
	.C2V_10 (C2V_24_613),
	.C2V_11 (C2V_24_769),
	.C2V_12 (C2V_24_845),
	.C2V_13 (C2V_24_878),
	.C2V_14 (C2V_24_940),
	.C2V_15 (C2V_24_975),
	.C2V_16 (C2V_24_1042),
	.C2V_17 (C2V_24_1058),
	.C2V_18 (C2V_24_1108),
	.C2V_19 (C2V_24_1175),
	.C2V_20 (C2V_24_1176),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU25 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_9_25),
	.V2C_2 (V2C_93_25),
	.V2C_3 (V2C_113_25),
	.V2C_4 (V2C_174_25),
	.V2C_5 (V2C_236_25),
	.V2C_6 (V2C_279_25),
	.V2C_7 (V2C_379_25),
	.V2C_8 (V2C_385_25),
	.V2C_9 (V2C_482_25),
	.V2C_10 (V2C_766_25),
	.V2C_11 (V2C_814_25),
	.V2C_12 (V2C_862_25),
	.V2C_13 (V2C_903_25),
	.V2C_14 (V2C_944_25),
	.V2C_15 (V2C_978_25),
	.V2C_16 (V2C_1017_25),
	.V2C_17 (V2C_1091_25),
	.V2C_18 (V2C_1150_25),
	.V2C_19 (V2C_1176_25),
	.V2C_20 (V2C_1177_25),
	.C2V_1 (C2V_25_9),
	.C2V_2 (C2V_25_93),
	.C2V_3 (C2V_25_113),
	.C2V_4 (C2V_25_174),
	.C2V_5 (C2V_25_236),
	.C2V_6 (C2V_25_279),
	.C2V_7 (C2V_25_379),
	.C2V_8 (C2V_25_385),
	.C2V_9 (C2V_25_482),
	.C2V_10 (C2V_25_766),
	.C2V_11 (C2V_25_814),
	.C2V_12 (C2V_25_862),
	.C2V_13 (C2V_25_903),
	.C2V_14 (C2V_25_944),
	.C2V_15 (C2V_25_978),
	.C2V_16 (C2V_25_1017),
	.C2V_17 (C2V_25_1091),
	.C2V_18 (C2V_25_1150),
	.C2V_19 (C2V_25_1176),
	.C2V_20 (C2V_25_1177),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU26 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_18_26),
	.V2C_2 (V2C_67_26),
	.V2C_3 (V2C_123_26),
	.V2C_4 (V2C_171_26),
	.V2C_5 (V2C_200_26),
	.V2C_6 (V2C_269_26),
	.V2C_7 (V2C_320_26),
	.V2C_8 (V2C_427_26),
	.V2C_9 (V2C_516_26),
	.V2C_10 (V2C_628_26),
	.V2C_11 (V2C_689_26),
	.V2C_12 (V2C_857_26),
	.V2C_13 (V2C_899_26),
	.V2C_14 (V2C_914_26),
	.V2C_15 (V2C_993_26),
	.V2C_16 (V2C_1025_26),
	.V2C_17 (V2C_1092_26),
	.V2C_18 (V2C_1123_26),
	.V2C_19 (V2C_1177_26),
	.V2C_20 (V2C_1178_26),
	.C2V_1 (C2V_26_18),
	.C2V_2 (C2V_26_67),
	.C2V_3 (C2V_26_123),
	.C2V_4 (C2V_26_171),
	.C2V_5 (C2V_26_200),
	.C2V_6 (C2V_26_269),
	.C2V_7 (C2V_26_320),
	.C2V_8 (C2V_26_427),
	.C2V_9 (C2V_26_516),
	.C2V_10 (C2V_26_628),
	.C2V_11 (C2V_26_689),
	.C2V_12 (C2V_26_857),
	.C2V_13 (C2V_26_899),
	.C2V_14 (C2V_26_914),
	.C2V_15 (C2V_26_993),
	.C2V_16 (C2V_26_1025),
	.C2V_17 (C2V_26_1092),
	.C2V_18 (C2V_26_1123),
	.C2V_19 (C2V_26_1177),
	.C2V_20 (C2V_26_1178),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU27 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_13_27),
	.V2C_2 (V2C_88_27),
	.V2C_3 (V2C_105_27),
	.V2C_4 (V2C_187_27),
	.V2C_5 (V2C_205_27),
	.V2C_6 (V2C_272_27),
	.V2C_7 (V2C_369_27),
	.V2C_8 (V2C_424_27),
	.V2C_9 (V2C_535_27),
	.V2C_10 (V2C_592_27),
	.V2C_11 (V2C_668_27),
	.V2C_12 (V2C_724_27),
	.V2C_13 (V2C_903_27),
	.V2C_14 (V2C_947_27),
	.V2C_15 (V2C_972_27),
	.V2C_16 (V2C_1032_27),
	.V2C_17 (V2C_1062_27),
	.V2C_18 (V2C_1107_27),
	.V2C_19 (V2C_1178_27),
	.V2C_20 (V2C_1179_27),
	.C2V_1 (C2V_27_13),
	.C2V_2 (C2V_27_88),
	.C2V_3 (C2V_27_105),
	.C2V_4 (C2V_27_187),
	.C2V_5 (C2V_27_205),
	.C2V_6 (C2V_27_272),
	.C2V_7 (C2V_27_369),
	.C2V_8 (C2V_27_424),
	.C2V_9 (C2V_27_535),
	.C2V_10 (C2V_27_592),
	.C2V_11 (C2V_27_668),
	.C2V_12 (C2V_27_724),
	.C2V_13 (C2V_27_903),
	.C2V_14 (C2V_27_947),
	.C2V_15 (C2V_27_972),
	.C2V_16 (C2V_27_1032),
	.C2V_17 (C2V_27_1062),
	.C2V_18 (C2V_27_1107),
	.C2V_19 (C2V_27_1178),
	.C2V_20 (C2V_27_1179),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU28 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_32_28),
	.V2C_2 (V2C_91_28),
	.V2C_3 (V2C_130_28),
	.V2C_4 (V2C_186_28),
	.V2C_5 (V2C_203_28),
	.V2C_6 (V2C_257_28),
	.V2C_7 (V2C_433_28),
	.V2C_8 (V2C_521_28),
	.V2C_9 (V2C_557_28),
	.V2C_10 (V2C_619_28),
	.V2C_11 (V2C_644_28),
	.V2C_12 (V2C_690_28),
	.V2C_13 (V2C_907_28),
	.V2C_14 (V2C_931_28),
	.V2C_15 (V2C_967_28),
	.V2C_16 (V2C_1045_28),
	.V2C_17 (V2C_1072_28),
	.V2C_18 (V2C_1136_28),
	.V2C_19 (V2C_1179_28),
	.V2C_20 (V2C_1180_28),
	.C2V_1 (C2V_28_32),
	.C2V_2 (C2V_28_91),
	.C2V_3 (C2V_28_130),
	.C2V_4 (C2V_28_186),
	.C2V_5 (C2V_28_203),
	.C2V_6 (C2V_28_257),
	.C2V_7 (C2V_28_433),
	.C2V_8 (C2V_28_521),
	.C2V_9 (C2V_28_557),
	.C2V_10 (C2V_28_619),
	.C2V_11 (C2V_28_644),
	.C2V_12 (C2V_28_690),
	.C2V_13 (C2V_28_907),
	.C2V_14 (C2V_28_931),
	.C2V_15 (C2V_28_967),
	.C2V_16 (C2V_28_1045),
	.C2V_17 (C2V_28_1072),
	.C2V_18 (C2V_28_1136),
	.C2V_19 (C2V_28_1179),
	.C2V_20 (C2V_28_1180),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU29 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_3_29),
	.V2C_2 (V2C_61_29),
	.V2C_3 (V2C_144_29),
	.V2C_4 (V2C_167_29),
	.V2C_5 (V2C_231_29),
	.V2C_6 (V2C_249_29),
	.V2C_7 (V2C_298_29),
	.V2C_8 (V2C_365_29),
	.V2C_9 (V2C_444_29),
	.V2C_10 (V2C_678_29),
	.V2C_11 (V2C_742_29),
	.V2C_12 (V2C_796_29),
	.V2C_13 (V2C_874_29),
	.V2C_14 (V2C_922_29),
	.V2C_15 (V2C_965_29),
	.V2C_16 (V2C_1017_29),
	.V2C_17 (V2C_1066_29),
	.V2C_18 (V2C_1114_29),
	.V2C_19 (V2C_1180_29),
	.V2C_20 (V2C_1181_29),
	.C2V_1 (C2V_29_3),
	.C2V_2 (C2V_29_61),
	.C2V_3 (C2V_29_144),
	.C2V_4 (C2V_29_167),
	.C2V_5 (C2V_29_231),
	.C2V_6 (C2V_29_249),
	.C2V_7 (C2V_29_298),
	.C2V_8 (C2V_29_365),
	.C2V_9 (C2V_29_444),
	.C2V_10 (C2V_29_678),
	.C2V_11 (C2V_29_742),
	.C2V_12 (C2V_29_796),
	.C2V_13 (C2V_29_874),
	.C2V_14 (C2V_29_922),
	.C2V_15 (C2V_29_965),
	.C2V_16 (C2V_29_1017),
	.C2V_17 (C2V_29_1066),
	.C2V_18 (C2V_29_1114),
	.C2V_19 (C2V_29_1180),
	.C2V_20 (C2V_29_1181),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU30 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_34_30),
	.V2C_2 (V2C_58_30),
	.V2C_3 (V2C_98_30),
	.V2C_4 (V2C_166_30),
	.V2C_5 (V2C_200_30),
	.V2C_6 (V2C_279_30),
	.V2C_7 (V2C_332_30),
	.V2C_8 (V2C_436_30),
	.V2C_9 (V2C_533_30),
	.V2C_10 (V2C_614_30),
	.V2C_11 (V2C_770_30),
	.V2C_12 (V2C_846_30),
	.V2C_13 (V2C_879_30),
	.V2C_14 (V2C_941_30),
	.V2C_15 (V2C_976_30),
	.V2C_16 (V2C_1043_30),
	.V2C_17 (V2C_1059_30),
	.V2C_18 (V2C_1109_30),
	.V2C_19 (V2C_1181_30),
	.V2C_20 (V2C_1182_30),
	.C2V_1 (C2V_30_34),
	.C2V_2 (C2V_30_58),
	.C2V_3 (C2V_30_98),
	.C2V_4 (C2V_30_166),
	.C2V_5 (C2V_30_200),
	.C2V_6 (C2V_30_279),
	.C2V_7 (C2V_30_332),
	.C2V_8 (C2V_30_436),
	.C2V_9 (C2V_30_533),
	.C2V_10 (C2V_30_614),
	.C2V_11 (C2V_30_770),
	.C2V_12 (C2V_30_846),
	.C2V_13 (C2V_30_879),
	.C2V_14 (C2V_30_941),
	.C2V_15 (C2V_30_976),
	.C2V_16 (C2V_30_1043),
	.C2V_17 (C2V_30_1059),
	.C2V_18 (C2V_30_1109),
	.C2V_19 (C2V_30_1181),
	.C2V_20 (C2V_30_1182),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU31 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_10_31),
	.V2C_2 (V2C_94_31),
	.V2C_3 (V2C_114_31),
	.V2C_4 (V2C_175_31),
	.V2C_5 (V2C_237_31),
	.V2C_6 (V2C_280_31),
	.V2C_7 (V2C_380_31),
	.V2C_8 (V2C_386_31),
	.V2C_9 (V2C_483_31),
	.V2C_10 (V2C_767_31),
	.V2C_11 (V2C_815_31),
	.V2C_12 (V2C_863_31),
	.V2C_13 (V2C_904_31),
	.V2C_14 (V2C_945_31),
	.V2C_15 (V2C_979_31),
	.V2C_16 (V2C_1018_31),
	.V2C_17 (V2C_1092_31),
	.V2C_18 (V2C_1151_31),
	.V2C_19 (V2C_1182_31),
	.V2C_20 (V2C_1183_31),
	.C2V_1 (C2V_31_10),
	.C2V_2 (C2V_31_94),
	.C2V_3 (C2V_31_114),
	.C2V_4 (C2V_31_175),
	.C2V_5 (C2V_31_237),
	.C2V_6 (C2V_31_280),
	.C2V_7 (C2V_31_380),
	.C2V_8 (C2V_31_386),
	.C2V_9 (C2V_31_483),
	.C2V_10 (C2V_31_767),
	.C2V_11 (C2V_31_815),
	.C2V_12 (C2V_31_863),
	.C2V_13 (C2V_31_904),
	.C2V_14 (C2V_31_945),
	.C2V_15 (C2V_31_979),
	.C2V_16 (C2V_31_1018),
	.C2V_17 (C2V_31_1092),
	.C2V_18 (C2V_31_1151),
	.C2V_19 (C2V_31_1182),
	.C2V_20 (C2V_31_1183),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU32 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_19_32),
	.V2C_2 (V2C_68_32),
	.V2C_3 (V2C_124_32),
	.V2C_4 (V2C_172_32),
	.V2C_5 (V2C_201_32),
	.V2C_6 (V2C_270_32),
	.V2C_7 (V2C_321_32),
	.V2C_8 (V2C_428_32),
	.V2C_9 (V2C_517_32),
	.V2C_10 (V2C_629_32),
	.V2C_11 (V2C_690_32),
	.V2C_12 (V2C_858_32),
	.V2C_13 (V2C_900_32),
	.V2C_14 (V2C_915_32),
	.V2C_15 (V2C_994_32),
	.V2C_16 (V2C_1026_32),
	.V2C_17 (V2C_1093_32),
	.V2C_18 (V2C_1124_32),
	.V2C_19 (V2C_1183_32),
	.V2C_20 (V2C_1184_32),
	.C2V_1 (C2V_32_19),
	.C2V_2 (C2V_32_68),
	.C2V_3 (C2V_32_124),
	.C2V_4 (C2V_32_172),
	.C2V_5 (C2V_32_201),
	.C2V_6 (C2V_32_270),
	.C2V_7 (C2V_32_321),
	.C2V_8 (C2V_32_428),
	.C2V_9 (C2V_32_517),
	.C2V_10 (C2V_32_629),
	.C2V_11 (C2V_32_690),
	.C2V_12 (C2V_32_858),
	.C2V_13 (C2V_32_900),
	.C2V_14 (C2V_32_915),
	.C2V_15 (C2V_32_994),
	.C2V_16 (C2V_32_1026),
	.C2V_17 (C2V_32_1093),
	.C2V_18 (C2V_32_1124),
	.C2V_19 (C2V_32_1183),
	.C2V_20 (C2V_32_1184),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU33 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_14_33),
	.V2C_2 (V2C_89_33),
	.V2C_3 (V2C_106_33),
	.V2C_4 (V2C_188_33),
	.V2C_5 (V2C_206_33),
	.V2C_6 (V2C_273_33),
	.V2C_7 (V2C_370_33),
	.V2C_8 (V2C_425_33),
	.V2C_9 (V2C_536_33),
	.V2C_10 (V2C_593_33),
	.V2C_11 (V2C_669_33),
	.V2C_12 (V2C_725_33),
	.V2C_13 (V2C_904_33),
	.V2C_14 (V2C_948_33),
	.V2C_15 (V2C_973_33),
	.V2C_16 (V2C_1033_33),
	.V2C_17 (V2C_1063_33),
	.V2C_18 (V2C_1108_33),
	.V2C_19 (V2C_1184_33),
	.V2C_20 (V2C_1185_33),
	.C2V_1 (C2V_33_14),
	.C2V_2 (C2V_33_89),
	.C2V_3 (C2V_33_106),
	.C2V_4 (C2V_33_188),
	.C2V_5 (C2V_33_206),
	.C2V_6 (C2V_33_273),
	.C2V_7 (C2V_33_370),
	.C2V_8 (C2V_33_425),
	.C2V_9 (C2V_33_536),
	.C2V_10 (C2V_33_593),
	.C2V_11 (C2V_33_669),
	.C2V_12 (C2V_33_725),
	.C2V_13 (C2V_33_904),
	.C2V_14 (C2V_33_948),
	.C2V_15 (C2V_33_973),
	.C2V_16 (C2V_33_1033),
	.C2V_17 (C2V_33_1063),
	.C2V_18 (C2V_33_1108),
	.C2V_19 (C2V_33_1184),
	.C2V_20 (C2V_33_1185),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU34 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_33_34),
	.V2C_2 (V2C_92_34),
	.V2C_3 (V2C_131_34),
	.V2C_4 (V2C_187_34),
	.V2C_5 (V2C_204_34),
	.V2C_6 (V2C_258_34),
	.V2C_7 (V2C_434_34),
	.V2C_8 (V2C_522_34),
	.V2C_9 (V2C_558_34),
	.V2C_10 (V2C_620_34),
	.V2C_11 (V2C_645_34),
	.V2C_12 (V2C_691_34),
	.V2C_13 (V2C_908_34),
	.V2C_14 (V2C_932_34),
	.V2C_15 (V2C_968_34),
	.V2C_16 (V2C_1046_34),
	.V2C_17 (V2C_1073_34),
	.V2C_18 (V2C_1137_34),
	.V2C_19 (V2C_1185_34),
	.V2C_20 (V2C_1186_34),
	.C2V_1 (C2V_34_33),
	.C2V_2 (C2V_34_92),
	.C2V_3 (C2V_34_131),
	.C2V_4 (C2V_34_187),
	.C2V_5 (C2V_34_204),
	.C2V_6 (C2V_34_258),
	.C2V_7 (C2V_34_434),
	.C2V_8 (C2V_34_522),
	.C2V_9 (C2V_34_558),
	.C2V_10 (C2V_34_620),
	.C2V_11 (C2V_34_645),
	.C2V_12 (C2V_34_691),
	.C2V_13 (C2V_34_908),
	.C2V_14 (C2V_34_932),
	.C2V_15 (C2V_34_968),
	.C2V_16 (C2V_34_1046),
	.C2V_17 (C2V_34_1073),
	.C2V_18 (C2V_34_1137),
	.C2V_19 (C2V_34_1185),
	.C2V_20 (C2V_34_1186),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU35 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_4_35),
	.V2C_2 (V2C_62_35),
	.V2C_3 (V2C_97_35),
	.V2C_4 (V2C_168_35),
	.V2C_5 (V2C_232_35),
	.V2C_6 (V2C_250_35),
	.V2C_7 (V2C_299_35),
	.V2C_8 (V2C_366_35),
	.V2C_9 (V2C_445_35),
	.V2C_10 (V2C_679_35),
	.V2C_11 (V2C_743_35),
	.V2C_12 (V2C_797_35),
	.V2C_13 (V2C_875_35),
	.V2C_14 (V2C_923_35),
	.V2C_15 (V2C_966_35),
	.V2C_16 (V2C_1018_35),
	.V2C_17 (V2C_1067_35),
	.V2C_18 (V2C_1115_35),
	.V2C_19 (V2C_1186_35),
	.V2C_20 (V2C_1187_35),
	.C2V_1 (C2V_35_4),
	.C2V_2 (C2V_35_62),
	.C2V_3 (C2V_35_97),
	.C2V_4 (C2V_35_168),
	.C2V_5 (C2V_35_232),
	.C2V_6 (C2V_35_250),
	.C2V_7 (C2V_35_299),
	.C2V_8 (C2V_35_366),
	.C2V_9 (C2V_35_445),
	.C2V_10 (C2V_35_679),
	.C2V_11 (C2V_35_743),
	.C2V_12 (C2V_35_797),
	.C2V_13 (C2V_35_875),
	.C2V_14 (C2V_35_923),
	.C2V_15 (C2V_35_966),
	.C2V_16 (C2V_35_1018),
	.C2V_17 (C2V_35_1067),
	.C2V_18 (C2V_35_1115),
	.C2V_19 (C2V_35_1186),
	.C2V_20 (C2V_35_1187),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU36 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_35_36),
	.V2C_2 (V2C_59_36),
	.V2C_3 (V2C_99_36),
	.V2C_4 (V2C_167_36),
	.V2C_5 (V2C_201_36),
	.V2C_6 (V2C_280_36),
	.V2C_7 (V2C_333_36),
	.V2C_8 (V2C_437_36),
	.V2C_9 (V2C_534_36),
	.V2C_10 (V2C_615_36),
	.V2C_11 (V2C_771_36),
	.V2C_12 (V2C_847_36),
	.V2C_13 (V2C_880_36),
	.V2C_14 (V2C_942_36),
	.V2C_15 (V2C_977_36),
	.V2C_16 (V2C_1044_36),
	.V2C_17 (V2C_1060_36),
	.V2C_18 (V2C_1110_36),
	.V2C_19 (V2C_1187_36),
	.V2C_20 (V2C_1188_36),
	.C2V_1 (C2V_36_35),
	.C2V_2 (C2V_36_59),
	.C2V_3 (C2V_36_99),
	.C2V_4 (C2V_36_167),
	.C2V_5 (C2V_36_201),
	.C2V_6 (C2V_36_280),
	.C2V_7 (C2V_36_333),
	.C2V_8 (C2V_36_437),
	.C2V_9 (C2V_36_534),
	.C2V_10 (C2V_36_615),
	.C2V_11 (C2V_36_771),
	.C2V_12 (C2V_36_847),
	.C2V_13 (C2V_36_880),
	.C2V_14 (C2V_36_942),
	.C2V_15 (C2V_36_977),
	.C2V_16 (C2V_36_1044),
	.C2V_17 (C2V_36_1060),
	.C2V_18 (C2V_36_1110),
	.C2V_19 (C2V_36_1187),
	.C2V_20 (C2V_36_1188),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU37 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_11_37),
	.V2C_2 (V2C_95_37),
	.V2C_3 (V2C_115_37),
	.V2C_4 (V2C_176_37),
	.V2C_5 (V2C_238_37),
	.V2C_6 (V2C_281_37),
	.V2C_7 (V2C_381_37),
	.V2C_8 (V2C_387_37),
	.V2C_9 (V2C_484_37),
	.V2C_10 (V2C_768_37),
	.V2C_11 (V2C_816_37),
	.V2C_12 (V2C_864_37),
	.V2C_13 (V2C_905_37),
	.V2C_14 (V2C_946_37),
	.V2C_15 (V2C_980_37),
	.V2C_16 (V2C_1019_37),
	.V2C_17 (V2C_1093_37),
	.V2C_18 (V2C_1152_37),
	.V2C_19 (V2C_1188_37),
	.V2C_20 (V2C_1189_37),
	.C2V_1 (C2V_37_11),
	.C2V_2 (C2V_37_95),
	.C2V_3 (C2V_37_115),
	.C2V_4 (C2V_37_176),
	.C2V_5 (C2V_37_238),
	.C2V_6 (C2V_37_281),
	.C2V_7 (C2V_37_381),
	.C2V_8 (C2V_37_387),
	.C2V_9 (C2V_37_484),
	.C2V_10 (C2V_37_768),
	.C2V_11 (C2V_37_816),
	.C2V_12 (C2V_37_864),
	.C2V_13 (C2V_37_905),
	.C2V_14 (C2V_37_946),
	.C2V_15 (C2V_37_980),
	.C2V_16 (C2V_37_1019),
	.C2V_17 (C2V_37_1093),
	.C2V_18 (C2V_37_1152),
	.C2V_19 (C2V_37_1188),
	.C2V_20 (C2V_37_1189),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU38 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_20_38),
	.V2C_2 (V2C_69_38),
	.V2C_3 (V2C_125_38),
	.V2C_4 (V2C_173_38),
	.V2C_5 (V2C_202_38),
	.V2C_6 (V2C_271_38),
	.V2C_7 (V2C_322_38),
	.V2C_8 (V2C_429_38),
	.V2C_9 (V2C_518_38),
	.V2C_10 (V2C_630_38),
	.V2C_11 (V2C_691_38),
	.V2C_12 (V2C_859_38),
	.V2C_13 (V2C_901_38),
	.V2C_14 (V2C_916_38),
	.V2C_15 (V2C_995_38),
	.V2C_16 (V2C_1027_38),
	.V2C_17 (V2C_1094_38),
	.V2C_18 (V2C_1125_38),
	.V2C_19 (V2C_1189_38),
	.V2C_20 (V2C_1190_38),
	.C2V_1 (C2V_38_20),
	.C2V_2 (C2V_38_69),
	.C2V_3 (C2V_38_125),
	.C2V_4 (C2V_38_173),
	.C2V_5 (C2V_38_202),
	.C2V_6 (C2V_38_271),
	.C2V_7 (C2V_38_322),
	.C2V_8 (C2V_38_429),
	.C2V_9 (C2V_38_518),
	.C2V_10 (C2V_38_630),
	.C2V_11 (C2V_38_691),
	.C2V_12 (C2V_38_859),
	.C2V_13 (C2V_38_901),
	.C2V_14 (C2V_38_916),
	.C2V_15 (C2V_38_995),
	.C2V_16 (C2V_38_1027),
	.C2V_17 (C2V_38_1094),
	.C2V_18 (C2V_38_1125),
	.C2V_19 (C2V_38_1189),
	.C2V_20 (C2V_38_1190),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU39 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_15_39),
	.V2C_2 (V2C_90_39),
	.V2C_3 (V2C_107_39),
	.V2C_4 (V2C_189_39),
	.V2C_5 (V2C_207_39),
	.V2C_6 (V2C_274_39),
	.V2C_7 (V2C_371_39),
	.V2C_8 (V2C_426_39),
	.V2C_9 (V2C_537_39),
	.V2C_10 (V2C_594_39),
	.V2C_11 (V2C_670_39),
	.V2C_12 (V2C_726_39),
	.V2C_13 (V2C_905_39),
	.V2C_14 (V2C_949_39),
	.V2C_15 (V2C_974_39),
	.V2C_16 (V2C_1034_39),
	.V2C_17 (V2C_1064_39),
	.V2C_18 (V2C_1109_39),
	.V2C_19 (V2C_1190_39),
	.V2C_20 (V2C_1191_39),
	.C2V_1 (C2V_39_15),
	.C2V_2 (C2V_39_90),
	.C2V_3 (C2V_39_107),
	.C2V_4 (C2V_39_189),
	.C2V_5 (C2V_39_207),
	.C2V_6 (C2V_39_274),
	.C2V_7 (C2V_39_371),
	.C2V_8 (C2V_39_426),
	.C2V_9 (C2V_39_537),
	.C2V_10 (C2V_39_594),
	.C2V_11 (C2V_39_670),
	.C2V_12 (C2V_39_726),
	.C2V_13 (C2V_39_905),
	.C2V_14 (C2V_39_949),
	.C2V_15 (C2V_39_974),
	.C2V_16 (C2V_39_1034),
	.C2V_17 (C2V_39_1064),
	.C2V_18 (C2V_39_1109),
	.C2V_19 (C2V_39_1190),
	.C2V_20 (C2V_39_1191),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU40 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_34_40),
	.V2C_2 (V2C_93_40),
	.V2C_3 (V2C_132_40),
	.V2C_4 (V2C_188_40),
	.V2C_5 (V2C_205_40),
	.V2C_6 (V2C_259_40),
	.V2C_7 (V2C_435_40),
	.V2C_8 (V2C_523_40),
	.V2C_9 (V2C_559_40),
	.V2C_10 (V2C_621_40),
	.V2C_11 (V2C_646_40),
	.V2C_12 (V2C_692_40),
	.V2C_13 (V2C_909_40),
	.V2C_14 (V2C_933_40),
	.V2C_15 (V2C_969_40),
	.V2C_16 (V2C_1047_40),
	.V2C_17 (V2C_1074_40),
	.V2C_18 (V2C_1138_40),
	.V2C_19 (V2C_1191_40),
	.V2C_20 (V2C_1192_40),
	.C2V_1 (C2V_40_34),
	.C2V_2 (C2V_40_93),
	.C2V_3 (C2V_40_132),
	.C2V_4 (C2V_40_188),
	.C2V_5 (C2V_40_205),
	.C2V_6 (C2V_40_259),
	.C2V_7 (C2V_40_435),
	.C2V_8 (C2V_40_523),
	.C2V_9 (C2V_40_559),
	.C2V_10 (C2V_40_621),
	.C2V_11 (C2V_40_646),
	.C2V_12 (C2V_40_692),
	.C2V_13 (C2V_40_909),
	.C2V_14 (C2V_40_933),
	.C2V_15 (C2V_40_969),
	.C2V_16 (C2V_40_1047),
	.C2V_17 (C2V_40_1074),
	.C2V_18 (C2V_40_1138),
	.C2V_19 (C2V_40_1191),
	.C2V_20 (C2V_40_1192),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU41 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_5_41),
	.V2C_2 (V2C_63_41),
	.V2C_3 (V2C_98_41),
	.V2C_4 (V2C_169_41),
	.V2C_5 (V2C_233_41),
	.V2C_6 (V2C_251_41),
	.V2C_7 (V2C_300_41),
	.V2C_8 (V2C_367_41),
	.V2C_9 (V2C_446_41),
	.V2C_10 (V2C_680_41),
	.V2C_11 (V2C_744_41),
	.V2C_12 (V2C_798_41),
	.V2C_13 (V2C_876_41),
	.V2C_14 (V2C_924_41),
	.V2C_15 (V2C_967_41),
	.V2C_16 (V2C_1019_41),
	.V2C_17 (V2C_1068_41),
	.V2C_18 (V2C_1116_41),
	.V2C_19 (V2C_1192_41),
	.V2C_20 (V2C_1193_41),
	.C2V_1 (C2V_41_5),
	.C2V_2 (C2V_41_63),
	.C2V_3 (C2V_41_98),
	.C2V_4 (C2V_41_169),
	.C2V_5 (C2V_41_233),
	.C2V_6 (C2V_41_251),
	.C2V_7 (C2V_41_300),
	.C2V_8 (C2V_41_367),
	.C2V_9 (C2V_41_446),
	.C2V_10 (C2V_41_680),
	.C2V_11 (C2V_41_744),
	.C2V_12 (C2V_41_798),
	.C2V_13 (C2V_41_876),
	.C2V_14 (C2V_41_924),
	.C2V_15 (C2V_41_967),
	.C2V_16 (C2V_41_1019),
	.C2V_17 (C2V_41_1068),
	.C2V_18 (C2V_41_1116),
	.C2V_19 (C2V_41_1192),
	.C2V_20 (C2V_41_1193),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU42 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_36_42),
	.V2C_2 (V2C_60_42),
	.V2C_3 (V2C_100_42),
	.V2C_4 (V2C_168_42),
	.V2C_5 (V2C_202_42),
	.V2C_6 (V2C_281_42),
	.V2C_7 (V2C_334_42),
	.V2C_8 (V2C_438_42),
	.V2C_9 (V2C_535_42),
	.V2C_10 (V2C_616_42),
	.V2C_11 (V2C_772_42),
	.V2C_12 (V2C_848_42),
	.V2C_13 (V2C_881_42),
	.V2C_14 (V2C_943_42),
	.V2C_15 (V2C_978_42),
	.V2C_16 (V2C_1045_42),
	.V2C_17 (V2C_1061_42),
	.V2C_18 (V2C_1111_42),
	.V2C_19 (V2C_1193_42),
	.V2C_20 (V2C_1194_42),
	.C2V_1 (C2V_42_36),
	.C2V_2 (C2V_42_60),
	.C2V_3 (C2V_42_100),
	.C2V_4 (C2V_42_168),
	.C2V_5 (C2V_42_202),
	.C2V_6 (C2V_42_281),
	.C2V_7 (C2V_42_334),
	.C2V_8 (C2V_42_438),
	.C2V_9 (C2V_42_535),
	.C2V_10 (C2V_42_616),
	.C2V_11 (C2V_42_772),
	.C2V_12 (C2V_42_848),
	.C2V_13 (C2V_42_881),
	.C2V_14 (C2V_42_943),
	.C2V_15 (C2V_42_978),
	.C2V_16 (C2V_42_1045),
	.C2V_17 (C2V_42_1061),
	.C2V_18 (C2V_42_1111),
	.C2V_19 (C2V_42_1193),
	.C2V_20 (C2V_42_1194),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU43 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_12_43),
	.V2C_2 (V2C_96_43),
	.V2C_3 (V2C_116_43),
	.V2C_4 (V2C_177_43),
	.V2C_5 (V2C_239_43),
	.V2C_6 (V2C_282_43),
	.V2C_7 (V2C_382_43),
	.V2C_8 (V2C_388_43),
	.V2C_9 (V2C_485_43),
	.V2C_10 (V2C_721_43),
	.V2C_11 (V2C_769_43),
	.V2C_12 (V2C_817_43),
	.V2C_13 (V2C_906_43),
	.V2C_14 (V2C_947_43),
	.V2C_15 (V2C_981_43),
	.V2C_16 (V2C_1020_43),
	.V2C_17 (V2C_1094_43),
	.V2C_18 (V2C_1105_43),
	.V2C_19 (V2C_1194_43),
	.V2C_20 (V2C_1195_43),
	.C2V_1 (C2V_43_12),
	.C2V_2 (C2V_43_96),
	.C2V_3 (C2V_43_116),
	.C2V_4 (C2V_43_177),
	.C2V_5 (C2V_43_239),
	.C2V_6 (C2V_43_282),
	.C2V_7 (C2V_43_382),
	.C2V_8 (C2V_43_388),
	.C2V_9 (C2V_43_485),
	.C2V_10 (C2V_43_721),
	.C2V_11 (C2V_43_769),
	.C2V_12 (C2V_43_817),
	.C2V_13 (C2V_43_906),
	.C2V_14 (C2V_43_947),
	.C2V_15 (C2V_43_981),
	.C2V_16 (C2V_43_1020),
	.C2V_17 (C2V_43_1094),
	.C2V_18 (C2V_43_1105),
	.C2V_19 (C2V_43_1194),
	.C2V_20 (C2V_43_1195),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU44 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_21_44),
	.V2C_2 (V2C_70_44),
	.V2C_3 (V2C_126_44),
	.V2C_4 (V2C_174_44),
	.V2C_5 (V2C_203_44),
	.V2C_6 (V2C_272_44),
	.V2C_7 (V2C_323_44),
	.V2C_8 (V2C_430_44),
	.V2C_9 (V2C_519_44),
	.V2C_10 (V2C_631_44),
	.V2C_11 (V2C_692_44),
	.V2C_12 (V2C_860_44),
	.V2C_13 (V2C_902_44),
	.V2C_14 (V2C_917_44),
	.V2C_15 (V2C_996_44),
	.V2C_16 (V2C_1028_44),
	.V2C_17 (V2C_1095_44),
	.V2C_18 (V2C_1126_44),
	.V2C_19 (V2C_1195_44),
	.V2C_20 (V2C_1196_44),
	.C2V_1 (C2V_44_21),
	.C2V_2 (C2V_44_70),
	.C2V_3 (C2V_44_126),
	.C2V_4 (C2V_44_174),
	.C2V_5 (C2V_44_203),
	.C2V_6 (C2V_44_272),
	.C2V_7 (C2V_44_323),
	.C2V_8 (C2V_44_430),
	.C2V_9 (C2V_44_519),
	.C2V_10 (C2V_44_631),
	.C2V_11 (C2V_44_692),
	.C2V_12 (C2V_44_860),
	.C2V_13 (C2V_44_902),
	.C2V_14 (C2V_44_917),
	.C2V_15 (C2V_44_996),
	.C2V_16 (C2V_44_1028),
	.C2V_17 (C2V_44_1095),
	.C2V_18 (C2V_44_1126),
	.C2V_19 (C2V_44_1195),
	.C2V_20 (C2V_44_1196),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU45 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_16_45),
	.V2C_2 (V2C_91_45),
	.V2C_3 (V2C_108_45),
	.V2C_4 (V2C_190_45),
	.V2C_5 (V2C_208_45),
	.V2C_6 (V2C_275_45),
	.V2C_7 (V2C_372_45),
	.V2C_8 (V2C_427_45),
	.V2C_9 (V2C_538_45),
	.V2C_10 (V2C_595_45),
	.V2C_11 (V2C_671_45),
	.V2C_12 (V2C_727_45),
	.V2C_13 (V2C_906_45),
	.V2C_14 (V2C_950_45),
	.V2C_15 (V2C_975_45),
	.V2C_16 (V2C_1035_45),
	.V2C_17 (V2C_1065_45),
	.V2C_18 (V2C_1110_45),
	.V2C_19 (V2C_1196_45),
	.V2C_20 (V2C_1197_45),
	.C2V_1 (C2V_45_16),
	.C2V_2 (C2V_45_91),
	.C2V_3 (C2V_45_108),
	.C2V_4 (C2V_45_190),
	.C2V_5 (C2V_45_208),
	.C2V_6 (C2V_45_275),
	.C2V_7 (C2V_45_372),
	.C2V_8 (C2V_45_427),
	.C2V_9 (C2V_45_538),
	.C2V_10 (C2V_45_595),
	.C2V_11 (C2V_45_671),
	.C2V_12 (C2V_45_727),
	.C2V_13 (C2V_45_906),
	.C2V_14 (C2V_45_950),
	.C2V_15 (C2V_45_975),
	.C2V_16 (C2V_45_1035),
	.C2V_17 (C2V_45_1065),
	.C2V_18 (C2V_45_1110),
	.C2V_19 (C2V_45_1196),
	.C2V_20 (C2V_45_1197),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU46 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_35_46),
	.V2C_2 (V2C_94_46),
	.V2C_3 (V2C_133_46),
	.V2C_4 (V2C_189_46),
	.V2C_5 (V2C_206_46),
	.V2C_6 (V2C_260_46),
	.V2C_7 (V2C_436_46),
	.V2C_8 (V2C_524_46),
	.V2C_9 (V2C_560_46),
	.V2C_10 (V2C_622_46),
	.V2C_11 (V2C_647_46),
	.V2C_12 (V2C_693_46),
	.V2C_13 (V2C_910_46),
	.V2C_14 (V2C_934_46),
	.V2C_15 (V2C_970_46),
	.V2C_16 (V2C_1048_46),
	.V2C_17 (V2C_1075_46),
	.V2C_18 (V2C_1139_46),
	.V2C_19 (V2C_1197_46),
	.V2C_20 (V2C_1198_46),
	.C2V_1 (C2V_46_35),
	.C2V_2 (C2V_46_94),
	.C2V_3 (C2V_46_133),
	.C2V_4 (C2V_46_189),
	.C2V_5 (C2V_46_206),
	.C2V_6 (C2V_46_260),
	.C2V_7 (C2V_46_436),
	.C2V_8 (C2V_46_524),
	.C2V_9 (C2V_46_560),
	.C2V_10 (C2V_46_622),
	.C2V_11 (C2V_46_647),
	.C2V_12 (C2V_46_693),
	.C2V_13 (C2V_46_910),
	.C2V_14 (C2V_46_934),
	.C2V_15 (C2V_46_970),
	.C2V_16 (C2V_46_1048),
	.C2V_17 (C2V_46_1075),
	.C2V_18 (C2V_46_1139),
	.C2V_19 (C2V_46_1197),
	.C2V_20 (C2V_46_1198),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU47 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_6_47),
	.V2C_2 (V2C_64_47),
	.V2C_3 (V2C_99_47),
	.V2C_4 (V2C_170_47),
	.V2C_5 (V2C_234_47),
	.V2C_6 (V2C_252_47),
	.V2C_7 (V2C_301_47),
	.V2C_8 (V2C_368_47),
	.V2C_9 (V2C_447_47),
	.V2C_10 (V2C_681_47),
	.V2C_11 (V2C_745_47),
	.V2C_12 (V2C_799_47),
	.V2C_13 (V2C_877_47),
	.V2C_14 (V2C_925_47),
	.V2C_15 (V2C_968_47),
	.V2C_16 (V2C_1020_47),
	.V2C_17 (V2C_1069_47),
	.V2C_18 (V2C_1117_47),
	.V2C_19 (V2C_1198_47),
	.V2C_20 (V2C_1199_47),
	.C2V_1 (C2V_47_6),
	.C2V_2 (C2V_47_64),
	.C2V_3 (C2V_47_99),
	.C2V_4 (C2V_47_170),
	.C2V_5 (C2V_47_234),
	.C2V_6 (C2V_47_252),
	.C2V_7 (C2V_47_301),
	.C2V_8 (C2V_47_368),
	.C2V_9 (C2V_47_447),
	.C2V_10 (C2V_47_681),
	.C2V_11 (C2V_47_745),
	.C2V_12 (C2V_47_799),
	.C2V_13 (C2V_47_877),
	.C2V_14 (C2V_47_925),
	.C2V_15 (C2V_47_968),
	.C2V_16 (C2V_47_1020),
	.C2V_17 (C2V_47_1069),
	.C2V_18 (C2V_47_1117),
	.C2V_19 (C2V_47_1198),
	.C2V_20 (C2V_47_1199),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU48 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_37_48),
	.V2C_2 (V2C_61_48),
	.V2C_3 (V2C_101_48),
	.V2C_4 (V2C_169_48),
	.V2C_5 (V2C_203_48),
	.V2C_6 (V2C_282_48),
	.V2C_7 (V2C_335_48),
	.V2C_8 (V2C_439_48),
	.V2C_9 (V2C_536_48),
	.V2C_10 (V2C_617_48),
	.V2C_11 (V2C_773_48),
	.V2C_12 (V2C_849_48),
	.V2C_13 (V2C_882_48),
	.V2C_14 (V2C_944_48),
	.V2C_15 (V2C_979_48),
	.V2C_16 (V2C_1046_48),
	.V2C_17 (V2C_1062_48),
	.V2C_18 (V2C_1112_48),
	.V2C_19 (V2C_1199_48),
	.V2C_20 (V2C_1200_48),
	.C2V_1 (C2V_48_37),
	.C2V_2 (C2V_48_61),
	.C2V_3 (C2V_48_101),
	.C2V_4 (C2V_48_169),
	.C2V_5 (C2V_48_203),
	.C2V_6 (C2V_48_282),
	.C2V_7 (C2V_48_335),
	.C2V_8 (C2V_48_439),
	.C2V_9 (C2V_48_536),
	.C2V_10 (C2V_48_617),
	.C2V_11 (C2V_48_773),
	.C2V_12 (C2V_48_849),
	.C2V_13 (C2V_48_882),
	.C2V_14 (C2V_48_944),
	.C2V_15 (C2V_48_979),
	.C2V_16 (C2V_48_1046),
	.C2V_17 (C2V_48_1062),
	.C2V_18 (C2V_48_1112),
	.C2V_19 (C2V_48_1199),
	.C2V_20 (C2V_48_1200),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU49 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_13_49),
	.V2C_2 (V2C_49_49),
	.V2C_3 (V2C_117_49),
	.V2C_4 (V2C_178_49),
	.V2C_5 (V2C_240_49),
	.V2C_6 (V2C_283_49),
	.V2C_7 (V2C_383_49),
	.V2C_8 (V2C_389_49),
	.V2C_9 (V2C_486_49),
	.V2C_10 (V2C_722_49),
	.V2C_11 (V2C_770_49),
	.V2C_12 (V2C_818_49),
	.V2C_13 (V2C_907_49),
	.V2C_14 (V2C_948_49),
	.V2C_15 (V2C_982_49),
	.V2C_16 (V2C_1021_49),
	.V2C_17 (V2C_1095_49),
	.V2C_18 (V2C_1106_49),
	.V2C_19 (V2C_1200_49),
	.V2C_20 (V2C_1201_49),
	.C2V_1 (C2V_49_13),
	.C2V_2 (C2V_49_49),
	.C2V_3 (C2V_49_117),
	.C2V_4 (C2V_49_178),
	.C2V_5 (C2V_49_240),
	.C2V_6 (C2V_49_283),
	.C2V_7 (C2V_49_383),
	.C2V_8 (C2V_49_389),
	.C2V_9 (C2V_49_486),
	.C2V_10 (C2V_49_722),
	.C2V_11 (C2V_49_770),
	.C2V_12 (C2V_49_818),
	.C2V_13 (C2V_49_907),
	.C2V_14 (C2V_49_948),
	.C2V_15 (C2V_49_982),
	.C2V_16 (C2V_49_1021),
	.C2V_17 (C2V_49_1095),
	.C2V_18 (C2V_49_1106),
	.C2V_19 (C2V_49_1200),
	.C2V_20 (C2V_49_1201),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU50 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_22_50),
	.V2C_2 (V2C_71_50),
	.V2C_3 (V2C_127_50),
	.V2C_4 (V2C_175_50),
	.V2C_5 (V2C_204_50),
	.V2C_6 (V2C_273_50),
	.V2C_7 (V2C_324_50),
	.V2C_8 (V2C_431_50),
	.V2C_9 (V2C_520_50),
	.V2C_10 (V2C_632_50),
	.V2C_11 (V2C_693_50),
	.V2C_12 (V2C_861_50),
	.V2C_13 (V2C_903_50),
	.V2C_14 (V2C_918_50),
	.V2C_15 (V2C_997_50),
	.V2C_16 (V2C_1029_50),
	.V2C_17 (V2C_1096_50),
	.V2C_18 (V2C_1127_50),
	.V2C_19 (V2C_1201_50),
	.V2C_20 (V2C_1202_50),
	.C2V_1 (C2V_50_22),
	.C2V_2 (C2V_50_71),
	.C2V_3 (C2V_50_127),
	.C2V_4 (C2V_50_175),
	.C2V_5 (C2V_50_204),
	.C2V_6 (C2V_50_273),
	.C2V_7 (C2V_50_324),
	.C2V_8 (C2V_50_431),
	.C2V_9 (C2V_50_520),
	.C2V_10 (C2V_50_632),
	.C2V_11 (C2V_50_693),
	.C2V_12 (C2V_50_861),
	.C2V_13 (C2V_50_903),
	.C2V_14 (C2V_50_918),
	.C2V_15 (C2V_50_997),
	.C2V_16 (C2V_50_1029),
	.C2V_17 (C2V_50_1096),
	.C2V_18 (C2V_50_1127),
	.C2V_19 (C2V_50_1201),
	.C2V_20 (C2V_50_1202),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU51 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_17_51),
	.V2C_2 (V2C_92_51),
	.V2C_3 (V2C_109_51),
	.V2C_4 (V2C_191_51),
	.V2C_5 (V2C_209_51),
	.V2C_6 (V2C_276_51),
	.V2C_7 (V2C_373_51),
	.V2C_8 (V2C_428_51),
	.V2C_9 (V2C_539_51),
	.V2C_10 (V2C_596_51),
	.V2C_11 (V2C_672_51),
	.V2C_12 (V2C_728_51),
	.V2C_13 (V2C_907_51),
	.V2C_14 (V2C_951_51),
	.V2C_15 (V2C_976_51),
	.V2C_16 (V2C_1036_51),
	.V2C_17 (V2C_1066_51),
	.V2C_18 (V2C_1111_51),
	.V2C_19 (V2C_1202_51),
	.V2C_20 (V2C_1203_51),
	.C2V_1 (C2V_51_17),
	.C2V_2 (C2V_51_92),
	.C2V_3 (C2V_51_109),
	.C2V_4 (C2V_51_191),
	.C2V_5 (C2V_51_209),
	.C2V_6 (C2V_51_276),
	.C2V_7 (C2V_51_373),
	.C2V_8 (C2V_51_428),
	.C2V_9 (C2V_51_539),
	.C2V_10 (C2V_51_596),
	.C2V_11 (C2V_51_672),
	.C2V_12 (C2V_51_728),
	.C2V_13 (C2V_51_907),
	.C2V_14 (C2V_51_951),
	.C2V_15 (C2V_51_976),
	.C2V_16 (C2V_51_1036),
	.C2V_17 (C2V_51_1066),
	.C2V_18 (C2V_51_1111),
	.C2V_19 (C2V_51_1202),
	.C2V_20 (C2V_51_1203),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU52 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_36_52),
	.V2C_2 (V2C_95_52),
	.V2C_3 (V2C_134_52),
	.V2C_4 (V2C_190_52),
	.V2C_5 (V2C_207_52),
	.V2C_6 (V2C_261_52),
	.V2C_7 (V2C_437_52),
	.V2C_8 (V2C_525_52),
	.V2C_9 (V2C_561_52),
	.V2C_10 (V2C_623_52),
	.V2C_11 (V2C_648_52),
	.V2C_12 (V2C_694_52),
	.V2C_13 (V2C_911_52),
	.V2C_14 (V2C_935_52),
	.V2C_15 (V2C_971_52),
	.V2C_16 (V2C_1049_52),
	.V2C_17 (V2C_1076_52),
	.V2C_18 (V2C_1140_52),
	.V2C_19 (V2C_1203_52),
	.V2C_20 (V2C_1204_52),
	.C2V_1 (C2V_52_36),
	.C2V_2 (C2V_52_95),
	.C2V_3 (C2V_52_134),
	.C2V_4 (C2V_52_190),
	.C2V_5 (C2V_52_207),
	.C2V_6 (C2V_52_261),
	.C2V_7 (C2V_52_437),
	.C2V_8 (C2V_52_525),
	.C2V_9 (C2V_52_561),
	.C2V_10 (C2V_52_623),
	.C2V_11 (C2V_52_648),
	.C2V_12 (C2V_52_694),
	.C2V_13 (C2V_52_911),
	.C2V_14 (C2V_52_935),
	.C2V_15 (C2V_52_971),
	.C2V_16 (C2V_52_1049),
	.C2V_17 (C2V_52_1076),
	.C2V_18 (C2V_52_1140),
	.C2V_19 (C2V_52_1203),
	.C2V_20 (C2V_52_1204),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU53 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_7_53),
	.V2C_2 (V2C_65_53),
	.V2C_3 (V2C_100_53),
	.V2C_4 (V2C_171_53),
	.V2C_5 (V2C_235_53),
	.V2C_6 (V2C_253_53),
	.V2C_7 (V2C_302_53),
	.V2C_8 (V2C_369_53),
	.V2C_9 (V2C_448_53),
	.V2C_10 (V2C_682_53),
	.V2C_11 (V2C_746_53),
	.V2C_12 (V2C_800_53),
	.V2C_13 (V2C_878_53),
	.V2C_14 (V2C_926_53),
	.V2C_15 (V2C_969_53),
	.V2C_16 (V2C_1021_53),
	.V2C_17 (V2C_1070_53),
	.V2C_18 (V2C_1118_53),
	.V2C_19 (V2C_1204_53),
	.V2C_20 (V2C_1205_53),
	.C2V_1 (C2V_53_7),
	.C2V_2 (C2V_53_65),
	.C2V_3 (C2V_53_100),
	.C2V_4 (C2V_53_171),
	.C2V_5 (C2V_53_235),
	.C2V_6 (C2V_53_253),
	.C2V_7 (C2V_53_302),
	.C2V_8 (C2V_53_369),
	.C2V_9 (C2V_53_448),
	.C2V_10 (C2V_53_682),
	.C2V_11 (C2V_53_746),
	.C2V_12 (C2V_53_800),
	.C2V_13 (C2V_53_878),
	.C2V_14 (C2V_53_926),
	.C2V_15 (C2V_53_969),
	.C2V_16 (C2V_53_1021),
	.C2V_17 (C2V_53_1070),
	.C2V_18 (C2V_53_1118),
	.C2V_19 (C2V_53_1204),
	.C2V_20 (C2V_53_1205),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU54 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_38_54),
	.V2C_2 (V2C_62_54),
	.V2C_3 (V2C_102_54),
	.V2C_4 (V2C_170_54),
	.V2C_5 (V2C_204_54),
	.V2C_6 (V2C_283_54),
	.V2C_7 (V2C_336_54),
	.V2C_8 (V2C_440_54),
	.V2C_9 (V2C_537_54),
	.V2C_10 (V2C_618_54),
	.V2C_11 (V2C_774_54),
	.V2C_12 (V2C_850_54),
	.V2C_13 (V2C_883_54),
	.V2C_14 (V2C_945_54),
	.V2C_15 (V2C_980_54),
	.V2C_16 (V2C_1047_54),
	.V2C_17 (V2C_1063_54),
	.V2C_18 (V2C_1113_54),
	.V2C_19 (V2C_1205_54),
	.V2C_20 (V2C_1206_54),
	.C2V_1 (C2V_54_38),
	.C2V_2 (C2V_54_62),
	.C2V_3 (C2V_54_102),
	.C2V_4 (C2V_54_170),
	.C2V_5 (C2V_54_204),
	.C2V_6 (C2V_54_283),
	.C2V_7 (C2V_54_336),
	.C2V_8 (C2V_54_440),
	.C2V_9 (C2V_54_537),
	.C2V_10 (C2V_54_618),
	.C2V_11 (C2V_54_774),
	.C2V_12 (C2V_54_850),
	.C2V_13 (C2V_54_883),
	.C2V_14 (C2V_54_945),
	.C2V_15 (C2V_54_980),
	.C2V_16 (C2V_54_1047),
	.C2V_17 (C2V_54_1063),
	.C2V_18 (C2V_54_1113),
	.C2V_19 (C2V_54_1205),
	.C2V_20 (C2V_54_1206),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU55 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_14_55),
	.V2C_2 (V2C_50_55),
	.V2C_3 (V2C_118_55),
	.V2C_4 (V2C_179_55),
	.V2C_5 (V2C_193_55),
	.V2C_6 (V2C_284_55),
	.V2C_7 (V2C_384_55),
	.V2C_8 (V2C_390_55),
	.V2C_9 (V2C_487_55),
	.V2C_10 (V2C_723_55),
	.V2C_11 (V2C_771_55),
	.V2C_12 (V2C_819_55),
	.V2C_13 (V2C_908_55),
	.V2C_14 (V2C_949_55),
	.V2C_15 (V2C_983_55),
	.V2C_16 (V2C_1022_55),
	.V2C_17 (V2C_1096_55),
	.V2C_18 (V2C_1107_55),
	.V2C_19 (V2C_1206_55),
	.V2C_20 (V2C_1207_55),
	.C2V_1 (C2V_55_14),
	.C2V_2 (C2V_55_50),
	.C2V_3 (C2V_55_118),
	.C2V_4 (C2V_55_179),
	.C2V_5 (C2V_55_193),
	.C2V_6 (C2V_55_284),
	.C2V_7 (C2V_55_384),
	.C2V_8 (C2V_55_390),
	.C2V_9 (C2V_55_487),
	.C2V_10 (C2V_55_723),
	.C2V_11 (C2V_55_771),
	.C2V_12 (C2V_55_819),
	.C2V_13 (C2V_55_908),
	.C2V_14 (C2V_55_949),
	.C2V_15 (C2V_55_983),
	.C2V_16 (C2V_55_1022),
	.C2V_17 (C2V_55_1096),
	.C2V_18 (C2V_55_1107),
	.C2V_19 (C2V_55_1206),
	.C2V_20 (C2V_55_1207),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU56 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_23_56),
	.V2C_2 (V2C_72_56),
	.V2C_3 (V2C_128_56),
	.V2C_4 (V2C_176_56),
	.V2C_5 (V2C_205_56),
	.V2C_6 (V2C_274_56),
	.V2C_7 (V2C_325_56),
	.V2C_8 (V2C_432_56),
	.V2C_9 (V2C_521_56),
	.V2C_10 (V2C_633_56),
	.V2C_11 (V2C_694_56),
	.V2C_12 (V2C_862_56),
	.V2C_13 (V2C_904_56),
	.V2C_14 (V2C_919_56),
	.V2C_15 (V2C_998_56),
	.V2C_16 (V2C_1030_56),
	.V2C_17 (V2C_1097_56),
	.V2C_18 (V2C_1128_56),
	.V2C_19 (V2C_1207_56),
	.V2C_20 (V2C_1208_56),
	.C2V_1 (C2V_56_23),
	.C2V_2 (C2V_56_72),
	.C2V_3 (C2V_56_128),
	.C2V_4 (C2V_56_176),
	.C2V_5 (C2V_56_205),
	.C2V_6 (C2V_56_274),
	.C2V_7 (C2V_56_325),
	.C2V_8 (C2V_56_432),
	.C2V_9 (C2V_56_521),
	.C2V_10 (C2V_56_633),
	.C2V_11 (C2V_56_694),
	.C2V_12 (C2V_56_862),
	.C2V_13 (C2V_56_904),
	.C2V_14 (C2V_56_919),
	.C2V_15 (C2V_56_998),
	.C2V_16 (C2V_56_1030),
	.C2V_17 (C2V_56_1097),
	.C2V_18 (C2V_56_1128),
	.C2V_19 (C2V_56_1207),
	.C2V_20 (C2V_56_1208),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU57 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_18_57),
	.V2C_2 (V2C_93_57),
	.V2C_3 (V2C_110_57),
	.V2C_4 (V2C_192_57),
	.V2C_5 (V2C_210_57),
	.V2C_6 (V2C_277_57),
	.V2C_7 (V2C_374_57),
	.V2C_8 (V2C_429_57),
	.V2C_9 (V2C_540_57),
	.V2C_10 (V2C_597_57),
	.V2C_11 (V2C_625_57),
	.V2C_12 (V2C_729_57),
	.V2C_13 (V2C_908_57),
	.V2C_14 (V2C_952_57),
	.V2C_15 (V2C_977_57),
	.V2C_16 (V2C_1037_57),
	.V2C_17 (V2C_1067_57),
	.V2C_18 (V2C_1112_57),
	.V2C_19 (V2C_1208_57),
	.V2C_20 (V2C_1209_57),
	.C2V_1 (C2V_57_18),
	.C2V_2 (C2V_57_93),
	.C2V_3 (C2V_57_110),
	.C2V_4 (C2V_57_192),
	.C2V_5 (C2V_57_210),
	.C2V_6 (C2V_57_277),
	.C2V_7 (C2V_57_374),
	.C2V_8 (C2V_57_429),
	.C2V_9 (C2V_57_540),
	.C2V_10 (C2V_57_597),
	.C2V_11 (C2V_57_625),
	.C2V_12 (C2V_57_729),
	.C2V_13 (C2V_57_908),
	.C2V_14 (C2V_57_952),
	.C2V_15 (C2V_57_977),
	.C2V_16 (C2V_57_1037),
	.C2V_17 (C2V_57_1067),
	.C2V_18 (C2V_57_1112),
	.C2V_19 (C2V_57_1208),
	.C2V_20 (C2V_57_1209),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU58 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_37_58),
	.V2C_2 (V2C_96_58),
	.V2C_3 (V2C_135_58),
	.V2C_4 (V2C_191_58),
	.V2C_5 (V2C_208_58),
	.V2C_6 (V2C_262_58),
	.V2C_7 (V2C_438_58),
	.V2C_8 (V2C_526_58),
	.V2C_9 (V2C_562_58),
	.V2C_10 (V2C_624_58),
	.V2C_11 (V2C_649_58),
	.V2C_12 (V2C_695_58),
	.V2C_13 (V2C_912_58),
	.V2C_14 (V2C_936_58),
	.V2C_15 (V2C_972_58),
	.V2C_16 (V2C_1050_58),
	.V2C_17 (V2C_1077_58),
	.V2C_18 (V2C_1141_58),
	.V2C_19 (V2C_1209_58),
	.V2C_20 (V2C_1210_58),
	.C2V_1 (C2V_58_37),
	.C2V_2 (C2V_58_96),
	.C2V_3 (C2V_58_135),
	.C2V_4 (C2V_58_191),
	.C2V_5 (C2V_58_208),
	.C2V_6 (C2V_58_262),
	.C2V_7 (C2V_58_438),
	.C2V_8 (C2V_58_526),
	.C2V_9 (C2V_58_562),
	.C2V_10 (C2V_58_624),
	.C2V_11 (C2V_58_649),
	.C2V_12 (C2V_58_695),
	.C2V_13 (C2V_58_912),
	.C2V_14 (C2V_58_936),
	.C2V_15 (C2V_58_972),
	.C2V_16 (C2V_58_1050),
	.C2V_17 (C2V_58_1077),
	.C2V_18 (C2V_58_1141),
	.C2V_19 (C2V_58_1209),
	.C2V_20 (C2V_58_1210),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU59 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_8_59),
	.V2C_2 (V2C_66_59),
	.V2C_3 (V2C_101_59),
	.V2C_4 (V2C_172_59),
	.V2C_5 (V2C_236_59),
	.V2C_6 (V2C_254_59),
	.V2C_7 (V2C_303_59),
	.V2C_8 (V2C_370_59),
	.V2C_9 (V2C_449_59),
	.V2C_10 (V2C_683_59),
	.V2C_11 (V2C_747_59),
	.V2C_12 (V2C_801_59),
	.V2C_13 (V2C_879_59),
	.V2C_14 (V2C_927_59),
	.V2C_15 (V2C_970_59),
	.V2C_16 (V2C_1022_59),
	.V2C_17 (V2C_1071_59),
	.V2C_18 (V2C_1119_59),
	.V2C_19 (V2C_1210_59),
	.V2C_20 (V2C_1211_59),
	.C2V_1 (C2V_59_8),
	.C2V_2 (C2V_59_66),
	.C2V_3 (C2V_59_101),
	.C2V_4 (C2V_59_172),
	.C2V_5 (C2V_59_236),
	.C2V_6 (C2V_59_254),
	.C2V_7 (C2V_59_303),
	.C2V_8 (C2V_59_370),
	.C2V_9 (C2V_59_449),
	.C2V_10 (C2V_59_683),
	.C2V_11 (C2V_59_747),
	.C2V_12 (C2V_59_801),
	.C2V_13 (C2V_59_879),
	.C2V_14 (C2V_59_927),
	.C2V_15 (C2V_59_970),
	.C2V_16 (C2V_59_1022),
	.C2V_17 (C2V_59_1071),
	.C2V_18 (C2V_59_1119),
	.C2V_19 (C2V_59_1210),
	.C2V_20 (C2V_59_1211),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU60 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_39_60),
	.V2C_2 (V2C_63_60),
	.V2C_3 (V2C_103_60),
	.V2C_4 (V2C_171_60),
	.V2C_5 (V2C_205_60),
	.V2C_6 (V2C_284_60),
	.V2C_7 (V2C_289_60),
	.V2C_8 (V2C_441_60),
	.V2C_9 (V2C_538_60),
	.V2C_10 (V2C_619_60),
	.V2C_11 (V2C_775_60),
	.V2C_12 (V2C_851_60),
	.V2C_13 (V2C_884_60),
	.V2C_14 (V2C_946_60),
	.V2C_15 (V2C_981_60),
	.V2C_16 (V2C_1048_60),
	.V2C_17 (V2C_1064_60),
	.V2C_18 (V2C_1114_60),
	.V2C_19 (V2C_1211_60),
	.V2C_20 (V2C_1212_60),
	.C2V_1 (C2V_60_39),
	.C2V_2 (C2V_60_63),
	.C2V_3 (C2V_60_103),
	.C2V_4 (C2V_60_171),
	.C2V_5 (C2V_60_205),
	.C2V_6 (C2V_60_284),
	.C2V_7 (C2V_60_289),
	.C2V_8 (C2V_60_441),
	.C2V_9 (C2V_60_538),
	.C2V_10 (C2V_60_619),
	.C2V_11 (C2V_60_775),
	.C2V_12 (C2V_60_851),
	.C2V_13 (C2V_60_884),
	.C2V_14 (C2V_60_946),
	.C2V_15 (C2V_60_981),
	.C2V_16 (C2V_60_1048),
	.C2V_17 (C2V_60_1064),
	.C2V_18 (C2V_60_1114),
	.C2V_19 (C2V_60_1211),
	.C2V_20 (C2V_60_1212),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU61 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_15_61),
	.V2C_2 (V2C_51_61),
	.V2C_3 (V2C_119_61),
	.V2C_4 (V2C_180_61),
	.V2C_5 (V2C_194_61),
	.V2C_6 (V2C_285_61),
	.V2C_7 (V2C_337_61),
	.V2C_8 (V2C_391_61),
	.V2C_9 (V2C_488_61),
	.V2C_10 (V2C_724_61),
	.V2C_11 (V2C_772_61),
	.V2C_12 (V2C_820_61),
	.V2C_13 (V2C_909_61),
	.V2C_14 (V2C_950_61),
	.V2C_15 (V2C_984_61),
	.V2C_16 (V2C_1023_61),
	.V2C_17 (V2C_1097_61),
	.V2C_18 (V2C_1108_61),
	.V2C_19 (V2C_1212_61),
	.V2C_20 (V2C_1213_61),
	.C2V_1 (C2V_61_15),
	.C2V_2 (C2V_61_51),
	.C2V_3 (C2V_61_119),
	.C2V_4 (C2V_61_180),
	.C2V_5 (C2V_61_194),
	.C2V_6 (C2V_61_285),
	.C2V_7 (C2V_61_337),
	.C2V_8 (C2V_61_391),
	.C2V_9 (C2V_61_488),
	.C2V_10 (C2V_61_724),
	.C2V_11 (C2V_61_772),
	.C2V_12 (C2V_61_820),
	.C2V_13 (C2V_61_909),
	.C2V_14 (C2V_61_950),
	.C2V_15 (C2V_61_984),
	.C2V_16 (C2V_61_1023),
	.C2V_17 (C2V_61_1097),
	.C2V_18 (C2V_61_1108),
	.C2V_19 (C2V_61_1212),
	.C2V_20 (C2V_61_1213),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU62 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_24_62),
	.V2C_2 (V2C_73_62),
	.V2C_3 (V2C_129_62),
	.V2C_4 (V2C_177_62),
	.V2C_5 (V2C_206_62),
	.V2C_6 (V2C_275_62),
	.V2C_7 (V2C_326_62),
	.V2C_8 (V2C_385_62),
	.V2C_9 (V2C_522_62),
	.V2C_10 (V2C_634_62),
	.V2C_11 (V2C_695_62),
	.V2C_12 (V2C_863_62),
	.V2C_13 (V2C_905_62),
	.V2C_14 (V2C_920_62),
	.V2C_15 (V2C_999_62),
	.V2C_16 (V2C_1031_62),
	.V2C_17 (V2C_1098_62),
	.V2C_18 (V2C_1129_62),
	.V2C_19 (V2C_1213_62),
	.V2C_20 (V2C_1214_62),
	.C2V_1 (C2V_62_24),
	.C2V_2 (C2V_62_73),
	.C2V_3 (C2V_62_129),
	.C2V_4 (C2V_62_177),
	.C2V_5 (C2V_62_206),
	.C2V_6 (C2V_62_275),
	.C2V_7 (C2V_62_326),
	.C2V_8 (C2V_62_385),
	.C2V_9 (C2V_62_522),
	.C2V_10 (C2V_62_634),
	.C2V_11 (C2V_62_695),
	.C2V_12 (C2V_62_863),
	.C2V_13 (C2V_62_905),
	.C2V_14 (C2V_62_920),
	.C2V_15 (C2V_62_999),
	.C2V_16 (C2V_62_1031),
	.C2V_17 (C2V_62_1098),
	.C2V_18 (C2V_62_1129),
	.C2V_19 (C2V_62_1213),
	.C2V_20 (C2V_62_1214),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU63 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_19_63),
	.V2C_2 (V2C_94_63),
	.V2C_3 (V2C_111_63),
	.V2C_4 (V2C_145_63),
	.V2C_5 (V2C_211_63),
	.V2C_6 (V2C_278_63),
	.V2C_7 (V2C_375_63),
	.V2C_8 (V2C_430_63),
	.V2C_9 (V2C_541_63),
	.V2C_10 (V2C_598_63),
	.V2C_11 (V2C_626_63),
	.V2C_12 (V2C_730_63),
	.V2C_13 (V2C_909_63),
	.V2C_14 (V2C_953_63),
	.V2C_15 (V2C_978_63),
	.V2C_16 (V2C_1038_63),
	.V2C_17 (V2C_1068_63),
	.V2C_18 (V2C_1113_63),
	.V2C_19 (V2C_1214_63),
	.V2C_20 (V2C_1215_63),
	.C2V_1 (C2V_63_19),
	.C2V_2 (C2V_63_94),
	.C2V_3 (C2V_63_111),
	.C2V_4 (C2V_63_145),
	.C2V_5 (C2V_63_211),
	.C2V_6 (C2V_63_278),
	.C2V_7 (C2V_63_375),
	.C2V_8 (C2V_63_430),
	.C2V_9 (C2V_63_541),
	.C2V_10 (C2V_63_598),
	.C2V_11 (C2V_63_626),
	.C2V_12 (C2V_63_730),
	.C2V_13 (C2V_63_909),
	.C2V_14 (C2V_63_953),
	.C2V_15 (C2V_63_978),
	.C2V_16 (C2V_63_1038),
	.C2V_17 (C2V_63_1068),
	.C2V_18 (C2V_63_1113),
	.C2V_19 (C2V_63_1214),
	.C2V_20 (C2V_63_1215),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU64 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_38_64),
	.V2C_2 (V2C_49_64),
	.V2C_3 (V2C_136_64),
	.V2C_4 (V2C_192_64),
	.V2C_5 (V2C_209_64),
	.V2C_6 (V2C_263_64),
	.V2C_7 (V2C_439_64),
	.V2C_8 (V2C_527_64),
	.V2C_9 (V2C_563_64),
	.V2C_10 (V2C_577_64),
	.V2C_11 (V2C_650_64),
	.V2C_12 (V2C_696_64),
	.V2C_13 (V2C_865_64),
	.V2C_14 (V2C_937_64),
	.V2C_15 (V2C_973_64),
	.V2C_16 (V2C_1051_64),
	.V2C_17 (V2C_1078_64),
	.V2C_18 (V2C_1142_64),
	.V2C_19 (V2C_1215_64),
	.V2C_20 (V2C_1216_64),
	.C2V_1 (C2V_64_38),
	.C2V_2 (C2V_64_49),
	.C2V_3 (C2V_64_136),
	.C2V_4 (C2V_64_192),
	.C2V_5 (C2V_64_209),
	.C2V_6 (C2V_64_263),
	.C2V_7 (C2V_64_439),
	.C2V_8 (C2V_64_527),
	.C2V_9 (C2V_64_563),
	.C2V_10 (C2V_64_577),
	.C2V_11 (C2V_64_650),
	.C2V_12 (C2V_64_696),
	.C2V_13 (C2V_64_865),
	.C2V_14 (C2V_64_937),
	.C2V_15 (C2V_64_973),
	.C2V_16 (C2V_64_1051),
	.C2V_17 (C2V_64_1078),
	.C2V_18 (C2V_64_1142),
	.C2V_19 (C2V_64_1215),
	.C2V_20 (C2V_64_1216),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU65 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_9_65),
	.V2C_2 (V2C_67_65),
	.V2C_3 (V2C_102_65),
	.V2C_4 (V2C_173_65),
	.V2C_5 (V2C_237_65),
	.V2C_6 (V2C_255_65),
	.V2C_7 (V2C_304_65),
	.V2C_8 (V2C_371_65),
	.V2C_9 (V2C_450_65),
	.V2C_10 (V2C_684_65),
	.V2C_11 (V2C_748_65),
	.V2C_12 (V2C_802_65),
	.V2C_13 (V2C_880_65),
	.V2C_14 (V2C_928_65),
	.V2C_15 (V2C_971_65),
	.V2C_16 (V2C_1023_65),
	.V2C_17 (V2C_1072_65),
	.V2C_18 (V2C_1120_65),
	.V2C_19 (V2C_1216_65),
	.V2C_20 (V2C_1217_65),
	.C2V_1 (C2V_65_9),
	.C2V_2 (C2V_65_67),
	.C2V_3 (C2V_65_102),
	.C2V_4 (C2V_65_173),
	.C2V_5 (C2V_65_237),
	.C2V_6 (C2V_65_255),
	.C2V_7 (C2V_65_304),
	.C2V_8 (C2V_65_371),
	.C2V_9 (C2V_65_450),
	.C2V_10 (C2V_65_684),
	.C2V_11 (C2V_65_748),
	.C2V_12 (C2V_65_802),
	.C2V_13 (C2V_65_880),
	.C2V_14 (C2V_65_928),
	.C2V_15 (C2V_65_971),
	.C2V_16 (C2V_65_1023),
	.C2V_17 (C2V_65_1072),
	.C2V_18 (C2V_65_1120),
	.C2V_19 (C2V_65_1216),
	.C2V_20 (C2V_65_1217),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU66 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_40_66),
	.V2C_2 (V2C_64_66),
	.V2C_3 (V2C_104_66),
	.V2C_4 (V2C_172_66),
	.V2C_5 (V2C_206_66),
	.V2C_6 (V2C_285_66),
	.V2C_7 (V2C_290_66),
	.V2C_8 (V2C_442_66),
	.V2C_9 (V2C_539_66),
	.V2C_10 (V2C_620_66),
	.V2C_11 (V2C_776_66),
	.V2C_12 (V2C_852_66),
	.V2C_13 (V2C_885_66),
	.V2C_14 (V2C_947_66),
	.V2C_15 (V2C_982_66),
	.V2C_16 (V2C_1049_66),
	.V2C_17 (V2C_1065_66),
	.V2C_18 (V2C_1115_66),
	.V2C_19 (V2C_1217_66),
	.V2C_20 (V2C_1218_66),
	.C2V_1 (C2V_66_40),
	.C2V_2 (C2V_66_64),
	.C2V_3 (C2V_66_104),
	.C2V_4 (C2V_66_172),
	.C2V_5 (C2V_66_206),
	.C2V_6 (C2V_66_285),
	.C2V_7 (C2V_66_290),
	.C2V_8 (C2V_66_442),
	.C2V_9 (C2V_66_539),
	.C2V_10 (C2V_66_620),
	.C2V_11 (C2V_66_776),
	.C2V_12 (C2V_66_852),
	.C2V_13 (C2V_66_885),
	.C2V_14 (C2V_66_947),
	.C2V_15 (C2V_66_982),
	.C2V_16 (C2V_66_1049),
	.C2V_17 (C2V_66_1065),
	.C2V_18 (C2V_66_1115),
	.C2V_19 (C2V_66_1217),
	.C2V_20 (C2V_66_1218),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU67 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_16_67),
	.V2C_2 (V2C_52_67),
	.V2C_3 (V2C_120_67),
	.V2C_4 (V2C_181_67),
	.V2C_5 (V2C_195_67),
	.V2C_6 (V2C_286_67),
	.V2C_7 (V2C_338_67),
	.V2C_8 (V2C_392_67),
	.V2C_9 (V2C_489_67),
	.V2C_10 (V2C_725_67),
	.V2C_11 (V2C_773_67),
	.V2C_12 (V2C_821_67),
	.V2C_13 (V2C_910_67),
	.V2C_14 (V2C_951_67),
	.V2C_15 (V2C_985_67),
	.V2C_16 (V2C_1024_67),
	.V2C_17 (V2C_1098_67),
	.V2C_18 (V2C_1109_67),
	.V2C_19 (V2C_1218_67),
	.V2C_20 (V2C_1219_67),
	.C2V_1 (C2V_67_16),
	.C2V_2 (C2V_67_52),
	.C2V_3 (C2V_67_120),
	.C2V_4 (C2V_67_181),
	.C2V_5 (C2V_67_195),
	.C2V_6 (C2V_67_286),
	.C2V_7 (C2V_67_338),
	.C2V_8 (C2V_67_392),
	.C2V_9 (C2V_67_489),
	.C2V_10 (C2V_67_725),
	.C2V_11 (C2V_67_773),
	.C2V_12 (C2V_67_821),
	.C2V_13 (C2V_67_910),
	.C2V_14 (C2V_67_951),
	.C2V_15 (C2V_67_985),
	.C2V_16 (C2V_67_1024),
	.C2V_17 (C2V_67_1098),
	.C2V_18 (C2V_67_1109),
	.C2V_19 (C2V_67_1218),
	.C2V_20 (C2V_67_1219),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU68 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_25_68),
	.V2C_2 (V2C_74_68),
	.V2C_3 (V2C_130_68),
	.V2C_4 (V2C_178_68),
	.V2C_5 (V2C_207_68),
	.V2C_6 (V2C_276_68),
	.V2C_7 (V2C_327_68),
	.V2C_8 (V2C_386_68),
	.V2C_9 (V2C_523_68),
	.V2C_10 (V2C_635_68),
	.V2C_11 (V2C_696_68),
	.V2C_12 (V2C_864_68),
	.V2C_13 (V2C_906_68),
	.V2C_14 (V2C_921_68),
	.V2C_15 (V2C_1000_68),
	.V2C_16 (V2C_1032_68),
	.V2C_17 (V2C_1099_68),
	.V2C_18 (V2C_1130_68),
	.V2C_19 (V2C_1219_68),
	.V2C_20 (V2C_1220_68),
	.C2V_1 (C2V_68_25),
	.C2V_2 (C2V_68_74),
	.C2V_3 (C2V_68_130),
	.C2V_4 (C2V_68_178),
	.C2V_5 (C2V_68_207),
	.C2V_6 (C2V_68_276),
	.C2V_7 (C2V_68_327),
	.C2V_8 (C2V_68_386),
	.C2V_9 (C2V_68_523),
	.C2V_10 (C2V_68_635),
	.C2V_11 (C2V_68_696),
	.C2V_12 (C2V_68_864),
	.C2V_13 (C2V_68_906),
	.C2V_14 (C2V_68_921),
	.C2V_15 (C2V_68_1000),
	.C2V_16 (C2V_68_1032),
	.C2V_17 (C2V_68_1099),
	.C2V_18 (C2V_68_1130),
	.C2V_19 (C2V_68_1219),
	.C2V_20 (C2V_68_1220),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU69 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_20_69),
	.V2C_2 (V2C_95_69),
	.V2C_3 (V2C_112_69),
	.V2C_4 (V2C_146_69),
	.V2C_5 (V2C_212_69),
	.V2C_6 (V2C_279_69),
	.V2C_7 (V2C_376_69),
	.V2C_8 (V2C_431_69),
	.V2C_9 (V2C_542_69),
	.V2C_10 (V2C_599_69),
	.V2C_11 (V2C_627_69),
	.V2C_12 (V2C_731_69),
	.V2C_13 (V2C_910_69),
	.V2C_14 (V2C_954_69),
	.V2C_15 (V2C_979_69),
	.V2C_16 (V2C_1039_69),
	.V2C_17 (V2C_1069_69),
	.V2C_18 (V2C_1114_69),
	.V2C_19 (V2C_1220_69),
	.V2C_20 (V2C_1221_69),
	.C2V_1 (C2V_69_20),
	.C2V_2 (C2V_69_95),
	.C2V_3 (C2V_69_112),
	.C2V_4 (C2V_69_146),
	.C2V_5 (C2V_69_212),
	.C2V_6 (C2V_69_279),
	.C2V_7 (C2V_69_376),
	.C2V_8 (C2V_69_431),
	.C2V_9 (C2V_69_542),
	.C2V_10 (C2V_69_599),
	.C2V_11 (C2V_69_627),
	.C2V_12 (C2V_69_731),
	.C2V_13 (C2V_69_910),
	.C2V_14 (C2V_69_954),
	.C2V_15 (C2V_69_979),
	.C2V_16 (C2V_69_1039),
	.C2V_17 (C2V_69_1069),
	.C2V_18 (C2V_69_1114),
	.C2V_19 (C2V_69_1220),
	.C2V_20 (C2V_69_1221),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU70 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_39_70),
	.V2C_2 (V2C_50_70),
	.V2C_3 (V2C_137_70),
	.V2C_4 (V2C_145_70),
	.V2C_5 (V2C_210_70),
	.V2C_6 (V2C_264_70),
	.V2C_7 (V2C_440_70),
	.V2C_8 (V2C_528_70),
	.V2C_9 (V2C_564_70),
	.V2C_10 (V2C_578_70),
	.V2C_11 (V2C_651_70),
	.V2C_12 (V2C_697_70),
	.V2C_13 (V2C_866_70),
	.V2C_14 (V2C_938_70),
	.V2C_15 (V2C_974_70),
	.V2C_16 (V2C_1052_70),
	.V2C_17 (V2C_1079_70),
	.V2C_18 (V2C_1143_70),
	.V2C_19 (V2C_1221_70),
	.V2C_20 (V2C_1222_70),
	.C2V_1 (C2V_70_39),
	.C2V_2 (C2V_70_50),
	.C2V_3 (C2V_70_137),
	.C2V_4 (C2V_70_145),
	.C2V_5 (C2V_70_210),
	.C2V_6 (C2V_70_264),
	.C2V_7 (C2V_70_440),
	.C2V_8 (C2V_70_528),
	.C2V_9 (C2V_70_564),
	.C2V_10 (C2V_70_578),
	.C2V_11 (C2V_70_651),
	.C2V_12 (C2V_70_697),
	.C2V_13 (C2V_70_866),
	.C2V_14 (C2V_70_938),
	.C2V_15 (C2V_70_974),
	.C2V_16 (C2V_70_1052),
	.C2V_17 (C2V_70_1079),
	.C2V_18 (C2V_70_1143),
	.C2V_19 (C2V_70_1221),
	.C2V_20 (C2V_70_1222),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU71 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_10_71),
	.V2C_2 (V2C_68_71),
	.V2C_3 (V2C_103_71),
	.V2C_4 (V2C_174_71),
	.V2C_5 (V2C_238_71),
	.V2C_6 (V2C_256_71),
	.V2C_7 (V2C_305_71),
	.V2C_8 (V2C_372_71),
	.V2C_9 (V2C_451_71),
	.V2C_10 (V2C_685_71),
	.V2C_11 (V2C_749_71),
	.V2C_12 (V2C_803_71),
	.V2C_13 (V2C_881_71),
	.V2C_14 (V2C_929_71),
	.V2C_15 (V2C_972_71),
	.V2C_16 (V2C_1024_71),
	.V2C_17 (V2C_1073_71),
	.V2C_18 (V2C_1121_71),
	.V2C_19 (V2C_1222_71),
	.V2C_20 (V2C_1223_71),
	.C2V_1 (C2V_71_10),
	.C2V_2 (C2V_71_68),
	.C2V_3 (C2V_71_103),
	.C2V_4 (C2V_71_174),
	.C2V_5 (C2V_71_238),
	.C2V_6 (C2V_71_256),
	.C2V_7 (C2V_71_305),
	.C2V_8 (C2V_71_372),
	.C2V_9 (C2V_71_451),
	.C2V_10 (C2V_71_685),
	.C2V_11 (C2V_71_749),
	.C2V_12 (C2V_71_803),
	.C2V_13 (C2V_71_881),
	.C2V_14 (C2V_71_929),
	.C2V_15 (C2V_71_972),
	.C2V_16 (C2V_71_1024),
	.C2V_17 (C2V_71_1073),
	.C2V_18 (C2V_71_1121),
	.C2V_19 (C2V_71_1222),
	.C2V_20 (C2V_71_1223),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU72 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_41_72),
	.V2C_2 (V2C_65_72),
	.V2C_3 (V2C_105_72),
	.V2C_4 (V2C_173_72),
	.V2C_5 (V2C_207_72),
	.V2C_6 (V2C_286_72),
	.V2C_7 (V2C_291_72),
	.V2C_8 (V2C_443_72),
	.V2C_9 (V2C_540_72),
	.V2C_10 (V2C_621_72),
	.V2C_11 (V2C_777_72),
	.V2C_12 (V2C_853_72),
	.V2C_13 (V2C_886_72),
	.V2C_14 (V2C_948_72),
	.V2C_15 (V2C_983_72),
	.V2C_16 (V2C_1050_72),
	.V2C_17 (V2C_1066_72),
	.V2C_18 (V2C_1116_72),
	.V2C_19 (V2C_1223_72),
	.V2C_20 (V2C_1224_72),
	.C2V_1 (C2V_72_41),
	.C2V_2 (C2V_72_65),
	.C2V_3 (C2V_72_105),
	.C2V_4 (C2V_72_173),
	.C2V_5 (C2V_72_207),
	.C2V_6 (C2V_72_286),
	.C2V_7 (C2V_72_291),
	.C2V_8 (C2V_72_443),
	.C2V_9 (C2V_72_540),
	.C2V_10 (C2V_72_621),
	.C2V_11 (C2V_72_777),
	.C2V_12 (C2V_72_853),
	.C2V_13 (C2V_72_886),
	.C2V_14 (C2V_72_948),
	.C2V_15 (C2V_72_983),
	.C2V_16 (C2V_72_1050),
	.C2V_17 (C2V_72_1066),
	.C2V_18 (C2V_72_1116),
	.C2V_19 (C2V_72_1223),
	.C2V_20 (C2V_72_1224),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU73 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_17_73),
	.V2C_2 (V2C_53_73),
	.V2C_3 (V2C_121_73),
	.V2C_4 (V2C_182_73),
	.V2C_5 (V2C_196_73),
	.V2C_6 (V2C_287_73),
	.V2C_7 (V2C_339_73),
	.V2C_8 (V2C_393_73),
	.V2C_9 (V2C_490_73),
	.V2C_10 (V2C_726_73),
	.V2C_11 (V2C_774_73),
	.V2C_12 (V2C_822_73),
	.V2C_13 (V2C_911_73),
	.V2C_14 (V2C_952_73),
	.V2C_15 (V2C_986_73),
	.V2C_16 (V2C_1025_73),
	.V2C_17 (V2C_1099_73),
	.V2C_18 (V2C_1110_73),
	.V2C_19 (V2C_1224_73),
	.V2C_20 (V2C_1225_73),
	.C2V_1 (C2V_73_17),
	.C2V_2 (C2V_73_53),
	.C2V_3 (C2V_73_121),
	.C2V_4 (C2V_73_182),
	.C2V_5 (C2V_73_196),
	.C2V_6 (C2V_73_287),
	.C2V_7 (C2V_73_339),
	.C2V_8 (C2V_73_393),
	.C2V_9 (C2V_73_490),
	.C2V_10 (C2V_73_726),
	.C2V_11 (C2V_73_774),
	.C2V_12 (C2V_73_822),
	.C2V_13 (C2V_73_911),
	.C2V_14 (C2V_73_952),
	.C2V_15 (C2V_73_986),
	.C2V_16 (C2V_73_1025),
	.C2V_17 (C2V_73_1099),
	.C2V_18 (C2V_73_1110),
	.C2V_19 (C2V_73_1224),
	.C2V_20 (C2V_73_1225),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU74 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_26_74),
	.V2C_2 (V2C_75_74),
	.V2C_3 (V2C_131_74),
	.V2C_4 (V2C_179_74),
	.V2C_5 (V2C_208_74),
	.V2C_6 (V2C_277_74),
	.V2C_7 (V2C_328_74),
	.V2C_8 (V2C_387_74),
	.V2C_9 (V2C_524_74),
	.V2C_10 (V2C_636_74),
	.V2C_11 (V2C_697_74),
	.V2C_12 (V2C_817_74),
	.V2C_13 (V2C_907_74),
	.V2C_14 (V2C_922_74),
	.V2C_15 (V2C_1001_74),
	.V2C_16 (V2C_1033_74),
	.V2C_17 (V2C_1100_74),
	.V2C_18 (V2C_1131_74),
	.V2C_19 (V2C_1225_74),
	.V2C_20 (V2C_1226_74),
	.C2V_1 (C2V_74_26),
	.C2V_2 (C2V_74_75),
	.C2V_3 (C2V_74_131),
	.C2V_4 (C2V_74_179),
	.C2V_5 (C2V_74_208),
	.C2V_6 (C2V_74_277),
	.C2V_7 (C2V_74_328),
	.C2V_8 (C2V_74_387),
	.C2V_9 (C2V_74_524),
	.C2V_10 (C2V_74_636),
	.C2V_11 (C2V_74_697),
	.C2V_12 (C2V_74_817),
	.C2V_13 (C2V_74_907),
	.C2V_14 (C2V_74_922),
	.C2V_15 (C2V_74_1001),
	.C2V_16 (C2V_74_1033),
	.C2V_17 (C2V_74_1100),
	.C2V_18 (C2V_74_1131),
	.C2V_19 (C2V_74_1225),
	.C2V_20 (C2V_74_1226),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU75 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_21_75),
	.V2C_2 (V2C_96_75),
	.V2C_3 (V2C_113_75),
	.V2C_4 (V2C_147_75),
	.V2C_5 (V2C_213_75),
	.V2C_6 (V2C_280_75),
	.V2C_7 (V2C_377_75),
	.V2C_8 (V2C_432_75),
	.V2C_9 (V2C_543_75),
	.V2C_10 (V2C_600_75),
	.V2C_11 (V2C_628_75),
	.V2C_12 (V2C_732_75),
	.V2C_13 (V2C_911_75),
	.V2C_14 (V2C_955_75),
	.V2C_15 (V2C_980_75),
	.V2C_16 (V2C_1040_75),
	.V2C_17 (V2C_1070_75),
	.V2C_18 (V2C_1115_75),
	.V2C_19 (V2C_1226_75),
	.V2C_20 (V2C_1227_75),
	.C2V_1 (C2V_75_21),
	.C2V_2 (C2V_75_96),
	.C2V_3 (C2V_75_113),
	.C2V_4 (C2V_75_147),
	.C2V_5 (C2V_75_213),
	.C2V_6 (C2V_75_280),
	.C2V_7 (C2V_75_377),
	.C2V_8 (C2V_75_432),
	.C2V_9 (C2V_75_543),
	.C2V_10 (C2V_75_600),
	.C2V_11 (C2V_75_628),
	.C2V_12 (C2V_75_732),
	.C2V_13 (C2V_75_911),
	.C2V_14 (C2V_75_955),
	.C2V_15 (C2V_75_980),
	.C2V_16 (C2V_75_1040),
	.C2V_17 (C2V_75_1070),
	.C2V_18 (C2V_75_1115),
	.C2V_19 (C2V_75_1226),
	.C2V_20 (C2V_75_1227),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU76 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_40_76),
	.V2C_2 (V2C_51_76),
	.V2C_3 (V2C_138_76),
	.V2C_4 (V2C_146_76),
	.V2C_5 (V2C_211_76),
	.V2C_6 (V2C_265_76),
	.V2C_7 (V2C_441_76),
	.V2C_8 (V2C_481_76),
	.V2C_9 (V2C_565_76),
	.V2C_10 (V2C_579_76),
	.V2C_11 (V2C_652_76),
	.V2C_12 (V2C_698_76),
	.V2C_13 (V2C_867_76),
	.V2C_14 (V2C_939_76),
	.V2C_15 (V2C_975_76),
	.V2C_16 (V2C_1053_76),
	.V2C_17 (V2C_1080_76),
	.V2C_18 (V2C_1144_76),
	.V2C_19 (V2C_1227_76),
	.V2C_20 (V2C_1228_76),
	.C2V_1 (C2V_76_40),
	.C2V_2 (C2V_76_51),
	.C2V_3 (C2V_76_138),
	.C2V_4 (C2V_76_146),
	.C2V_5 (C2V_76_211),
	.C2V_6 (C2V_76_265),
	.C2V_7 (C2V_76_441),
	.C2V_8 (C2V_76_481),
	.C2V_9 (C2V_76_565),
	.C2V_10 (C2V_76_579),
	.C2V_11 (C2V_76_652),
	.C2V_12 (C2V_76_698),
	.C2V_13 (C2V_76_867),
	.C2V_14 (C2V_76_939),
	.C2V_15 (C2V_76_975),
	.C2V_16 (C2V_76_1053),
	.C2V_17 (C2V_76_1080),
	.C2V_18 (C2V_76_1144),
	.C2V_19 (C2V_76_1227),
	.C2V_20 (C2V_76_1228),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU77 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_11_77),
	.V2C_2 (V2C_69_77),
	.V2C_3 (V2C_104_77),
	.V2C_4 (V2C_175_77),
	.V2C_5 (V2C_239_77),
	.V2C_6 (V2C_257_77),
	.V2C_7 (V2C_306_77),
	.V2C_8 (V2C_373_77),
	.V2C_9 (V2C_452_77),
	.V2C_10 (V2C_686_77),
	.V2C_11 (V2C_750_77),
	.V2C_12 (V2C_804_77),
	.V2C_13 (V2C_882_77),
	.V2C_14 (V2C_930_77),
	.V2C_15 (V2C_973_77),
	.V2C_16 (V2C_1025_77),
	.V2C_17 (V2C_1074_77),
	.V2C_18 (V2C_1122_77),
	.V2C_19 (V2C_1228_77),
	.V2C_20 (V2C_1229_77),
	.C2V_1 (C2V_77_11),
	.C2V_2 (C2V_77_69),
	.C2V_3 (C2V_77_104),
	.C2V_4 (C2V_77_175),
	.C2V_5 (C2V_77_239),
	.C2V_6 (C2V_77_257),
	.C2V_7 (C2V_77_306),
	.C2V_8 (C2V_77_373),
	.C2V_9 (C2V_77_452),
	.C2V_10 (C2V_77_686),
	.C2V_11 (C2V_77_750),
	.C2V_12 (C2V_77_804),
	.C2V_13 (C2V_77_882),
	.C2V_14 (C2V_77_930),
	.C2V_15 (C2V_77_973),
	.C2V_16 (C2V_77_1025),
	.C2V_17 (C2V_77_1074),
	.C2V_18 (C2V_77_1122),
	.C2V_19 (C2V_77_1228),
	.C2V_20 (C2V_77_1229),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU78 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_42_78),
	.V2C_2 (V2C_66_78),
	.V2C_3 (V2C_106_78),
	.V2C_4 (V2C_174_78),
	.V2C_5 (V2C_208_78),
	.V2C_6 (V2C_287_78),
	.V2C_7 (V2C_292_78),
	.V2C_8 (V2C_444_78),
	.V2C_9 (V2C_541_78),
	.V2C_10 (V2C_622_78),
	.V2C_11 (V2C_778_78),
	.V2C_12 (V2C_854_78),
	.V2C_13 (V2C_887_78),
	.V2C_14 (V2C_949_78),
	.V2C_15 (V2C_984_78),
	.V2C_16 (V2C_1051_78),
	.V2C_17 (V2C_1067_78),
	.V2C_18 (V2C_1117_78),
	.V2C_19 (V2C_1229_78),
	.V2C_20 (V2C_1230_78),
	.C2V_1 (C2V_78_42),
	.C2V_2 (C2V_78_66),
	.C2V_3 (C2V_78_106),
	.C2V_4 (C2V_78_174),
	.C2V_5 (C2V_78_208),
	.C2V_6 (C2V_78_287),
	.C2V_7 (C2V_78_292),
	.C2V_8 (C2V_78_444),
	.C2V_9 (C2V_78_541),
	.C2V_10 (C2V_78_622),
	.C2V_11 (C2V_78_778),
	.C2V_12 (C2V_78_854),
	.C2V_13 (C2V_78_887),
	.C2V_14 (C2V_78_949),
	.C2V_15 (C2V_78_984),
	.C2V_16 (C2V_78_1051),
	.C2V_17 (C2V_78_1067),
	.C2V_18 (C2V_78_1117),
	.C2V_19 (C2V_78_1229),
	.C2V_20 (C2V_78_1230),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU79 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_18_79),
	.V2C_2 (V2C_54_79),
	.V2C_3 (V2C_122_79),
	.V2C_4 (V2C_183_79),
	.V2C_5 (V2C_197_79),
	.V2C_6 (V2C_288_79),
	.V2C_7 (V2C_340_79),
	.V2C_8 (V2C_394_79),
	.V2C_9 (V2C_491_79),
	.V2C_10 (V2C_727_79),
	.V2C_11 (V2C_775_79),
	.V2C_12 (V2C_823_79),
	.V2C_13 (V2C_912_79),
	.V2C_14 (V2C_953_79),
	.V2C_15 (V2C_987_79),
	.V2C_16 (V2C_1026_79),
	.V2C_17 (V2C_1100_79),
	.V2C_18 (V2C_1111_79),
	.V2C_19 (V2C_1230_79),
	.V2C_20 (V2C_1231_79),
	.C2V_1 (C2V_79_18),
	.C2V_2 (C2V_79_54),
	.C2V_3 (C2V_79_122),
	.C2V_4 (C2V_79_183),
	.C2V_5 (C2V_79_197),
	.C2V_6 (C2V_79_288),
	.C2V_7 (C2V_79_340),
	.C2V_8 (C2V_79_394),
	.C2V_9 (C2V_79_491),
	.C2V_10 (C2V_79_727),
	.C2V_11 (C2V_79_775),
	.C2V_12 (C2V_79_823),
	.C2V_13 (C2V_79_912),
	.C2V_14 (C2V_79_953),
	.C2V_15 (C2V_79_987),
	.C2V_16 (C2V_79_1026),
	.C2V_17 (C2V_79_1100),
	.C2V_18 (C2V_79_1111),
	.C2V_19 (C2V_79_1230),
	.C2V_20 (C2V_79_1231),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU80 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_27_80),
	.V2C_2 (V2C_76_80),
	.V2C_3 (V2C_132_80),
	.V2C_4 (V2C_180_80),
	.V2C_5 (V2C_209_80),
	.V2C_6 (V2C_278_80),
	.V2C_7 (V2C_329_80),
	.V2C_8 (V2C_388_80),
	.V2C_9 (V2C_525_80),
	.V2C_10 (V2C_637_80),
	.V2C_11 (V2C_698_80),
	.V2C_12 (V2C_818_80),
	.V2C_13 (V2C_908_80),
	.V2C_14 (V2C_923_80),
	.V2C_15 (V2C_1002_80),
	.V2C_16 (V2C_1034_80),
	.V2C_17 (V2C_1101_80),
	.V2C_18 (V2C_1132_80),
	.V2C_19 (V2C_1231_80),
	.V2C_20 (V2C_1232_80),
	.C2V_1 (C2V_80_27),
	.C2V_2 (C2V_80_76),
	.C2V_3 (C2V_80_132),
	.C2V_4 (C2V_80_180),
	.C2V_5 (C2V_80_209),
	.C2V_6 (C2V_80_278),
	.C2V_7 (C2V_80_329),
	.C2V_8 (C2V_80_388),
	.C2V_9 (C2V_80_525),
	.C2V_10 (C2V_80_637),
	.C2V_11 (C2V_80_698),
	.C2V_12 (C2V_80_818),
	.C2V_13 (C2V_80_908),
	.C2V_14 (C2V_80_923),
	.C2V_15 (C2V_80_1002),
	.C2V_16 (C2V_80_1034),
	.C2V_17 (C2V_80_1101),
	.C2V_18 (C2V_80_1132),
	.C2V_19 (C2V_80_1231),
	.C2V_20 (C2V_80_1232),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU81 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_22_81),
	.V2C_2 (V2C_49_81),
	.V2C_3 (V2C_114_81),
	.V2C_4 (V2C_148_81),
	.V2C_5 (V2C_214_81),
	.V2C_6 (V2C_281_81),
	.V2C_7 (V2C_378_81),
	.V2C_8 (V2C_385_81),
	.V2C_9 (V2C_544_81),
	.V2C_10 (V2C_601_81),
	.V2C_11 (V2C_629_81),
	.V2C_12 (V2C_733_81),
	.V2C_13 (V2C_912_81),
	.V2C_14 (V2C_956_81),
	.V2C_15 (V2C_981_81),
	.V2C_16 (V2C_1041_81),
	.V2C_17 (V2C_1071_81),
	.V2C_18 (V2C_1116_81),
	.V2C_19 (V2C_1232_81),
	.V2C_20 (V2C_1233_81),
	.C2V_1 (C2V_81_22),
	.C2V_2 (C2V_81_49),
	.C2V_3 (C2V_81_114),
	.C2V_4 (C2V_81_148),
	.C2V_5 (C2V_81_214),
	.C2V_6 (C2V_81_281),
	.C2V_7 (C2V_81_378),
	.C2V_8 (C2V_81_385),
	.C2V_9 (C2V_81_544),
	.C2V_10 (C2V_81_601),
	.C2V_11 (C2V_81_629),
	.C2V_12 (C2V_81_733),
	.C2V_13 (C2V_81_912),
	.C2V_14 (C2V_81_956),
	.C2V_15 (C2V_81_981),
	.C2V_16 (C2V_81_1041),
	.C2V_17 (C2V_81_1071),
	.C2V_18 (C2V_81_1116),
	.C2V_19 (C2V_81_1232),
	.C2V_20 (C2V_81_1233),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU82 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_41_82),
	.V2C_2 (V2C_52_82),
	.V2C_3 (V2C_139_82),
	.V2C_4 (V2C_147_82),
	.V2C_5 (V2C_212_82),
	.V2C_6 (V2C_266_82),
	.V2C_7 (V2C_442_82),
	.V2C_8 (V2C_482_82),
	.V2C_9 (V2C_566_82),
	.V2C_10 (V2C_580_82),
	.V2C_11 (V2C_653_82),
	.V2C_12 (V2C_699_82),
	.V2C_13 (V2C_868_82),
	.V2C_14 (V2C_940_82),
	.V2C_15 (V2C_976_82),
	.V2C_16 (V2C_1054_82),
	.V2C_17 (V2C_1081_82),
	.V2C_18 (V2C_1145_82),
	.V2C_19 (V2C_1233_82),
	.V2C_20 (V2C_1234_82),
	.C2V_1 (C2V_82_41),
	.C2V_2 (C2V_82_52),
	.C2V_3 (C2V_82_139),
	.C2V_4 (C2V_82_147),
	.C2V_5 (C2V_82_212),
	.C2V_6 (C2V_82_266),
	.C2V_7 (C2V_82_442),
	.C2V_8 (C2V_82_482),
	.C2V_9 (C2V_82_566),
	.C2V_10 (C2V_82_580),
	.C2V_11 (C2V_82_653),
	.C2V_12 (C2V_82_699),
	.C2V_13 (C2V_82_868),
	.C2V_14 (C2V_82_940),
	.C2V_15 (C2V_82_976),
	.C2V_16 (C2V_82_1054),
	.C2V_17 (C2V_82_1081),
	.C2V_18 (C2V_82_1145),
	.C2V_19 (C2V_82_1233),
	.C2V_20 (C2V_82_1234),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU83 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_12_83),
	.V2C_2 (V2C_70_83),
	.V2C_3 (V2C_105_83),
	.V2C_4 (V2C_176_83),
	.V2C_5 (V2C_240_83),
	.V2C_6 (V2C_258_83),
	.V2C_7 (V2C_307_83),
	.V2C_8 (V2C_374_83),
	.V2C_9 (V2C_453_83),
	.V2C_10 (V2C_687_83),
	.V2C_11 (V2C_751_83),
	.V2C_12 (V2C_805_83),
	.V2C_13 (V2C_883_83),
	.V2C_14 (V2C_931_83),
	.V2C_15 (V2C_974_83),
	.V2C_16 (V2C_1026_83),
	.V2C_17 (V2C_1075_83),
	.V2C_18 (V2C_1123_83),
	.V2C_19 (V2C_1234_83),
	.V2C_20 (V2C_1235_83),
	.C2V_1 (C2V_83_12),
	.C2V_2 (C2V_83_70),
	.C2V_3 (C2V_83_105),
	.C2V_4 (C2V_83_176),
	.C2V_5 (C2V_83_240),
	.C2V_6 (C2V_83_258),
	.C2V_7 (C2V_83_307),
	.C2V_8 (C2V_83_374),
	.C2V_9 (C2V_83_453),
	.C2V_10 (C2V_83_687),
	.C2V_11 (C2V_83_751),
	.C2V_12 (C2V_83_805),
	.C2V_13 (C2V_83_883),
	.C2V_14 (C2V_83_931),
	.C2V_15 (C2V_83_974),
	.C2V_16 (C2V_83_1026),
	.C2V_17 (C2V_83_1075),
	.C2V_18 (C2V_83_1123),
	.C2V_19 (C2V_83_1234),
	.C2V_20 (C2V_83_1235),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU84 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_43_84),
	.V2C_2 (V2C_67_84),
	.V2C_3 (V2C_107_84),
	.V2C_4 (V2C_175_84),
	.V2C_5 (V2C_209_84),
	.V2C_6 (V2C_288_84),
	.V2C_7 (V2C_293_84),
	.V2C_8 (V2C_445_84),
	.V2C_9 (V2C_542_84),
	.V2C_10 (V2C_623_84),
	.V2C_11 (V2C_779_84),
	.V2C_12 (V2C_855_84),
	.V2C_13 (V2C_888_84),
	.V2C_14 (V2C_950_84),
	.V2C_15 (V2C_985_84),
	.V2C_16 (V2C_1052_84),
	.V2C_17 (V2C_1068_84),
	.V2C_18 (V2C_1118_84),
	.V2C_19 (V2C_1235_84),
	.V2C_20 (V2C_1236_84),
	.C2V_1 (C2V_84_43),
	.C2V_2 (C2V_84_67),
	.C2V_3 (C2V_84_107),
	.C2V_4 (C2V_84_175),
	.C2V_5 (C2V_84_209),
	.C2V_6 (C2V_84_288),
	.C2V_7 (C2V_84_293),
	.C2V_8 (C2V_84_445),
	.C2V_9 (C2V_84_542),
	.C2V_10 (C2V_84_623),
	.C2V_11 (C2V_84_779),
	.C2V_12 (C2V_84_855),
	.C2V_13 (C2V_84_888),
	.C2V_14 (C2V_84_950),
	.C2V_15 (C2V_84_985),
	.C2V_16 (C2V_84_1052),
	.C2V_17 (C2V_84_1068),
	.C2V_18 (C2V_84_1118),
	.C2V_19 (C2V_84_1235),
	.C2V_20 (C2V_84_1236),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU85 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_19_85),
	.V2C_2 (V2C_55_85),
	.V2C_3 (V2C_123_85),
	.V2C_4 (V2C_184_85),
	.V2C_5 (V2C_198_85),
	.V2C_6 (V2C_241_85),
	.V2C_7 (V2C_341_85),
	.V2C_8 (V2C_395_85),
	.V2C_9 (V2C_492_85),
	.V2C_10 (V2C_728_85),
	.V2C_11 (V2C_776_85),
	.V2C_12 (V2C_824_85),
	.V2C_13 (V2C_865_85),
	.V2C_14 (V2C_954_85),
	.V2C_15 (V2C_988_85),
	.V2C_16 (V2C_1027_85),
	.V2C_17 (V2C_1101_85),
	.V2C_18 (V2C_1112_85),
	.V2C_19 (V2C_1236_85),
	.V2C_20 (V2C_1237_85),
	.C2V_1 (C2V_85_19),
	.C2V_2 (C2V_85_55),
	.C2V_3 (C2V_85_123),
	.C2V_4 (C2V_85_184),
	.C2V_5 (C2V_85_198),
	.C2V_6 (C2V_85_241),
	.C2V_7 (C2V_85_341),
	.C2V_8 (C2V_85_395),
	.C2V_9 (C2V_85_492),
	.C2V_10 (C2V_85_728),
	.C2V_11 (C2V_85_776),
	.C2V_12 (C2V_85_824),
	.C2V_13 (C2V_85_865),
	.C2V_14 (C2V_85_954),
	.C2V_15 (C2V_85_988),
	.C2V_16 (C2V_85_1027),
	.C2V_17 (C2V_85_1101),
	.C2V_18 (C2V_85_1112),
	.C2V_19 (C2V_85_1236),
	.C2V_20 (C2V_85_1237),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU86 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_28_86),
	.V2C_2 (V2C_77_86),
	.V2C_3 (V2C_133_86),
	.V2C_4 (V2C_181_86),
	.V2C_5 (V2C_210_86),
	.V2C_6 (V2C_279_86),
	.V2C_7 (V2C_330_86),
	.V2C_8 (V2C_389_86),
	.V2C_9 (V2C_526_86),
	.V2C_10 (V2C_638_86),
	.V2C_11 (V2C_699_86),
	.V2C_12 (V2C_819_86),
	.V2C_13 (V2C_909_86),
	.V2C_14 (V2C_924_86),
	.V2C_15 (V2C_1003_86),
	.V2C_16 (V2C_1035_86),
	.V2C_17 (V2C_1102_86),
	.V2C_18 (V2C_1133_86),
	.V2C_19 (V2C_1237_86),
	.V2C_20 (V2C_1238_86),
	.C2V_1 (C2V_86_28),
	.C2V_2 (C2V_86_77),
	.C2V_3 (C2V_86_133),
	.C2V_4 (C2V_86_181),
	.C2V_5 (C2V_86_210),
	.C2V_6 (C2V_86_279),
	.C2V_7 (C2V_86_330),
	.C2V_8 (C2V_86_389),
	.C2V_9 (C2V_86_526),
	.C2V_10 (C2V_86_638),
	.C2V_11 (C2V_86_699),
	.C2V_12 (C2V_86_819),
	.C2V_13 (C2V_86_909),
	.C2V_14 (C2V_86_924),
	.C2V_15 (C2V_86_1003),
	.C2V_16 (C2V_86_1035),
	.C2V_17 (C2V_86_1102),
	.C2V_18 (C2V_86_1133),
	.C2V_19 (C2V_86_1237),
	.C2V_20 (C2V_86_1238),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU87 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_23_87),
	.V2C_2 (V2C_50_87),
	.V2C_3 (V2C_115_87),
	.V2C_4 (V2C_149_87),
	.V2C_5 (V2C_215_87),
	.V2C_6 (V2C_282_87),
	.V2C_7 (V2C_379_87),
	.V2C_8 (V2C_386_87),
	.V2C_9 (V2C_545_87),
	.V2C_10 (V2C_602_87),
	.V2C_11 (V2C_630_87),
	.V2C_12 (V2C_734_87),
	.V2C_13 (V2C_865_87),
	.V2C_14 (V2C_957_87),
	.V2C_15 (V2C_982_87),
	.V2C_16 (V2C_1042_87),
	.V2C_17 (V2C_1072_87),
	.V2C_18 (V2C_1117_87),
	.V2C_19 (V2C_1238_87),
	.V2C_20 (V2C_1239_87),
	.C2V_1 (C2V_87_23),
	.C2V_2 (C2V_87_50),
	.C2V_3 (C2V_87_115),
	.C2V_4 (C2V_87_149),
	.C2V_5 (C2V_87_215),
	.C2V_6 (C2V_87_282),
	.C2V_7 (C2V_87_379),
	.C2V_8 (C2V_87_386),
	.C2V_9 (C2V_87_545),
	.C2V_10 (C2V_87_602),
	.C2V_11 (C2V_87_630),
	.C2V_12 (C2V_87_734),
	.C2V_13 (C2V_87_865),
	.C2V_14 (C2V_87_957),
	.C2V_15 (C2V_87_982),
	.C2V_16 (C2V_87_1042),
	.C2V_17 (C2V_87_1072),
	.C2V_18 (C2V_87_1117),
	.C2V_19 (C2V_87_1238),
	.C2V_20 (C2V_87_1239),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU88 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_42_88),
	.V2C_2 (V2C_53_88),
	.V2C_3 (V2C_140_88),
	.V2C_4 (V2C_148_88),
	.V2C_5 (V2C_213_88),
	.V2C_6 (V2C_267_88),
	.V2C_7 (V2C_443_88),
	.V2C_8 (V2C_483_88),
	.V2C_9 (V2C_567_88),
	.V2C_10 (V2C_581_88),
	.V2C_11 (V2C_654_88),
	.V2C_12 (V2C_700_88),
	.V2C_13 (V2C_869_88),
	.V2C_14 (V2C_941_88),
	.V2C_15 (V2C_977_88),
	.V2C_16 (V2C_1055_88),
	.V2C_17 (V2C_1082_88),
	.V2C_18 (V2C_1146_88),
	.V2C_19 (V2C_1239_88),
	.V2C_20 (V2C_1240_88),
	.C2V_1 (C2V_88_42),
	.C2V_2 (C2V_88_53),
	.C2V_3 (C2V_88_140),
	.C2V_4 (C2V_88_148),
	.C2V_5 (C2V_88_213),
	.C2V_6 (C2V_88_267),
	.C2V_7 (C2V_88_443),
	.C2V_8 (C2V_88_483),
	.C2V_9 (C2V_88_567),
	.C2V_10 (C2V_88_581),
	.C2V_11 (C2V_88_654),
	.C2V_12 (C2V_88_700),
	.C2V_13 (C2V_88_869),
	.C2V_14 (C2V_88_941),
	.C2V_15 (C2V_88_977),
	.C2V_16 (C2V_88_1055),
	.C2V_17 (C2V_88_1082),
	.C2V_18 (C2V_88_1146),
	.C2V_19 (C2V_88_1239),
	.C2V_20 (C2V_88_1240),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU89 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_13_89),
	.V2C_2 (V2C_71_89),
	.V2C_3 (V2C_106_89),
	.V2C_4 (V2C_177_89),
	.V2C_5 (V2C_193_89),
	.V2C_6 (V2C_259_89),
	.V2C_7 (V2C_308_89),
	.V2C_8 (V2C_375_89),
	.V2C_9 (V2C_454_89),
	.V2C_10 (V2C_688_89),
	.V2C_11 (V2C_752_89),
	.V2C_12 (V2C_806_89),
	.V2C_13 (V2C_884_89),
	.V2C_14 (V2C_932_89),
	.V2C_15 (V2C_975_89),
	.V2C_16 (V2C_1027_89),
	.V2C_17 (V2C_1076_89),
	.V2C_18 (V2C_1124_89),
	.V2C_19 (V2C_1240_89),
	.V2C_20 (V2C_1241_89),
	.C2V_1 (C2V_89_13),
	.C2V_2 (C2V_89_71),
	.C2V_3 (C2V_89_106),
	.C2V_4 (C2V_89_177),
	.C2V_5 (C2V_89_193),
	.C2V_6 (C2V_89_259),
	.C2V_7 (C2V_89_308),
	.C2V_8 (C2V_89_375),
	.C2V_9 (C2V_89_454),
	.C2V_10 (C2V_89_688),
	.C2V_11 (C2V_89_752),
	.C2V_12 (C2V_89_806),
	.C2V_13 (C2V_89_884),
	.C2V_14 (C2V_89_932),
	.C2V_15 (C2V_89_975),
	.C2V_16 (C2V_89_1027),
	.C2V_17 (C2V_89_1076),
	.C2V_18 (C2V_89_1124),
	.C2V_19 (C2V_89_1240),
	.C2V_20 (C2V_89_1241),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU90 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_44_90),
	.V2C_2 (V2C_68_90),
	.V2C_3 (V2C_108_90),
	.V2C_4 (V2C_176_90),
	.V2C_5 (V2C_210_90),
	.V2C_6 (V2C_241_90),
	.V2C_7 (V2C_294_90),
	.V2C_8 (V2C_446_90),
	.V2C_9 (V2C_543_90),
	.V2C_10 (V2C_624_90),
	.V2C_11 (V2C_780_90),
	.V2C_12 (V2C_856_90),
	.V2C_13 (V2C_889_90),
	.V2C_14 (V2C_951_90),
	.V2C_15 (V2C_986_90),
	.V2C_16 (V2C_1053_90),
	.V2C_17 (V2C_1069_90),
	.V2C_18 (V2C_1119_90),
	.V2C_19 (V2C_1241_90),
	.V2C_20 (V2C_1242_90),
	.C2V_1 (C2V_90_44),
	.C2V_2 (C2V_90_68),
	.C2V_3 (C2V_90_108),
	.C2V_4 (C2V_90_176),
	.C2V_5 (C2V_90_210),
	.C2V_6 (C2V_90_241),
	.C2V_7 (C2V_90_294),
	.C2V_8 (C2V_90_446),
	.C2V_9 (C2V_90_543),
	.C2V_10 (C2V_90_624),
	.C2V_11 (C2V_90_780),
	.C2V_12 (C2V_90_856),
	.C2V_13 (C2V_90_889),
	.C2V_14 (C2V_90_951),
	.C2V_15 (C2V_90_986),
	.C2V_16 (C2V_90_1053),
	.C2V_17 (C2V_90_1069),
	.C2V_18 (C2V_90_1119),
	.C2V_19 (C2V_90_1241),
	.C2V_20 (C2V_90_1242),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU91 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_20_91),
	.V2C_2 (V2C_56_91),
	.V2C_3 (V2C_124_91),
	.V2C_4 (V2C_185_91),
	.V2C_5 (V2C_199_91),
	.V2C_6 (V2C_242_91),
	.V2C_7 (V2C_342_91),
	.V2C_8 (V2C_396_91),
	.V2C_9 (V2C_493_91),
	.V2C_10 (V2C_729_91),
	.V2C_11 (V2C_777_91),
	.V2C_12 (V2C_825_91),
	.V2C_13 (V2C_866_91),
	.V2C_14 (V2C_955_91),
	.V2C_15 (V2C_989_91),
	.V2C_16 (V2C_1028_91),
	.V2C_17 (V2C_1102_91),
	.V2C_18 (V2C_1113_91),
	.V2C_19 (V2C_1242_91),
	.V2C_20 (V2C_1243_91),
	.C2V_1 (C2V_91_20),
	.C2V_2 (C2V_91_56),
	.C2V_3 (C2V_91_124),
	.C2V_4 (C2V_91_185),
	.C2V_5 (C2V_91_199),
	.C2V_6 (C2V_91_242),
	.C2V_7 (C2V_91_342),
	.C2V_8 (C2V_91_396),
	.C2V_9 (C2V_91_493),
	.C2V_10 (C2V_91_729),
	.C2V_11 (C2V_91_777),
	.C2V_12 (C2V_91_825),
	.C2V_13 (C2V_91_866),
	.C2V_14 (C2V_91_955),
	.C2V_15 (C2V_91_989),
	.C2V_16 (C2V_91_1028),
	.C2V_17 (C2V_91_1102),
	.C2V_18 (C2V_91_1113),
	.C2V_19 (C2V_91_1242),
	.C2V_20 (C2V_91_1243),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU92 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_29_92),
	.V2C_2 (V2C_78_92),
	.V2C_3 (V2C_134_92),
	.V2C_4 (V2C_182_92),
	.V2C_5 (V2C_211_92),
	.V2C_6 (V2C_280_92),
	.V2C_7 (V2C_331_92),
	.V2C_8 (V2C_390_92),
	.V2C_9 (V2C_527_92),
	.V2C_10 (V2C_639_92),
	.V2C_11 (V2C_700_92),
	.V2C_12 (V2C_820_92),
	.V2C_13 (V2C_910_92),
	.V2C_14 (V2C_925_92),
	.V2C_15 (V2C_1004_92),
	.V2C_16 (V2C_1036_92),
	.V2C_17 (V2C_1103_92),
	.V2C_18 (V2C_1134_92),
	.V2C_19 (V2C_1243_92),
	.V2C_20 (V2C_1244_92),
	.C2V_1 (C2V_92_29),
	.C2V_2 (C2V_92_78),
	.C2V_3 (C2V_92_134),
	.C2V_4 (C2V_92_182),
	.C2V_5 (C2V_92_211),
	.C2V_6 (C2V_92_280),
	.C2V_7 (C2V_92_331),
	.C2V_8 (C2V_92_390),
	.C2V_9 (C2V_92_527),
	.C2V_10 (C2V_92_639),
	.C2V_11 (C2V_92_700),
	.C2V_12 (C2V_92_820),
	.C2V_13 (C2V_92_910),
	.C2V_14 (C2V_92_925),
	.C2V_15 (C2V_92_1004),
	.C2V_16 (C2V_92_1036),
	.C2V_17 (C2V_92_1103),
	.C2V_18 (C2V_92_1134),
	.C2V_19 (C2V_92_1243),
	.C2V_20 (C2V_92_1244),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU93 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_24_93),
	.V2C_2 (V2C_51_93),
	.V2C_3 (V2C_116_93),
	.V2C_4 (V2C_150_93),
	.V2C_5 (V2C_216_93),
	.V2C_6 (V2C_283_93),
	.V2C_7 (V2C_380_93),
	.V2C_8 (V2C_387_93),
	.V2C_9 (V2C_546_93),
	.V2C_10 (V2C_603_93),
	.V2C_11 (V2C_631_93),
	.V2C_12 (V2C_735_93),
	.V2C_13 (V2C_866_93),
	.V2C_14 (V2C_958_93),
	.V2C_15 (V2C_983_93),
	.V2C_16 (V2C_1043_93),
	.V2C_17 (V2C_1073_93),
	.V2C_18 (V2C_1118_93),
	.V2C_19 (V2C_1244_93),
	.V2C_20 (V2C_1245_93),
	.C2V_1 (C2V_93_24),
	.C2V_2 (C2V_93_51),
	.C2V_3 (C2V_93_116),
	.C2V_4 (C2V_93_150),
	.C2V_5 (C2V_93_216),
	.C2V_6 (C2V_93_283),
	.C2V_7 (C2V_93_380),
	.C2V_8 (C2V_93_387),
	.C2V_9 (C2V_93_546),
	.C2V_10 (C2V_93_603),
	.C2V_11 (C2V_93_631),
	.C2V_12 (C2V_93_735),
	.C2V_13 (C2V_93_866),
	.C2V_14 (C2V_93_958),
	.C2V_15 (C2V_93_983),
	.C2V_16 (C2V_93_1043),
	.C2V_17 (C2V_93_1073),
	.C2V_18 (C2V_93_1118),
	.C2V_19 (C2V_93_1244),
	.C2V_20 (C2V_93_1245),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU94 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_43_94),
	.V2C_2 (V2C_54_94),
	.V2C_3 (V2C_141_94),
	.V2C_4 (V2C_149_94),
	.V2C_5 (V2C_214_94),
	.V2C_6 (V2C_268_94),
	.V2C_7 (V2C_444_94),
	.V2C_8 (V2C_484_94),
	.V2C_9 (V2C_568_94),
	.V2C_10 (V2C_582_94),
	.V2C_11 (V2C_655_94),
	.V2C_12 (V2C_701_94),
	.V2C_13 (V2C_870_94),
	.V2C_14 (V2C_942_94),
	.V2C_15 (V2C_978_94),
	.V2C_16 (V2C_1056_94),
	.V2C_17 (V2C_1083_94),
	.V2C_18 (V2C_1147_94),
	.V2C_19 (V2C_1245_94),
	.V2C_20 (V2C_1246_94),
	.C2V_1 (C2V_94_43),
	.C2V_2 (C2V_94_54),
	.C2V_3 (C2V_94_141),
	.C2V_4 (C2V_94_149),
	.C2V_5 (C2V_94_214),
	.C2V_6 (C2V_94_268),
	.C2V_7 (C2V_94_444),
	.C2V_8 (C2V_94_484),
	.C2V_9 (C2V_94_568),
	.C2V_10 (C2V_94_582),
	.C2V_11 (C2V_94_655),
	.C2V_12 (C2V_94_701),
	.C2V_13 (C2V_94_870),
	.C2V_14 (C2V_94_942),
	.C2V_15 (C2V_94_978),
	.C2V_16 (C2V_94_1056),
	.C2V_17 (C2V_94_1083),
	.C2V_18 (C2V_94_1147),
	.C2V_19 (C2V_94_1245),
	.C2V_20 (C2V_94_1246),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU95 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_14_95),
	.V2C_2 (V2C_72_95),
	.V2C_3 (V2C_107_95),
	.V2C_4 (V2C_178_95),
	.V2C_5 (V2C_194_95),
	.V2C_6 (V2C_260_95),
	.V2C_7 (V2C_309_95),
	.V2C_8 (V2C_376_95),
	.V2C_9 (V2C_455_95),
	.V2C_10 (V2C_689_95),
	.V2C_11 (V2C_753_95),
	.V2C_12 (V2C_807_95),
	.V2C_13 (V2C_885_95),
	.V2C_14 (V2C_933_95),
	.V2C_15 (V2C_976_95),
	.V2C_16 (V2C_1028_95),
	.V2C_17 (V2C_1077_95),
	.V2C_18 (V2C_1125_95),
	.V2C_19 (V2C_1246_95),
	.V2C_20 (V2C_1247_95),
	.C2V_1 (C2V_95_14),
	.C2V_2 (C2V_95_72),
	.C2V_3 (C2V_95_107),
	.C2V_4 (C2V_95_178),
	.C2V_5 (C2V_95_194),
	.C2V_6 (C2V_95_260),
	.C2V_7 (C2V_95_309),
	.C2V_8 (C2V_95_376),
	.C2V_9 (C2V_95_455),
	.C2V_10 (C2V_95_689),
	.C2V_11 (C2V_95_753),
	.C2V_12 (C2V_95_807),
	.C2V_13 (C2V_95_885),
	.C2V_14 (C2V_95_933),
	.C2V_15 (C2V_95_976),
	.C2V_16 (C2V_95_1028),
	.C2V_17 (C2V_95_1077),
	.C2V_18 (C2V_95_1125),
	.C2V_19 (C2V_95_1246),
	.C2V_20 (C2V_95_1247),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU96 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_45_96),
	.V2C_2 (V2C_69_96),
	.V2C_3 (V2C_109_96),
	.V2C_4 (V2C_177_96),
	.V2C_5 (V2C_211_96),
	.V2C_6 (V2C_242_96),
	.V2C_7 (V2C_295_96),
	.V2C_8 (V2C_447_96),
	.V2C_9 (V2C_544_96),
	.V2C_10 (V2C_577_96),
	.V2C_11 (V2C_781_96),
	.V2C_12 (V2C_857_96),
	.V2C_13 (V2C_890_96),
	.V2C_14 (V2C_952_96),
	.V2C_15 (V2C_987_96),
	.V2C_16 (V2C_1054_96),
	.V2C_17 (V2C_1070_96),
	.V2C_18 (V2C_1120_96),
	.V2C_19 (V2C_1247_96),
	.V2C_20 (V2C_1248_96),
	.C2V_1 (C2V_96_45),
	.C2V_2 (C2V_96_69),
	.C2V_3 (C2V_96_109),
	.C2V_4 (C2V_96_177),
	.C2V_5 (C2V_96_211),
	.C2V_6 (C2V_96_242),
	.C2V_7 (C2V_96_295),
	.C2V_8 (C2V_96_447),
	.C2V_9 (C2V_96_544),
	.C2V_10 (C2V_96_577),
	.C2V_11 (C2V_96_781),
	.C2V_12 (C2V_96_857),
	.C2V_13 (C2V_96_890),
	.C2V_14 (C2V_96_952),
	.C2V_15 (C2V_96_987),
	.C2V_16 (C2V_96_1054),
	.C2V_17 (C2V_96_1070),
	.C2V_18 (C2V_96_1120),
	.C2V_19 (C2V_96_1247),
	.C2V_20 (C2V_96_1248),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU97 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_21_97),
	.V2C_2 (V2C_57_97),
	.V2C_3 (V2C_125_97),
	.V2C_4 (V2C_186_97),
	.V2C_5 (V2C_200_97),
	.V2C_6 (V2C_243_97),
	.V2C_7 (V2C_343_97),
	.V2C_8 (V2C_397_97),
	.V2C_9 (V2C_494_97),
	.V2C_10 (V2C_730_97),
	.V2C_11 (V2C_778_97),
	.V2C_12 (V2C_826_97),
	.V2C_13 (V2C_867_97),
	.V2C_14 (V2C_956_97),
	.V2C_15 (V2C_990_97),
	.V2C_16 (V2C_1029_97),
	.V2C_17 (V2C_1103_97),
	.V2C_18 (V2C_1114_97),
	.V2C_19 (V2C_1248_97),
	.V2C_20 (V2C_1249_97),
	.C2V_1 (C2V_97_21),
	.C2V_2 (C2V_97_57),
	.C2V_3 (C2V_97_125),
	.C2V_4 (C2V_97_186),
	.C2V_5 (C2V_97_200),
	.C2V_6 (C2V_97_243),
	.C2V_7 (C2V_97_343),
	.C2V_8 (C2V_97_397),
	.C2V_9 (C2V_97_494),
	.C2V_10 (C2V_97_730),
	.C2V_11 (C2V_97_778),
	.C2V_12 (C2V_97_826),
	.C2V_13 (C2V_97_867),
	.C2V_14 (C2V_97_956),
	.C2V_15 (C2V_97_990),
	.C2V_16 (C2V_97_1029),
	.C2V_17 (C2V_97_1103),
	.C2V_18 (C2V_97_1114),
	.C2V_19 (C2V_97_1248),
	.C2V_20 (C2V_97_1249),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU98 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_30_98),
	.V2C_2 (V2C_79_98),
	.V2C_3 (V2C_135_98),
	.V2C_4 (V2C_183_98),
	.V2C_5 (V2C_212_98),
	.V2C_6 (V2C_281_98),
	.V2C_7 (V2C_332_98),
	.V2C_8 (V2C_391_98),
	.V2C_9 (V2C_528_98),
	.V2C_10 (V2C_640_98),
	.V2C_11 (V2C_701_98),
	.V2C_12 (V2C_821_98),
	.V2C_13 (V2C_911_98),
	.V2C_14 (V2C_926_98),
	.V2C_15 (V2C_1005_98),
	.V2C_16 (V2C_1037_98),
	.V2C_17 (V2C_1104_98),
	.V2C_18 (V2C_1135_98),
	.V2C_19 (V2C_1249_98),
	.V2C_20 (V2C_1250_98),
	.C2V_1 (C2V_98_30),
	.C2V_2 (C2V_98_79),
	.C2V_3 (C2V_98_135),
	.C2V_4 (C2V_98_183),
	.C2V_5 (C2V_98_212),
	.C2V_6 (C2V_98_281),
	.C2V_7 (C2V_98_332),
	.C2V_8 (C2V_98_391),
	.C2V_9 (C2V_98_528),
	.C2V_10 (C2V_98_640),
	.C2V_11 (C2V_98_701),
	.C2V_12 (C2V_98_821),
	.C2V_13 (C2V_98_911),
	.C2V_14 (C2V_98_926),
	.C2V_15 (C2V_98_1005),
	.C2V_16 (C2V_98_1037),
	.C2V_17 (C2V_98_1104),
	.C2V_18 (C2V_98_1135),
	.C2V_19 (C2V_98_1249),
	.C2V_20 (C2V_98_1250),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU99 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_25_99),
	.V2C_2 (V2C_52_99),
	.V2C_3 (V2C_117_99),
	.V2C_4 (V2C_151_99),
	.V2C_5 (V2C_217_99),
	.V2C_6 (V2C_284_99),
	.V2C_7 (V2C_381_99),
	.V2C_8 (V2C_388_99),
	.V2C_9 (V2C_547_99),
	.V2C_10 (V2C_604_99),
	.V2C_11 (V2C_632_99),
	.V2C_12 (V2C_736_99),
	.V2C_13 (V2C_867_99),
	.V2C_14 (V2C_959_99),
	.V2C_15 (V2C_984_99),
	.V2C_16 (V2C_1044_99),
	.V2C_17 (V2C_1074_99),
	.V2C_18 (V2C_1119_99),
	.V2C_19 (V2C_1250_99),
	.V2C_20 (V2C_1251_99),
	.C2V_1 (C2V_99_25),
	.C2V_2 (C2V_99_52),
	.C2V_3 (C2V_99_117),
	.C2V_4 (C2V_99_151),
	.C2V_5 (C2V_99_217),
	.C2V_6 (C2V_99_284),
	.C2V_7 (C2V_99_381),
	.C2V_8 (C2V_99_388),
	.C2V_9 (C2V_99_547),
	.C2V_10 (C2V_99_604),
	.C2V_11 (C2V_99_632),
	.C2V_12 (C2V_99_736),
	.C2V_13 (C2V_99_867),
	.C2V_14 (C2V_99_959),
	.C2V_15 (C2V_99_984),
	.C2V_16 (C2V_99_1044),
	.C2V_17 (C2V_99_1074),
	.C2V_18 (C2V_99_1119),
	.C2V_19 (C2V_99_1250),
	.C2V_20 (C2V_99_1251),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU100 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_44_100),
	.V2C_2 (V2C_55_100),
	.V2C_3 (V2C_142_100),
	.V2C_4 (V2C_150_100),
	.V2C_5 (V2C_215_100),
	.V2C_6 (V2C_269_100),
	.V2C_7 (V2C_445_100),
	.V2C_8 (V2C_485_100),
	.V2C_9 (V2C_569_100),
	.V2C_10 (V2C_583_100),
	.V2C_11 (V2C_656_100),
	.V2C_12 (V2C_702_100),
	.V2C_13 (V2C_871_100),
	.V2C_14 (V2C_943_100),
	.V2C_15 (V2C_979_100),
	.V2C_16 (V2C_1009_100),
	.V2C_17 (V2C_1084_100),
	.V2C_18 (V2C_1148_100),
	.V2C_19 (V2C_1251_100),
	.V2C_20 (V2C_1252_100),
	.C2V_1 (C2V_100_44),
	.C2V_2 (C2V_100_55),
	.C2V_3 (C2V_100_142),
	.C2V_4 (C2V_100_150),
	.C2V_5 (C2V_100_215),
	.C2V_6 (C2V_100_269),
	.C2V_7 (C2V_100_445),
	.C2V_8 (C2V_100_485),
	.C2V_9 (C2V_100_569),
	.C2V_10 (C2V_100_583),
	.C2V_11 (C2V_100_656),
	.C2V_12 (C2V_100_702),
	.C2V_13 (C2V_100_871),
	.C2V_14 (C2V_100_943),
	.C2V_15 (C2V_100_979),
	.C2V_16 (C2V_100_1009),
	.C2V_17 (C2V_100_1084),
	.C2V_18 (C2V_100_1148),
	.C2V_19 (C2V_100_1251),
	.C2V_20 (C2V_100_1252),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU101 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_15_101),
	.V2C_2 (V2C_73_101),
	.V2C_3 (V2C_108_101),
	.V2C_4 (V2C_179_101),
	.V2C_5 (V2C_195_101),
	.V2C_6 (V2C_261_101),
	.V2C_7 (V2C_310_101),
	.V2C_8 (V2C_377_101),
	.V2C_9 (V2C_456_101),
	.V2C_10 (V2C_690_101),
	.V2C_11 (V2C_754_101),
	.V2C_12 (V2C_808_101),
	.V2C_13 (V2C_886_101),
	.V2C_14 (V2C_934_101),
	.V2C_15 (V2C_977_101),
	.V2C_16 (V2C_1029_101),
	.V2C_17 (V2C_1078_101),
	.V2C_18 (V2C_1126_101),
	.V2C_19 (V2C_1252_101),
	.V2C_20 (V2C_1253_101),
	.C2V_1 (C2V_101_15),
	.C2V_2 (C2V_101_73),
	.C2V_3 (C2V_101_108),
	.C2V_4 (C2V_101_179),
	.C2V_5 (C2V_101_195),
	.C2V_6 (C2V_101_261),
	.C2V_7 (C2V_101_310),
	.C2V_8 (C2V_101_377),
	.C2V_9 (C2V_101_456),
	.C2V_10 (C2V_101_690),
	.C2V_11 (C2V_101_754),
	.C2V_12 (C2V_101_808),
	.C2V_13 (C2V_101_886),
	.C2V_14 (C2V_101_934),
	.C2V_15 (C2V_101_977),
	.C2V_16 (C2V_101_1029),
	.C2V_17 (C2V_101_1078),
	.C2V_18 (C2V_101_1126),
	.C2V_19 (C2V_101_1252),
	.C2V_20 (C2V_101_1253),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU102 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_46_102),
	.V2C_2 (V2C_70_102),
	.V2C_3 (V2C_110_102),
	.V2C_4 (V2C_178_102),
	.V2C_5 (V2C_212_102),
	.V2C_6 (V2C_243_102),
	.V2C_7 (V2C_296_102),
	.V2C_8 (V2C_448_102),
	.V2C_9 (V2C_545_102),
	.V2C_10 (V2C_578_102),
	.V2C_11 (V2C_782_102),
	.V2C_12 (V2C_858_102),
	.V2C_13 (V2C_891_102),
	.V2C_14 (V2C_953_102),
	.V2C_15 (V2C_988_102),
	.V2C_16 (V2C_1055_102),
	.V2C_17 (V2C_1071_102),
	.V2C_18 (V2C_1121_102),
	.V2C_19 (V2C_1253_102),
	.V2C_20 (V2C_1254_102),
	.C2V_1 (C2V_102_46),
	.C2V_2 (C2V_102_70),
	.C2V_3 (C2V_102_110),
	.C2V_4 (C2V_102_178),
	.C2V_5 (C2V_102_212),
	.C2V_6 (C2V_102_243),
	.C2V_7 (C2V_102_296),
	.C2V_8 (C2V_102_448),
	.C2V_9 (C2V_102_545),
	.C2V_10 (C2V_102_578),
	.C2V_11 (C2V_102_782),
	.C2V_12 (C2V_102_858),
	.C2V_13 (C2V_102_891),
	.C2V_14 (C2V_102_953),
	.C2V_15 (C2V_102_988),
	.C2V_16 (C2V_102_1055),
	.C2V_17 (C2V_102_1071),
	.C2V_18 (C2V_102_1121),
	.C2V_19 (C2V_102_1253),
	.C2V_20 (C2V_102_1254),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU103 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_22_103),
	.V2C_2 (V2C_58_103),
	.V2C_3 (V2C_126_103),
	.V2C_4 (V2C_187_103),
	.V2C_5 (V2C_201_103),
	.V2C_6 (V2C_244_103),
	.V2C_7 (V2C_344_103),
	.V2C_8 (V2C_398_103),
	.V2C_9 (V2C_495_103),
	.V2C_10 (V2C_731_103),
	.V2C_11 (V2C_779_103),
	.V2C_12 (V2C_827_103),
	.V2C_13 (V2C_868_103),
	.V2C_14 (V2C_957_103),
	.V2C_15 (V2C_991_103),
	.V2C_16 (V2C_1030_103),
	.V2C_17 (V2C_1104_103),
	.V2C_18 (V2C_1115_103),
	.V2C_19 (V2C_1254_103),
	.V2C_20 (V2C_1255_103),
	.C2V_1 (C2V_103_22),
	.C2V_2 (C2V_103_58),
	.C2V_3 (C2V_103_126),
	.C2V_4 (C2V_103_187),
	.C2V_5 (C2V_103_201),
	.C2V_6 (C2V_103_244),
	.C2V_7 (C2V_103_344),
	.C2V_8 (C2V_103_398),
	.C2V_9 (C2V_103_495),
	.C2V_10 (C2V_103_731),
	.C2V_11 (C2V_103_779),
	.C2V_12 (C2V_103_827),
	.C2V_13 (C2V_103_868),
	.C2V_14 (C2V_103_957),
	.C2V_15 (C2V_103_991),
	.C2V_16 (C2V_103_1030),
	.C2V_17 (C2V_103_1104),
	.C2V_18 (C2V_103_1115),
	.C2V_19 (C2V_103_1254),
	.C2V_20 (C2V_103_1255),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU104 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_31_104),
	.V2C_2 (V2C_80_104),
	.V2C_3 (V2C_136_104),
	.V2C_4 (V2C_184_104),
	.V2C_5 (V2C_213_104),
	.V2C_6 (V2C_282_104),
	.V2C_7 (V2C_333_104),
	.V2C_8 (V2C_392_104),
	.V2C_9 (V2C_481_104),
	.V2C_10 (V2C_641_104),
	.V2C_11 (V2C_702_104),
	.V2C_12 (V2C_822_104),
	.V2C_13 (V2C_912_104),
	.V2C_14 (V2C_927_104),
	.V2C_15 (V2C_1006_104),
	.V2C_16 (V2C_1038_104),
	.V2C_17 (V2C_1057_104),
	.V2C_18 (V2C_1136_104),
	.V2C_19 (V2C_1255_104),
	.V2C_20 (V2C_1256_104),
	.C2V_1 (C2V_104_31),
	.C2V_2 (C2V_104_80),
	.C2V_3 (C2V_104_136),
	.C2V_4 (C2V_104_184),
	.C2V_5 (C2V_104_213),
	.C2V_6 (C2V_104_282),
	.C2V_7 (C2V_104_333),
	.C2V_8 (C2V_104_392),
	.C2V_9 (C2V_104_481),
	.C2V_10 (C2V_104_641),
	.C2V_11 (C2V_104_702),
	.C2V_12 (C2V_104_822),
	.C2V_13 (C2V_104_912),
	.C2V_14 (C2V_104_927),
	.C2V_15 (C2V_104_1006),
	.C2V_16 (C2V_104_1038),
	.C2V_17 (C2V_104_1057),
	.C2V_18 (C2V_104_1136),
	.C2V_19 (C2V_104_1255),
	.C2V_20 (C2V_104_1256),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU105 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_26_105),
	.V2C_2 (V2C_53_105),
	.V2C_3 (V2C_118_105),
	.V2C_4 (V2C_152_105),
	.V2C_5 (V2C_218_105),
	.V2C_6 (V2C_285_105),
	.V2C_7 (V2C_382_105),
	.V2C_8 (V2C_389_105),
	.V2C_9 (V2C_548_105),
	.V2C_10 (V2C_605_105),
	.V2C_11 (V2C_633_105),
	.V2C_12 (V2C_737_105),
	.V2C_13 (V2C_868_105),
	.V2C_14 (V2C_960_105),
	.V2C_15 (V2C_985_105),
	.V2C_16 (V2C_1045_105),
	.V2C_17 (V2C_1075_105),
	.V2C_18 (V2C_1120_105),
	.V2C_19 (V2C_1256_105),
	.V2C_20 (V2C_1257_105),
	.C2V_1 (C2V_105_26),
	.C2V_2 (C2V_105_53),
	.C2V_3 (C2V_105_118),
	.C2V_4 (C2V_105_152),
	.C2V_5 (C2V_105_218),
	.C2V_6 (C2V_105_285),
	.C2V_7 (C2V_105_382),
	.C2V_8 (C2V_105_389),
	.C2V_9 (C2V_105_548),
	.C2V_10 (C2V_105_605),
	.C2V_11 (C2V_105_633),
	.C2V_12 (C2V_105_737),
	.C2V_13 (C2V_105_868),
	.C2V_14 (C2V_105_960),
	.C2V_15 (C2V_105_985),
	.C2V_16 (C2V_105_1045),
	.C2V_17 (C2V_105_1075),
	.C2V_18 (C2V_105_1120),
	.C2V_19 (C2V_105_1256),
	.C2V_20 (C2V_105_1257),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU106 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_45_106),
	.V2C_2 (V2C_56_106),
	.V2C_3 (V2C_143_106),
	.V2C_4 (V2C_151_106),
	.V2C_5 (V2C_216_106),
	.V2C_6 (V2C_270_106),
	.V2C_7 (V2C_446_106),
	.V2C_8 (V2C_486_106),
	.V2C_9 (V2C_570_106),
	.V2C_10 (V2C_584_106),
	.V2C_11 (V2C_657_106),
	.V2C_12 (V2C_703_106),
	.V2C_13 (V2C_872_106),
	.V2C_14 (V2C_944_106),
	.V2C_15 (V2C_980_106),
	.V2C_16 (V2C_1010_106),
	.V2C_17 (V2C_1085_106),
	.V2C_18 (V2C_1149_106),
	.V2C_19 (V2C_1257_106),
	.V2C_20 (V2C_1258_106),
	.C2V_1 (C2V_106_45),
	.C2V_2 (C2V_106_56),
	.C2V_3 (C2V_106_143),
	.C2V_4 (C2V_106_151),
	.C2V_5 (C2V_106_216),
	.C2V_6 (C2V_106_270),
	.C2V_7 (C2V_106_446),
	.C2V_8 (C2V_106_486),
	.C2V_9 (C2V_106_570),
	.C2V_10 (C2V_106_584),
	.C2V_11 (C2V_106_657),
	.C2V_12 (C2V_106_703),
	.C2V_13 (C2V_106_872),
	.C2V_14 (C2V_106_944),
	.C2V_15 (C2V_106_980),
	.C2V_16 (C2V_106_1010),
	.C2V_17 (C2V_106_1085),
	.C2V_18 (C2V_106_1149),
	.C2V_19 (C2V_106_1257),
	.C2V_20 (C2V_106_1258),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU107 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_16_107),
	.V2C_2 (V2C_74_107),
	.V2C_3 (V2C_109_107),
	.V2C_4 (V2C_180_107),
	.V2C_5 (V2C_196_107),
	.V2C_6 (V2C_262_107),
	.V2C_7 (V2C_311_107),
	.V2C_8 (V2C_378_107),
	.V2C_9 (V2C_457_107),
	.V2C_10 (V2C_691_107),
	.V2C_11 (V2C_755_107),
	.V2C_12 (V2C_809_107),
	.V2C_13 (V2C_887_107),
	.V2C_14 (V2C_935_107),
	.V2C_15 (V2C_978_107),
	.V2C_16 (V2C_1030_107),
	.V2C_17 (V2C_1079_107),
	.V2C_18 (V2C_1127_107),
	.V2C_19 (V2C_1258_107),
	.V2C_20 (V2C_1259_107),
	.C2V_1 (C2V_107_16),
	.C2V_2 (C2V_107_74),
	.C2V_3 (C2V_107_109),
	.C2V_4 (C2V_107_180),
	.C2V_5 (C2V_107_196),
	.C2V_6 (C2V_107_262),
	.C2V_7 (C2V_107_311),
	.C2V_8 (C2V_107_378),
	.C2V_9 (C2V_107_457),
	.C2V_10 (C2V_107_691),
	.C2V_11 (C2V_107_755),
	.C2V_12 (C2V_107_809),
	.C2V_13 (C2V_107_887),
	.C2V_14 (C2V_107_935),
	.C2V_15 (C2V_107_978),
	.C2V_16 (C2V_107_1030),
	.C2V_17 (C2V_107_1079),
	.C2V_18 (C2V_107_1127),
	.C2V_19 (C2V_107_1258),
	.C2V_20 (C2V_107_1259),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU108 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_47_108),
	.V2C_2 (V2C_71_108),
	.V2C_3 (V2C_111_108),
	.V2C_4 (V2C_179_108),
	.V2C_5 (V2C_213_108),
	.V2C_6 (V2C_244_108),
	.V2C_7 (V2C_297_108),
	.V2C_8 (V2C_449_108),
	.V2C_9 (V2C_546_108),
	.V2C_10 (V2C_579_108),
	.V2C_11 (V2C_783_108),
	.V2C_12 (V2C_859_108),
	.V2C_13 (V2C_892_108),
	.V2C_14 (V2C_954_108),
	.V2C_15 (V2C_989_108),
	.V2C_16 (V2C_1056_108),
	.V2C_17 (V2C_1072_108),
	.V2C_18 (V2C_1122_108),
	.V2C_19 (V2C_1259_108),
	.V2C_20 (V2C_1260_108),
	.C2V_1 (C2V_108_47),
	.C2V_2 (C2V_108_71),
	.C2V_3 (C2V_108_111),
	.C2V_4 (C2V_108_179),
	.C2V_5 (C2V_108_213),
	.C2V_6 (C2V_108_244),
	.C2V_7 (C2V_108_297),
	.C2V_8 (C2V_108_449),
	.C2V_9 (C2V_108_546),
	.C2V_10 (C2V_108_579),
	.C2V_11 (C2V_108_783),
	.C2V_12 (C2V_108_859),
	.C2V_13 (C2V_108_892),
	.C2V_14 (C2V_108_954),
	.C2V_15 (C2V_108_989),
	.C2V_16 (C2V_108_1056),
	.C2V_17 (C2V_108_1072),
	.C2V_18 (C2V_108_1122),
	.C2V_19 (C2V_108_1259),
	.C2V_20 (C2V_108_1260),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU109 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_23_109),
	.V2C_2 (V2C_59_109),
	.V2C_3 (V2C_127_109),
	.V2C_4 (V2C_188_109),
	.V2C_5 (V2C_202_109),
	.V2C_6 (V2C_245_109),
	.V2C_7 (V2C_345_109),
	.V2C_8 (V2C_399_109),
	.V2C_9 (V2C_496_109),
	.V2C_10 (V2C_732_109),
	.V2C_11 (V2C_780_109),
	.V2C_12 (V2C_828_109),
	.V2C_13 (V2C_869_109),
	.V2C_14 (V2C_958_109),
	.V2C_15 (V2C_992_109),
	.V2C_16 (V2C_1031_109),
	.V2C_17 (V2C_1057_109),
	.V2C_18 (V2C_1116_109),
	.V2C_19 (V2C_1260_109),
	.V2C_20 (V2C_1261_109),
	.C2V_1 (C2V_109_23),
	.C2V_2 (C2V_109_59),
	.C2V_3 (C2V_109_127),
	.C2V_4 (C2V_109_188),
	.C2V_5 (C2V_109_202),
	.C2V_6 (C2V_109_245),
	.C2V_7 (C2V_109_345),
	.C2V_8 (C2V_109_399),
	.C2V_9 (C2V_109_496),
	.C2V_10 (C2V_109_732),
	.C2V_11 (C2V_109_780),
	.C2V_12 (C2V_109_828),
	.C2V_13 (C2V_109_869),
	.C2V_14 (C2V_109_958),
	.C2V_15 (C2V_109_992),
	.C2V_16 (C2V_109_1031),
	.C2V_17 (C2V_109_1057),
	.C2V_18 (C2V_109_1116),
	.C2V_19 (C2V_109_1260),
	.C2V_20 (C2V_109_1261),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU110 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_32_110),
	.V2C_2 (V2C_81_110),
	.V2C_3 (V2C_137_110),
	.V2C_4 (V2C_185_110),
	.V2C_5 (V2C_214_110),
	.V2C_6 (V2C_283_110),
	.V2C_7 (V2C_334_110),
	.V2C_8 (V2C_393_110),
	.V2C_9 (V2C_482_110),
	.V2C_10 (V2C_642_110),
	.V2C_11 (V2C_703_110),
	.V2C_12 (V2C_823_110),
	.V2C_13 (V2C_865_110),
	.V2C_14 (V2C_928_110),
	.V2C_15 (V2C_1007_110),
	.V2C_16 (V2C_1039_110),
	.V2C_17 (V2C_1058_110),
	.V2C_18 (V2C_1137_110),
	.V2C_19 (V2C_1261_110),
	.V2C_20 (V2C_1262_110),
	.C2V_1 (C2V_110_32),
	.C2V_2 (C2V_110_81),
	.C2V_3 (C2V_110_137),
	.C2V_4 (C2V_110_185),
	.C2V_5 (C2V_110_214),
	.C2V_6 (C2V_110_283),
	.C2V_7 (C2V_110_334),
	.C2V_8 (C2V_110_393),
	.C2V_9 (C2V_110_482),
	.C2V_10 (C2V_110_642),
	.C2V_11 (C2V_110_703),
	.C2V_12 (C2V_110_823),
	.C2V_13 (C2V_110_865),
	.C2V_14 (C2V_110_928),
	.C2V_15 (C2V_110_1007),
	.C2V_16 (C2V_110_1039),
	.C2V_17 (C2V_110_1058),
	.C2V_18 (C2V_110_1137),
	.C2V_19 (C2V_110_1261),
	.C2V_20 (C2V_110_1262),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU111 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_27_111),
	.V2C_2 (V2C_54_111),
	.V2C_3 (V2C_119_111),
	.V2C_4 (V2C_153_111),
	.V2C_5 (V2C_219_111),
	.V2C_6 (V2C_286_111),
	.V2C_7 (V2C_383_111),
	.V2C_8 (V2C_390_111),
	.V2C_9 (V2C_549_111),
	.V2C_10 (V2C_606_111),
	.V2C_11 (V2C_634_111),
	.V2C_12 (V2C_738_111),
	.V2C_13 (V2C_869_111),
	.V2C_14 (V2C_913_111),
	.V2C_15 (V2C_986_111),
	.V2C_16 (V2C_1046_111),
	.V2C_17 (V2C_1076_111),
	.V2C_18 (V2C_1121_111),
	.V2C_19 (V2C_1262_111),
	.V2C_20 (V2C_1263_111),
	.C2V_1 (C2V_111_27),
	.C2V_2 (C2V_111_54),
	.C2V_3 (C2V_111_119),
	.C2V_4 (C2V_111_153),
	.C2V_5 (C2V_111_219),
	.C2V_6 (C2V_111_286),
	.C2V_7 (C2V_111_383),
	.C2V_8 (C2V_111_390),
	.C2V_9 (C2V_111_549),
	.C2V_10 (C2V_111_606),
	.C2V_11 (C2V_111_634),
	.C2V_12 (C2V_111_738),
	.C2V_13 (C2V_111_869),
	.C2V_14 (C2V_111_913),
	.C2V_15 (C2V_111_986),
	.C2V_16 (C2V_111_1046),
	.C2V_17 (C2V_111_1076),
	.C2V_18 (C2V_111_1121),
	.C2V_19 (C2V_111_1262),
	.C2V_20 (C2V_111_1263),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU112 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_46_112),
	.V2C_2 (V2C_57_112),
	.V2C_3 (V2C_144_112),
	.V2C_4 (V2C_152_112),
	.V2C_5 (V2C_217_112),
	.V2C_6 (V2C_271_112),
	.V2C_7 (V2C_447_112),
	.V2C_8 (V2C_487_112),
	.V2C_9 (V2C_571_112),
	.V2C_10 (V2C_585_112),
	.V2C_11 (V2C_658_112),
	.V2C_12 (V2C_704_112),
	.V2C_13 (V2C_873_112),
	.V2C_14 (V2C_945_112),
	.V2C_15 (V2C_981_112),
	.V2C_16 (V2C_1011_112),
	.V2C_17 (V2C_1086_112),
	.V2C_18 (V2C_1150_112),
	.V2C_19 (V2C_1263_112),
	.V2C_20 (V2C_1264_112),
	.C2V_1 (C2V_112_46),
	.C2V_2 (C2V_112_57),
	.C2V_3 (C2V_112_144),
	.C2V_4 (C2V_112_152),
	.C2V_5 (C2V_112_217),
	.C2V_6 (C2V_112_271),
	.C2V_7 (C2V_112_447),
	.C2V_8 (C2V_112_487),
	.C2V_9 (C2V_112_571),
	.C2V_10 (C2V_112_585),
	.C2V_11 (C2V_112_658),
	.C2V_12 (C2V_112_704),
	.C2V_13 (C2V_112_873),
	.C2V_14 (C2V_112_945),
	.C2V_15 (C2V_112_981),
	.C2V_16 (C2V_112_1011),
	.C2V_17 (C2V_112_1086),
	.C2V_18 (C2V_112_1150),
	.C2V_19 (C2V_112_1263),
	.C2V_20 (C2V_112_1264),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU113 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_17_113),
	.V2C_2 (V2C_75_113),
	.V2C_3 (V2C_110_113),
	.V2C_4 (V2C_181_113),
	.V2C_5 (V2C_197_113),
	.V2C_6 (V2C_263_113),
	.V2C_7 (V2C_312_113),
	.V2C_8 (V2C_379_113),
	.V2C_9 (V2C_458_113),
	.V2C_10 (V2C_692_113),
	.V2C_11 (V2C_756_113),
	.V2C_12 (V2C_810_113),
	.V2C_13 (V2C_888_113),
	.V2C_14 (V2C_936_113),
	.V2C_15 (V2C_979_113),
	.V2C_16 (V2C_1031_113),
	.V2C_17 (V2C_1080_113),
	.V2C_18 (V2C_1128_113),
	.V2C_19 (V2C_1264_113),
	.V2C_20 (V2C_1265_113),
	.C2V_1 (C2V_113_17),
	.C2V_2 (C2V_113_75),
	.C2V_3 (C2V_113_110),
	.C2V_4 (C2V_113_181),
	.C2V_5 (C2V_113_197),
	.C2V_6 (C2V_113_263),
	.C2V_7 (C2V_113_312),
	.C2V_8 (C2V_113_379),
	.C2V_9 (C2V_113_458),
	.C2V_10 (C2V_113_692),
	.C2V_11 (C2V_113_756),
	.C2V_12 (C2V_113_810),
	.C2V_13 (C2V_113_888),
	.C2V_14 (C2V_113_936),
	.C2V_15 (C2V_113_979),
	.C2V_16 (C2V_113_1031),
	.C2V_17 (C2V_113_1080),
	.C2V_18 (C2V_113_1128),
	.C2V_19 (C2V_113_1264),
	.C2V_20 (C2V_113_1265),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU114 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_48_114),
	.V2C_2 (V2C_72_114),
	.V2C_3 (V2C_112_114),
	.V2C_4 (V2C_180_114),
	.V2C_5 (V2C_214_114),
	.V2C_6 (V2C_245_114),
	.V2C_7 (V2C_298_114),
	.V2C_8 (V2C_450_114),
	.V2C_9 (V2C_547_114),
	.V2C_10 (V2C_580_114),
	.V2C_11 (V2C_784_114),
	.V2C_12 (V2C_860_114),
	.V2C_13 (V2C_893_114),
	.V2C_14 (V2C_955_114),
	.V2C_15 (V2C_990_114),
	.V2C_16 (V2C_1009_114),
	.V2C_17 (V2C_1073_114),
	.V2C_18 (V2C_1123_114),
	.V2C_19 (V2C_1265_114),
	.V2C_20 (V2C_1266_114),
	.C2V_1 (C2V_114_48),
	.C2V_2 (C2V_114_72),
	.C2V_3 (C2V_114_112),
	.C2V_4 (C2V_114_180),
	.C2V_5 (C2V_114_214),
	.C2V_6 (C2V_114_245),
	.C2V_7 (C2V_114_298),
	.C2V_8 (C2V_114_450),
	.C2V_9 (C2V_114_547),
	.C2V_10 (C2V_114_580),
	.C2V_11 (C2V_114_784),
	.C2V_12 (C2V_114_860),
	.C2V_13 (C2V_114_893),
	.C2V_14 (C2V_114_955),
	.C2V_15 (C2V_114_990),
	.C2V_16 (C2V_114_1009),
	.C2V_17 (C2V_114_1073),
	.C2V_18 (C2V_114_1123),
	.C2V_19 (C2V_114_1265),
	.C2V_20 (C2V_114_1266),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU115 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_24_115),
	.V2C_2 (V2C_60_115),
	.V2C_3 (V2C_128_115),
	.V2C_4 (V2C_189_115),
	.V2C_5 (V2C_203_115),
	.V2C_6 (V2C_246_115),
	.V2C_7 (V2C_346_115),
	.V2C_8 (V2C_400_115),
	.V2C_9 (V2C_497_115),
	.V2C_10 (V2C_733_115),
	.V2C_11 (V2C_781_115),
	.V2C_12 (V2C_829_115),
	.V2C_13 (V2C_870_115),
	.V2C_14 (V2C_959_115),
	.V2C_15 (V2C_993_115),
	.V2C_16 (V2C_1032_115),
	.V2C_17 (V2C_1058_115),
	.V2C_18 (V2C_1117_115),
	.V2C_19 (V2C_1266_115),
	.V2C_20 (V2C_1267_115),
	.C2V_1 (C2V_115_24),
	.C2V_2 (C2V_115_60),
	.C2V_3 (C2V_115_128),
	.C2V_4 (C2V_115_189),
	.C2V_5 (C2V_115_203),
	.C2V_6 (C2V_115_246),
	.C2V_7 (C2V_115_346),
	.C2V_8 (C2V_115_400),
	.C2V_9 (C2V_115_497),
	.C2V_10 (C2V_115_733),
	.C2V_11 (C2V_115_781),
	.C2V_12 (C2V_115_829),
	.C2V_13 (C2V_115_870),
	.C2V_14 (C2V_115_959),
	.C2V_15 (C2V_115_993),
	.C2V_16 (C2V_115_1032),
	.C2V_17 (C2V_115_1058),
	.C2V_18 (C2V_115_1117),
	.C2V_19 (C2V_115_1266),
	.C2V_20 (C2V_115_1267),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU116 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_33_116),
	.V2C_2 (V2C_82_116),
	.V2C_3 (V2C_138_116),
	.V2C_4 (V2C_186_116),
	.V2C_5 (V2C_215_116),
	.V2C_6 (V2C_284_116),
	.V2C_7 (V2C_335_116),
	.V2C_8 (V2C_394_116),
	.V2C_9 (V2C_483_116),
	.V2C_10 (V2C_643_116),
	.V2C_11 (V2C_704_116),
	.V2C_12 (V2C_824_116),
	.V2C_13 (V2C_866_116),
	.V2C_14 (V2C_929_116),
	.V2C_15 (V2C_1008_116),
	.V2C_16 (V2C_1040_116),
	.V2C_17 (V2C_1059_116),
	.V2C_18 (V2C_1138_116),
	.V2C_19 (V2C_1267_116),
	.V2C_20 (V2C_1268_116),
	.C2V_1 (C2V_116_33),
	.C2V_2 (C2V_116_82),
	.C2V_3 (C2V_116_138),
	.C2V_4 (C2V_116_186),
	.C2V_5 (C2V_116_215),
	.C2V_6 (C2V_116_284),
	.C2V_7 (C2V_116_335),
	.C2V_8 (C2V_116_394),
	.C2V_9 (C2V_116_483),
	.C2V_10 (C2V_116_643),
	.C2V_11 (C2V_116_704),
	.C2V_12 (C2V_116_824),
	.C2V_13 (C2V_116_866),
	.C2V_14 (C2V_116_929),
	.C2V_15 (C2V_116_1008),
	.C2V_16 (C2V_116_1040),
	.C2V_17 (C2V_116_1059),
	.C2V_18 (C2V_116_1138),
	.C2V_19 (C2V_116_1267),
	.C2V_20 (C2V_116_1268),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU117 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_28_117),
	.V2C_2 (V2C_55_117),
	.V2C_3 (V2C_120_117),
	.V2C_4 (V2C_154_117),
	.V2C_5 (V2C_220_117),
	.V2C_6 (V2C_287_117),
	.V2C_7 (V2C_384_117),
	.V2C_8 (V2C_391_117),
	.V2C_9 (V2C_550_117),
	.V2C_10 (V2C_607_117),
	.V2C_11 (V2C_635_117),
	.V2C_12 (V2C_739_117),
	.V2C_13 (V2C_870_117),
	.V2C_14 (V2C_914_117),
	.V2C_15 (V2C_987_117),
	.V2C_16 (V2C_1047_117),
	.V2C_17 (V2C_1077_117),
	.V2C_18 (V2C_1122_117),
	.V2C_19 (V2C_1268_117),
	.V2C_20 (V2C_1269_117),
	.C2V_1 (C2V_117_28),
	.C2V_2 (C2V_117_55),
	.C2V_3 (C2V_117_120),
	.C2V_4 (C2V_117_154),
	.C2V_5 (C2V_117_220),
	.C2V_6 (C2V_117_287),
	.C2V_7 (C2V_117_384),
	.C2V_8 (C2V_117_391),
	.C2V_9 (C2V_117_550),
	.C2V_10 (C2V_117_607),
	.C2V_11 (C2V_117_635),
	.C2V_12 (C2V_117_739),
	.C2V_13 (C2V_117_870),
	.C2V_14 (C2V_117_914),
	.C2V_15 (C2V_117_987),
	.C2V_16 (C2V_117_1047),
	.C2V_17 (C2V_117_1077),
	.C2V_18 (C2V_117_1122),
	.C2V_19 (C2V_117_1268),
	.C2V_20 (C2V_117_1269),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU118 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_47_118),
	.V2C_2 (V2C_58_118),
	.V2C_3 (V2C_97_118),
	.V2C_4 (V2C_153_118),
	.V2C_5 (V2C_218_118),
	.V2C_6 (V2C_272_118),
	.V2C_7 (V2C_448_118),
	.V2C_8 (V2C_488_118),
	.V2C_9 (V2C_572_118),
	.V2C_10 (V2C_586_118),
	.V2C_11 (V2C_659_118),
	.V2C_12 (V2C_705_118),
	.V2C_13 (V2C_874_118),
	.V2C_14 (V2C_946_118),
	.V2C_15 (V2C_982_118),
	.V2C_16 (V2C_1012_118),
	.V2C_17 (V2C_1087_118),
	.V2C_18 (V2C_1151_118),
	.V2C_19 (V2C_1269_118),
	.V2C_20 (V2C_1270_118),
	.C2V_1 (C2V_118_47),
	.C2V_2 (C2V_118_58),
	.C2V_3 (C2V_118_97),
	.C2V_4 (C2V_118_153),
	.C2V_5 (C2V_118_218),
	.C2V_6 (C2V_118_272),
	.C2V_7 (C2V_118_448),
	.C2V_8 (C2V_118_488),
	.C2V_9 (C2V_118_572),
	.C2V_10 (C2V_118_586),
	.C2V_11 (C2V_118_659),
	.C2V_12 (C2V_118_705),
	.C2V_13 (C2V_118_874),
	.C2V_14 (C2V_118_946),
	.C2V_15 (C2V_118_982),
	.C2V_16 (C2V_118_1012),
	.C2V_17 (C2V_118_1087),
	.C2V_18 (C2V_118_1151),
	.C2V_19 (C2V_118_1269),
	.C2V_20 (C2V_118_1270),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU119 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_18_119),
	.V2C_2 (V2C_76_119),
	.V2C_3 (V2C_111_119),
	.V2C_4 (V2C_182_119),
	.V2C_5 (V2C_198_119),
	.V2C_6 (V2C_264_119),
	.V2C_7 (V2C_313_119),
	.V2C_8 (V2C_380_119),
	.V2C_9 (V2C_459_119),
	.V2C_10 (V2C_693_119),
	.V2C_11 (V2C_757_119),
	.V2C_12 (V2C_811_119),
	.V2C_13 (V2C_889_119),
	.V2C_14 (V2C_937_119),
	.V2C_15 (V2C_980_119),
	.V2C_16 (V2C_1032_119),
	.V2C_17 (V2C_1081_119),
	.V2C_18 (V2C_1129_119),
	.V2C_19 (V2C_1270_119),
	.V2C_20 (V2C_1271_119),
	.C2V_1 (C2V_119_18),
	.C2V_2 (C2V_119_76),
	.C2V_3 (C2V_119_111),
	.C2V_4 (C2V_119_182),
	.C2V_5 (C2V_119_198),
	.C2V_6 (C2V_119_264),
	.C2V_7 (C2V_119_313),
	.C2V_8 (C2V_119_380),
	.C2V_9 (C2V_119_459),
	.C2V_10 (C2V_119_693),
	.C2V_11 (C2V_119_757),
	.C2V_12 (C2V_119_811),
	.C2V_13 (C2V_119_889),
	.C2V_14 (C2V_119_937),
	.C2V_15 (C2V_119_980),
	.C2V_16 (C2V_119_1032),
	.C2V_17 (C2V_119_1081),
	.C2V_18 (C2V_119_1129),
	.C2V_19 (C2V_119_1270),
	.C2V_20 (C2V_119_1271),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU120 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_1_120),
	.V2C_2 (V2C_73_120),
	.V2C_3 (V2C_113_120),
	.V2C_4 (V2C_181_120),
	.V2C_5 (V2C_215_120),
	.V2C_6 (V2C_246_120),
	.V2C_7 (V2C_299_120),
	.V2C_8 (V2C_451_120),
	.V2C_9 (V2C_548_120),
	.V2C_10 (V2C_581_120),
	.V2C_11 (V2C_785_120),
	.V2C_12 (V2C_861_120),
	.V2C_13 (V2C_894_120),
	.V2C_14 (V2C_956_120),
	.V2C_15 (V2C_991_120),
	.V2C_16 (V2C_1010_120),
	.V2C_17 (V2C_1074_120),
	.V2C_18 (V2C_1124_120),
	.V2C_19 (V2C_1271_120),
	.V2C_20 (V2C_1272_120),
	.C2V_1 (C2V_120_1),
	.C2V_2 (C2V_120_73),
	.C2V_3 (C2V_120_113),
	.C2V_4 (C2V_120_181),
	.C2V_5 (C2V_120_215),
	.C2V_6 (C2V_120_246),
	.C2V_7 (C2V_120_299),
	.C2V_8 (C2V_120_451),
	.C2V_9 (C2V_120_548),
	.C2V_10 (C2V_120_581),
	.C2V_11 (C2V_120_785),
	.C2V_12 (C2V_120_861),
	.C2V_13 (C2V_120_894),
	.C2V_14 (C2V_120_956),
	.C2V_15 (C2V_120_991),
	.C2V_16 (C2V_120_1010),
	.C2V_17 (C2V_120_1074),
	.C2V_18 (C2V_120_1124),
	.C2V_19 (C2V_120_1271),
	.C2V_20 (C2V_120_1272),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU121 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_25_121),
	.V2C_2 (V2C_61_121),
	.V2C_3 (V2C_129_121),
	.V2C_4 (V2C_190_121),
	.V2C_5 (V2C_204_121),
	.V2C_6 (V2C_247_121),
	.V2C_7 (V2C_347_121),
	.V2C_8 (V2C_401_121),
	.V2C_9 (V2C_498_121),
	.V2C_10 (V2C_734_121),
	.V2C_11 (V2C_782_121),
	.V2C_12 (V2C_830_121),
	.V2C_13 (V2C_871_121),
	.V2C_14 (V2C_960_121),
	.V2C_15 (V2C_994_121),
	.V2C_16 (V2C_1033_121),
	.V2C_17 (V2C_1059_121),
	.V2C_18 (V2C_1118_121),
	.V2C_19 (V2C_1272_121),
	.V2C_20 (V2C_1273_121),
	.C2V_1 (C2V_121_25),
	.C2V_2 (C2V_121_61),
	.C2V_3 (C2V_121_129),
	.C2V_4 (C2V_121_190),
	.C2V_5 (C2V_121_204),
	.C2V_6 (C2V_121_247),
	.C2V_7 (C2V_121_347),
	.C2V_8 (C2V_121_401),
	.C2V_9 (C2V_121_498),
	.C2V_10 (C2V_121_734),
	.C2V_11 (C2V_121_782),
	.C2V_12 (C2V_121_830),
	.C2V_13 (C2V_121_871),
	.C2V_14 (C2V_121_960),
	.C2V_15 (C2V_121_994),
	.C2V_16 (C2V_121_1033),
	.C2V_17 (C2V_121_1059),
	.C2V_18 (C2V_121_1118),
	.C2V_19 (C2V_121_1272),
	.C2V_20 (C2V_121_1273),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU122 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_34_122),
	.V2C_2 (V2C_83_122),
	.V2C_3 (V2C_139_122),
	.V2C_4 (V2C_187_122),
	.V2C_5 (V2C_216_122),
	.V2C_6 (V2C_285_122),
	.V2C_7 (V2C_336_122),
	.V2C_8 (V2C_395_122),
	.V2C_9 (V2C_484_122),
	.V2C_10 (V2C_644_122),
	.V2C_11 (V2C_705_122),
	.V2C_12 (V2C_825_122),
	.V2C_13 (V2C_867_122),
	.V2C_14 (V2C_930_122),
	.V2C_15 (V2C_961_122),
	.V2C_16 (V2C_1041_122),
	.V2C_17 (V2C_1060_122),
	.V2C_18 (V2C_1139_122),
	.V2C_19 (V2C_1273_122),
	.V2C_20 (V2C_1274_122),
	.C2V_1 (C2V_122_34),
	.C2V_2 (C2V_122_83),
	.C2V_3 (C2V_122_139),
	.C2V_4 (C2V_122_187),
	.C2V_5 (C2V_122_216),
	.C2V_6 (C2V_122_285),
	.C2V_7 (C2V_122_336),
	.C2V_8 (C2V_122_395),
	.C2V_9 (C2V_122_484),
	.C2V_10 (C2V_122_644),
	.C2V_11 (C2V_122_705),
	.C2V_12 (C2V_122_825),
	.C2V_13 (C2V_122_867),
	.C2V_14 (C2V_122_930),
	.C2V_15 (C2V_122_961),
	.C2V_16 (C2V_122_1041),
	.C2V_17 (C2V_122_1060),
	.C2V_18 (C2V_122_1139),
	.C2V_19 (C2V_122_1273),
	.C2V_20 (C2V_122_1274),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU123 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_29_123),
	.V2C_2 (V2C_56_123),
	.V2C_3 (V2C_121_123),
	.V2C_4 (V2C_155_123),
	.V2C_5 (V2C_221_123),
	.V2C_6 (V2C_288_123),
	.V2C_7 (V2C_337_123),
	.V2C_8 (V2C_392_123),
	.V2C_9 (V2C_551_123),
	.V2C_10 (V2C_608_123),
	.V2C_11 (V2C_636_123),
	.V2C_12 (V2C_740_123),
	.V2C_13 (V2C_871_123),
	.V2C_14 (V2C_915_123),
	.V2C_15 (V2C_988_123),
	.V2C_16 (V2C_1048_123),
	.V2C_17 (V2C_1078_123),
	.V2C_18 (V2C_1123_123),
	.V2C_19 (V2C_1274_123),
	.V2C_20 (V2C_1275_123),
	.C2V_1 (C2V_123_29),
	.C2V_2 (C2V_123_56),
	.C2V_3 (C2V_123_121),
	.C2V_4 (C2V_123_155),
	.C2V_5 (C2V_123_221),
	.C2V_6 (C2V_123_288),
	.C2V_7 (C2V_123_337),
	.C2V_8 (C2V_123_392),
	.C2V_9 (C2V_123_551),
	.C2V_10 (C2V_123_608),
	.C2V_11 (C2V_123_636),
	.C2V_12 (C2V_123_740),
	.C2V_13 (C2V_123_871),
	.C2V_14 (C2V_123_915),
	.C2V_15 (C2V_123_988),
	.C2V_16 (C2V_123_1048),
	.C2V_17 (C2V_123_1078),
	.C2V_18 (C2V_123_1123),
	.C2V_19 (C2V_123_1274),
	.C2V_20 (C2V_123_1275),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU124 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_48_124),
	.V2C_2 (V2C_59_124),
	.V2C_3 (V2C_98_124),
	.V2C_4 (V2C_154_124),
	.V2C_5 (V2C_219_124),
	.V2C_6 (V2C_273_124),
	.V2C_7 (V2C_449_124),
	.V2C_8 (V2C_489_124),
	.V2C_9 (V2C_573_124),
	.V2C_10 (V2C_587_124),
	.V2C_11 (V2C_660_124),
	.V2C_12 (V2C_706_124),
	.V2C_13 (V2C_875_124),
	.V2C_14 (V2C_947_124),
	.V2C_15 (V2C_983_124),
	.V2C_16 (V2C_1013_124),
	.V2C_17 (V2C_1088_124),
	.V2C_18 (V2C_1152_124),
	.V2C_19 (V2C_1275_124),
	.V2C_20 (V2C_1276_124),
	.C2V_1 (C2V_124_48),
	.C2V_2 (C2V_124_59),
	.C2V_3 (C2V_124_98),
	.C2V_4 (C2V_124_154),
	.C2V_5 (C2V_124_219),
	.C2V_6 (C2V_124_273),
	.C2V_7 (C2V_124_449),
	.C2V_8 (C2V_124_489),
	.C2V_9 (C2V_124_573),
	.C2V_10 (C2V_124_587),
	.C2V_11 (C2V_124_660),
	.C2V_12 (C2V_124_706),
	.C2V_13 (C2V_124_875),
	.C2V_14 (C2V_124_947),
	.C2V_15 (C2V_124_983),
	.C2V_16 (C2V_124_1013),
	.C2V_17 (C2V_124_1088),
	.C2V_18 (C2V_124_1152),
	.C2V_19 (C2V_124_1275),
	.C2V_20 (C2V_124_1276),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU125 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_19_125),
	.V2C_2 (V2C_77_125),
	.V2C_3 (V2C_112_125),
	.V2C_4 (V2C_183_125),
	.V2C_5 (V2C_199_125),
	.V2C_6 (V2C_265_125),
	.V2C_7 (V2C_314_125),
	.V2C_8 (V2C_381_125),
	.V2C_9 (V2C_460_125),
	.V2C_10 (V2C_694_125),
	.V2C_11 (V2C_758_125),
	.V2C_12 (V2C_812_125),
	.V2C_13 (V2C_890_125),
	.V2C_14 (V2C_938_125),
	.V2C_15 (V2C_981_125),
	.V2C_16 (V2C_1033_125),
	.V2C_17 (V2C_1082_125),
	.V2C_18 (V2C_1130_125),
	.V2C_19 (V2C_1276_125),
	.V2C_20 (V2C_1277_125),
	.C2V_1 (C2V_125_19),
	.C2V_2 (C2V_125_77),
	.C2V_3 (C2V_125_112),
	.C2V_4 (C2V_125_183),
	.C2V_5 (C2V_125_199),
	.C2V_6 (C2V_125_265),
	.C2V_7 (C2V_125_314),
	.C2V_8 (C2V_125_381),
	.C2V_9 (C2V_125_460),
	.C2V_10 (C2V_125_694),
	.C2V_11 (C2V_125_758),
	.C2V_12 (C2V_125_812),
	.C2V_13 (C2V_125_890),
	.C2V_14 (C2V_125_938),
	.C2V_15 (C2V_125_981),
	.C2V_16 (C2V_125_1033),
	.C2V_17 (C2V_125_1082),
	.C2V_18 (C2V_125_1130),
	.C2V_19 (C2V_125_1276),
	.C2V_20 (C2V_125_1277),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU126 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_2_126),
	.V2C_2 (V2C_74_126),
	.V2C_3 (V2C_114_126),
	.V2C_4 (V2C_182_126),
	.V2C_5 (V2C_216_126),
	.V2C_6 (V2C_247_126),
	.V2C_7 (V2C_300_126),
	.V2C_8 (V2C_452_126),
	.V2C_9 (V2C_549_126),
	.V2C_10 (V2C_582_126),
	.V2C_11 (V2C_786_126),
	.V2C_12 (V2C_862_126),
	.V2C_13 (V2C_895_126),
	.V2C_14 (V2C_957_126),
	.V2C_15 (V2C_992_126),
	.V2C_16 (V2C_1011_126),
	.V2C_17 (V2C_1075_126),
	.V2C_18 (V2C_1125_126),
	.V2C_19 (V2C_1277_126),
	.V2C_20 (V2C_1278_126),
	.C2V_1 (C2V_126_2),
	.C2V_2 (C2V_126_74),
	.C2V_3 (C2V_126_114),
	.C2V_4 (C2V_126_182),
	.C2V_5 (C2V_126_216),
	.C2V_6 (C2V_126_247),
	.C2V_7 (C2V_126_300),
	.C2V_8 (C2V_126_452),
	.C2V_9 (C2V_126_549),
	.C2V_10 (C2V_126_582),
	.C2V_11 (C2V_126_786),
	.C2V_12 (C2V_126_862),
	.C2V_13 (C2V_126_895),
	.C2V_14 (C2V_126_957),
	.C2V_15 (C2V_126_992),
	.C2V_16 (C2V_126_1011),
	.C2V_17 (C2V_126_1075),
	.C2V_18 (C2V_126_1125),
	.C2V_19 (C2V_126_1277),
	.C2V_20 (C2V_126_1278),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU127 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_26_127),
	.V2C_2 (V2C_62_127),
	.V2C_3 (V2C_130_127),
	.V2C_4 (V2C_191_127),
	.V2C_5 (V2C_205_127),
	.V2C_6 (V2C_248_127),
	.V2C_7 (V2C_348_127),
	.V2C_8 (V2C_402_127),
	.V2C_9 (V2C_499_127),
	.V2C_10 (V2C_735_127),
	.V2C_11 (V2C_783_127),
	.V2C_12 (V2C_831_127),
	.V2C_13 (V2C_872_127),
	.V2C_14 (V2C_913_127),
	.V2C_15 (V2C_995_127),
	.V2C_16 (V2C_1034_127),
	.V2C_17 (V2C_1060_127),
	.V2C_18 (V2C_1119_127),
	.V2C_19 (V2C_1278_127),
	.V2C_20 (V2C_1279_127),
	.C2V_1 (C2V_127_26),
	.C2V_2 (C2V_127_62),
	.C2V_3 (C2V_127_130),
	.C2V_4 (C2V_127_191),
	.C2V_5 (C2V_127_205),
	.C2V_6 (C2V_127_248),
	.C2V_7 (C2V_127_348),
	.C2V_8 (C2V_127_402),
	.C2V_9 (C2V_127_499),
	.C2V_10 (C2V_127_735),
	.C2V_11 (C2V_127_783),
	.C2V_12 (C2V_127_831),
	.C2V_13 (C2V_127_872),
	.C2V_14 (C2V_127_913),
	.C2V_15 (C2V_127_995),
	.C2V_16 (C2V_127_1034),
	.C2V_17 (C2V_127_1060),
	.C2V_18 (C2V_127_1119),
	.C2V_19 (C2V_127_1278),
	.C2V_20 (C2V_127_1279),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU128 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_35_128),
	.V2C_2 (V2C_84_128),
	.V2C_3 (V2C_140_128),
	.V2C_4 (V2C_188_128),
	.V2C_5 (V2C_217_128),
	.V2C_6 (V2C_286_128),
	.V2C_7 (V2C_289_128),
	.V2C_8 (V2C_396_128),
	.V2C_9 (V2C_485_128),
	.V2C_10 (V2C_645_128),
	.V2C_11 (V2C_706_128),
	.V2C_12 (V2C_826_128),
	.V2C_13 (V2C_868_128),
	.V2C_14 (V2C_931_128),
	.V2C_15 (V2C_962_128),
	.V2C_16 (V2C_1042_128),
	.V2C_17 (V2C_1061_128),
	.V2C_18 (V2C_1140_128),
	.V2C_19 (V2C_1279_128),
	.V2C_20 (V2C_1280_128),
	.C2V_1 (C2V_128_35),
	.C2V_2 (C2V_128_84),
	.C2V_3 (C2V_128_140),
	.C2V_4 (C2V_128_188),
	.C2V_5 (C2V_128_217),
	.C2V_6 (C2V_128_286),
	.C2V_7 (C2V_128_289),
	.C2V_8 (C2V_128_396),
	.C2V_9 (C2V_128_485),
	.C2V_10 (C2V_128_645),
	.C2V_11 (C2V_128_706),
	.C2V_12 (C2V_128_826),
	.C2V_13 (C2V_128_868),
	.C2V_14 (C2V_128_931),
	.C2V_15 (C2V_128_962),
	.C2V_16 (C2V_128_1042),
	.C2V_17 (C2V_128_1061),
	.C2V_18 (C2V_128_1140),
	.C2V_19 (C2V_128_1279),
	.C2V_20 (C2V_128_1280),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU129 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_30_129),
	.V2C_2 (V2C_57_129),
	.V2C_3 (V2C_122_129),
	.V2C_4 (V2C_156_129),
	.V2C_5 (V2C_222_129),
	.V2C_6 (V2C_241_129),
	.V2C_7 (V2C_338_129),
	.V2C_8 (V2C_393_129),
	.V2C_9 (V2C_552_129),
	.V2C_10 (V2C_609_129),
	.V2C_11 (V2C_637_129),
	.V2C_12 (V2C_741_129),
	.V2C_13 (V2C_872_129),
	.V2C_14 (V2C_916_129),
	.V2C_15 (V2C_989_129),
	.V2C_16 (V2C_1049_129),
	.V2C_17 (V2C_1079_129),
	.V2C_18 (V2C_1124_129),
	.V2C_19 (V2C_1280_129),
	.V2C_20 (V2C_1281_129),
	.C2V_1 (C2V_129_30),
	.C2V_2 (C2V_129_57),
	.C2V_3 (C2V_129_122),
	.C2V_4 (C2V_129_156),
	.C2V_5 (C2V_129_222),
	.C2V_6 (C2V_129_241),
	.C2V_7 (C2V_129_338),
	.C2V_8 (C2V_129_393),
	.C2V_9 (C2V_129_552),
	.C2V_10 (C2V_129_609),
	.C2V_11 (C2V_129_637),
	.C2V_12 (C2V_129_741),
	.C2V_13 (C2V_129_872),
	.C2V_14 (C2V_129_916),
	.C2V_15 (C2V_129_989),
	.C2V_16 (C2V_129_1049),
	.C2V_17 (C2V_129_1079),
	.C2V_18 (C2V_129_1124),
	.C2V_19 (C2V_129_1280),
	.C2V_20 (C2V_129_1281),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU130 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_1_130),
	.V2C_2 (V2C_60_130),
	.V2C_3 (V2C_99_130),
	.V2C_4 (V2C_155_130),
	.V2C_5 (V2C_220_130),
	.V2C_6 (V2C_274_130),
	.V2C_7 (V2C_450_130),
	.V2C_8 (V2C_490_130),
	.V2C_9 (V2C_574_130),
	.V2C_10 (V2C_588_130),
	.V2C_11 (V2C_661_130),
	.V2C_12 (V2C_707_130),
	.V2C_13 (V2C_876_130),
	.V2C_14 (V2C_948_130),
	.V2C_15 (V2C_984_130),
	.V2C_16 (V2C_1014_130),
	.V2C_17 (V2C_1089_130),
	.V2C_18 (V2C_1105_130),
	.V2C_19 (V2C_1281_130),
	.V2C_20 (V2C_1282_130),
	.C2V_1 (C2V_130_1),
	.C2V_2 (C2V_130_60),
	.C2V_3 (C2V_130_99),
	.C2V_4 (C2V_130_155),
	.C2V_5 (C2V_130_220),
	.C2V_6 (C2V_130_274),
	.C2V_7 (C2V_130_450),
	.C2V_8 (C2V_130_490),
	.C2V_9 (C2V_130_574),
	.C2V_10 (C2V_130_588),
	.C2V_11 (C2V_130_661),
	.C2V_12 (C2V_130_707),
	.C2V_13 (C2V_130_876),
	.C2V_14 (C2V_130_948),
	.C2V_15 (C2V_130_984),
	.C2V_16 (C2V_130_1014),
	.C2V_17 (C2V_130_1089),
	.C2V_18 (C2V_130_1105),
	.C2V_19 (C2V_130_1281),
	.C2V_20 (C2V_130_1282),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU131 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_20_131),
	.V2C_2 (V2C_78_131),
	.V2C_3 (V2C_113_131),
	.V2C_4 (V2C_184_131),
	.V2C_5 (V2C_200_131),
	.V2C_6 (V2C_266_131),
	.V2C_7 (V2C_315_131),
	.V2C_8 (V2C_382_131),
	.V2C_9 (V2C_461_131),
	.V2C_10 (V2C_695_131),
	.V2C_11 (V2C_759_131),
	.V2C_12 (V2C_813_131),
	.V2C_13 (V2C_891_131),
	.V2C_14 (V2C_939_131),
	.V2C_15 (V2C_982_131),
	.V2C_16 (V2C_1034_131),
	.V2C_17 (V2C_1083_131),
	.V2C_18 (V2C_1131_131),
	.V2C_19 (V2C_1282_131),
	.V2C_20 (V2C_1283_131),
	.C2V_1 (C2V_131_20),
	.C2V_2 (C2V_131_78),
	.C2V_3 (C2V_131_113),
	.C2V_4 (C2V_131_184),
	.C2V_5 (C2V_131_200),
	.C2V_6 (C2V_131_266),
	.C2V_7 (C2V_131_315),
	.C2V_8 (C2V_131_382),
	.C2V_9 (C2V_131_461),
	.C2V_10 (C2V_131_695),
	.C2V_11 (C2V_131_759),
	.C2V_12 (C2V_131_813),
	.C2V_13 (C2V_131_891),
	.C2V_14 (C2V_131_939),
	.C2V_15 (C2V_131_982),
	.C2V_16 (C2V_131_1034),
	.C2V_17 (C2V_131_1083),
	.C2V_18 (C2V_131_1131),
	.C2V_19 (C2V_131_1282),
	.C2V_20 (C2V_131_1283),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU132 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_3_132),
	.V2C_2 (V2C_75_132),
	.V2C_3 (V2C_115_132),
	.V2C_4 (V2C_183_132),
	.V2C_5 (V2C_217_132),
	.V2C_6 (V2C_248_132),
	.V2C_7 (V2C_301_132),
	.V2C_8 (V2C_453_132),
	.V2C_9 (V2C_550_132),
	.V2C_10 (V2C_583_132),
	.V2C_11 (V2C_787_132),
	.V2C_12 (V2C_863_132),
	.V2C_13 (V2C_896_132),
	.V2C_14 (V2C_958_132),
	.V2C_15 (V2C_993_132),
	.V2C_16 (V2C_1012_132),
	.V2C_17 (V2C_1076_132),
	.V2C_18 (V2C_1126_132),
	.V2C_19 (V2C_1283_132),
	.V2C_20 (V2C_1284_132),
	.C2V_1 (C2V_132_3),
	.C2V_2 (C2V_132_75),
	.C2V_3 (C2V_132_115),
	.C2V_4 (C2V_132_183),
	.C2V_5 (C2V_132_217),
	.C2V_6 (C2V_132_248),
	.C2V_7 (C2V_132_301),
	.C2V_8 (C2V_132_453),
	.C2V_9 (C2V_132_550),
	.C2V_10 (C2V_132_583),
	.C2V_11 (C2V_132_787),
	.C2V_12 (C2V_132_863),
	.C2V_13 (C2V_132_896),
	.C2V_14 (C2V_132_958),
	.C2V_15 (C2V_132_993),
	.C2V_16 (C2V_132_1012),
	.C2V_17 (C2V_132_1076),
	.C2V_18 (C2V_132_1126),
	.C2V_19 (C2V_132_1283),
	.C2V_20 (C2V_132_1284),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU133 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_27_133),
	.V2C_2 (V2C_63_133),
	.V2C_3 (V2C_131_133),
	.V2C_4 (V2C_192_133),
	.V2C_5 (V2C_206_133),
	.V2C_6 (V2C_249_133),
	.V2C_7 (V2C_349_133),
	.V2C_8 (V2C_403_133),
	.V2C_9 (V2C_500_133),
	.V2C_10 (V2C_736_133),
	.V2C_11 (V2C_784_133),
	.V2C_12 (V2C_832_133),
	.V2C_13 (V2C_873_133),
	.V2C_14 (V2C_914_133),
	.V2C_15 (V2C_996_133),
	.V2C_16 (V2C_1035_133),
	.V2C_17 (V2C_1061_133),
	.V2C_18 (V2C_1120_133),
	.V2C_19 (V2C_1284_133),
	.V2C_20 (V2C_1285_133),
	.C2V_1 (C2V_133_27),
	.C2V_2 (C2V_133_63),
	.C2V_3 (C2V_133_131),
	.C2V_4 (C2V_133_192),
	.C2V_5 (C2V_133_206),
	.C2V_6 (C2V_133_249),
	.C2V_7 (C2V_133_349),
	.C2V_8 (C2V_133_403),
	.C2V_9 (C2V_133_500),
	.C2V_10 (C2V_133_736),
	.C2V_11 (C2V_133_784),
	.C2V_12 (C2V_133_832),
	.C2V_13 (C2V_133_873),
	.C2V_14 (C2V_133_914),
	.C2V_15 (C2V_133_996),
	.C2V_16 (C2V_133_1035),
	.C2V_17 (C2V_133_1061),
	.C2V_18 (C2V_133_1120),
	.C2V_19 (C2V_133_1284),
	.C2V_20 (C2V_133_1285),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU134 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_36_134),
	.V2C_2 (V2C_85_134),
	.V2C_3 (V2C_141_134),
	.V2C_4 (V2C_189_134),
	.V2C_5 (V2C_218_134),
	.V2C_6 (V2C_287_134),
	.V2C_7 (V2C_290_134),
	.V2C_8 (V2C_397_134),
	.V2C_9 (V2C_486_134),
	.V2C_10 (V2C_646_134),
	.V2C_11 (V2C_707_134),
	.V2C_12 (V2C_827_134),
	.V2C_13 (V2C_869_134),
	.V2C_14 (V2C_932_134),
	.V2C_15 (V2C_963_134),
	.V2C_16 (V2C_1043_134),
	.V2C_17 (V2C_1062_134),
	.V2C_18 (V2C_1141_134),
	.V2C_19 (V2C_1285_134),
	.V2C_20 (V2C_1286_134),
	.C2V_1 (C2V_134_36),
	.C2V_2 (C2V_134_85),
	.C2V_3 (C2V_134_141),
	.C2V_4 (C2V_134_189),
	.C2V_5 (C2V_134_218),
	.C2V_6 (C2V_134_287),
	.C2V_7 (C2V_134_290),
	.C2V_8 (C2V_134_397),
	.C2V_9 (C2V_134_486),
	.C2V_10 (C2V_134_646),
	.C2V_11 (C2V_134_707),
	.C2V_12 (C2V_134_827),
	.C2V_13 (C2V_134_869),
	.C2V_14 (C2V_134_932),
	.C2V_15 (C2V_134_963),
	.C2V_16 (C2V_134_1043),
	.C2V_17 (C2V_134_1062),
	.C2V_18 (C2V_134_1141),
	.C2V_19 (C2V_134_1285),
	.C2V_20 (C2V_134_1286),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU135 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_31_135),
	.V2C_2 (V2C_58_135),
	.V2C_3 (V2C_123_135),
	.V2C_4 (V2C_157_135),
	.V2C_5 (V2C_223_135),
	.V2C_6 (V2C_242_135),
	.V2C_7 (V2C_339_135),
	.V2C_8 (V2C_394_135),
	.V2C_9 (V2C_553_135),
	.V2C_10 (V2C_610_135),
	.V2C_11 (V2C_638_135),
	.V2C_12 (V2C_742_135),
	.V2C_13 (V2C_873_135),
	.V2C_14 (V2C_917_135),
	.V2C_15 (V2C_990_135),
	.V2C_16 (V2C_1050_135),
	.V2C_17 (V2C_1080_135),
	.V2C_18 (V2C_1125_135),
	.V2C_19 (V2C_1286_135),
	.V2C_20 (V2C_1287_135),
	.C2V_1 (C2V_135_31),
	.C2V_2 (C2V_135_58),
	.C2V_3 (C2V_135_123),
	.C2V_4 (C2V_135_157),
	.C2V_5 (C2V_135_223),
	.C2V_6 (C2V_135_242),
	.C2V_7 (C2V_135_339),
	.C2V_8 (C2V_135_394),
	.C2V_9 (C2V_135_553),
	.C2V_10 (C2V_135_610),
	.C2V_11 (C2V_135_638),
	.C2V_12 (C2V_135_742),
	.C2V_13 (C2V_135_873),
	.C2V_14 (C2V_135_917),
	.C2V_15 (C2V_135_990),
	.C2V_16 (C2V_135_1050),
	.C2V_17 (C2V_135_1080),
	.C2V_18 (C2V_135_1125),
	.C2V_19 (C2V_135_1286),
	.C2V_20 (C2V_135_1287),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU136 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_2_136),
	.V2C_2 (V2C_61_136),
	.V2C_3 (V2C_100_136),
	.V2C_4 (V2C_156_136),
	.V2C_5 (V2C_221_136),
	.V2C_6 (V2C_275_136),
	.V2C_7 (V2C_451_136),
	.V2C_8 (V2C_491_136),
	.V2C_9 (V2C_575_136),
	.V2C_10 (V2C_589_136),
	.V2C_11 (V2C_662_136),
	.V2C_12 (V2C_708_136),
	.V2C_13 (V2C_877_136),
	.V2C_14 (V2C_949_136),
	.V2C_15 (V2C_985_136),
	.V2C_16 (V2C_1015_136),
	.V2C_17 (V2C_1090_136),
	.V2C_18 (V2C_1106_136),
	.V2C_19 (V2C_1287_136),
	.V2C_20 (V2C_1288_136),
	.C2V_1 (C2V_136_2),
	.C2V_2 (C2V_136_61),
	.C2V_3 (C2V_136_100),
	.C2V_4 (C2V_136_156),
	.C2V_5 (C2V_136_221),
	.C2V_6 (C2V_136_275),
	.C2V_7 (C2V_136_451),
	.C2V_8 (C2V_136_491),
	.C2V_9 (C2V_136_575),
	.C2V_10 (C2V_136_589),
	.C2V_11 (C2V_136_662),
	.C2V_12 (C2V_136_708),
	.C2V_13 (C2V_136_877),
	.C2V_14 (C2V_136_949),
	.C2V_15 (C2V_136_985),
	.C2V_16 (C2V_136_1015),
	.C2V_17 (C2V_136_1090),
	.C2V_18 (C2V_136_1106),
	.C2V_19 (C2V_136_1287),
	.C2V_20 (C2V_136_1288),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU137 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_21_137),
	.V2C_2 (V2C_79_137),
	.V2C_3 (V2C_114_137),
	.V2C_4 (V2C_185_137),
	.V2C_5 (V2C_201_137),
	.V2C_6 (V2C_267_137),
	.V2C_7 (V2C_316_137),
	.V2C_8 (V2C_383_137),
	.V2C_9 (V2C_462_137),
	.V2C_10 (V2C_696_137),
	.V2C_11 (V2C_760_137),
	.V2C_12 (V2C_814_137),
	.V2C_13 (V2C_892_137),
	.V2C_14 (V2C_940_137),
	.V2C_15 (V2C_983_137),
	.V2C_16 (V2C_1035_137),
	.V2C_17 (V2C_1084_137),
	.V2C_18 (V2C_1132_137),
	.V2C_19 (V2C_1288_137),
	.V2C_20 (V2C_1289_137),
	.C2V_1 (C2V_137_21),
	.C2V_2 (C2V_137_79),
	.C2V_3 (C2V_137_114),
	.C2V_4 (C2V_137_185),
	.C2V_5 (C2V_137_201),
	.C2V_6 (C2V_137_267),
	.C2V_7 (C2V_137_316),
	.C2V_8 (C2V_137_383),
	.C2V_9 (C2V_137_462),
	.C2V_10 (C2V_137_696),
	.C2V_11 (C2V_137_760),
	.C2V_12 (C2V_137_814),
	.C2V_13 (C2V_137_892),
	.C2V_14 (C2V_137_940),
	.C2V_15 (C2V_137_983),
	.C2V_16 (C2V_137_1035),
	.C2V_17 (C2V_137_1084),
	.C2V_18 (C2V_137_1132),
	.C2V_19 (C2V_137_1288),
	.C2V_20 (C2V_137_1289),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU138 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_4_138),
	.V2C_2 (V2C_76_138),
	.V2C_3 (V2C_116_138),
	.V2C_4 (V2C_184_138),
	.V2C_5 (V2C_218_138),
	.V2C_6 (V2C_249_138),
	.V2C_7 (V2C_302_138),
	.V2C_8 (V2C_454_138),
	.V2C_9 (V2C_551_138),
	.V2C_10 (V2C_584_138),
	.V2C_11 (V2C_788_138),
	.V2C_12 (V2C_864_138),
	.V2C_13 (V2C_897_138),
	.V2C_14 (V2C_959_138),
	.V2C_15 (V2C_994_138),
	.V2C_16 (V2C_1013_138),
	.V2C_17 (V2C_1077_138),
	.V2C_18 (V2C_1127_138),
	.V2C_19 (V2C_1289_138),
	.V2C_20 (V2C_1290_138),
	.C2V_1 (C2V_138_4),
	.C2V_2 (C2V_138_76),
	.C2V_3 (C2V_138_116),
	.C2V_4 (C2V_138_184),
	.C2V_5 (C2V_138_218),
	.C2V_6 (C2V_138_249),
	.C2V_7 (C2V_138_302),
	.C2V_8 (C2V_138_454),
	.C2V_9 (C2V_138_551),
	.C2V_10 (C2V_138_584),
	.C2V_11 (C2V_138_788),
	.C2V_12 (C2V_138_864),
	.C2V_13 (C2V_138_897),
	.C2V_14 (C2V_138_959),
	.C2V_15 (C2V_138_994),
	.C2V_16 (C2V_138_1013),
	.C2V_17 (C2V_138_1077),
	.C2V_18 (C2V_138_1127),
	.C2V_19 (C2V_138_1289),
	.C2V_20 (C2V_138_1290),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU139 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_28_139),
	.V2C_2 (V2C_64_139),
	.V2C_3 (V2C_132_139),
	.V2C_4 (V2C_145_139),
	.V2C_5 (V2C_207_139),
	.V2C_6 (V2C_250_139),
	.V2C_7 (V2C_350_139),
	.V2C_8 (V2C_404_139),
	.V2C_9 (V2C_501_139),
	.V2C_10 (V2C_737_139),
	.V2C_11 (V2C_785_139),
	.V2C_12 (V2C_833_139),
	.V2C_13 (V2C_874_139),
	.V2C_14 (V2C_915_139),
	.V2C_15 (V2C_997_139),
	.V2C_16 (V2C_1036_139),
	.V2C_17 (V2C_1062_139),
	.V2C_18 (V2C_1121_139),
	.V2C_19 (V2C_1290_139),
	.V2C_20 (V2C_1291_139),
	.C2V_1 (C2V_139_28),
	.C2V_2 (C2V_139_64),
	.C2V_3 (C2V_139_132),
	.C2V_4 (C2V_139_145),
	.C2V_5 (C2V_139_207),
	.C2V_6 (C2V_139_250),
	.C2V_7 (C2V_139_350),
	.C2V_8 (C2V_139_404),
	.C2V_9 (C2V_139_501),
	.C2V_10 (C2V_139_737),
	.C2V_11 (C2V_139_785),
	.C2V_12 (C2V_139_833),
	.C2V_13 (C2V_139_874),
	.C2V_14 (C2V_139_915),
	.C2V_15 (C2V_139_997),
	.C2V_16 (C2V_139_1036),
	.C2V_17 (C2V_139_1062),
	.C2V_18 (C2V_139_1121),
	.C2V_19 (C2V_139_1290),
	.C2V_20 (C2V_139_1291),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU140 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_37_140),
	.V2C_2 (V2C_86_140),
	.V2C_3 (V2C_142_140),
	.V2C_4 (V2C_190_140),
	.V2C_5 (V2C_219_140),
	.V2C_6 (V2C_288_140),
	.V2C_7 (V2C_291_140),
	.V2C_8 (V2C_398_140),
	.V2C_9 (V2C_487_140),
	.V2C_10 (V2C_647_140),
	.V2C_11 (V2C_708_140),
	.V2C_12 (V2C_828_140),
	.V2C_13 (V2C_870_140),
	.V2C_14 (V2C_933_140),
	.V2C_15 (V2C_964_140),
	.V2C_16 (V2C_1044_140),
	.V2C_17 (V2C_1063_140),
	.V2C_18 (V2C_1142_140),
	.V2C_19 (V2C_1291_140),
	.V2C_20 (V2C_1292_140),
	.C2V_1 (C2V_140_37),
	.C2V_2 (C2V_140_86),
	.C2V_3 (C2V_140_142),
	.C2V_4 (C2V_140_190),
	.C2V_5 (C2V_140_219),
	.C2V_6 (C2V_140_288),
	.C2V_7 (C2V_140_291),
	.C2V_8 (C2V_140_398),
	.C2V_9 (C2V_140_487),
	.C2V_10 (C2V_140_647),
	.C2V_11 (C2V_140_708),
	.C2V_12 (C2V_140_828),
	.C2V_13 (C2V_140_870),
	.C2V_14 (C2V_140_933),
	.C2V_15 (C2V_140_964),
	.C2V_16 (C2V_140_1044),
	.C2V_17 (C2V_140_1063),
	.C2V_18 (C2V_140_1142),
	.C2V_19 (C2V_140_1291),
	.C2V_20 (C2V_140_1292),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU141 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_32_141),
	.V2C_2 (V2C_59_141),
	.V2C_3 (V2C_124_141),
	.V2C_4 (V2C_158_141),
	.V2C_5 (V2C_224_141),
	.V2C_6 (V2C_243_141),
	.V2C_7 (V2C_340_141),
	.V2C_8 (V2C_395_141),
	.V2C_9 (V2C_554_141),
	.V2C_10 (V2C_611_141),
	.V2C_11 (V2C_639_141),
	.V2C_12 (V2C_743_141),
	.V2C_13 (V2C_874_141),
	.V2C_14 (V2C_918_141),
	.V2C_15 (V2C_991_141),
	.V2C_16 (V2C_1051_141),
	.V2C_17 (V2C_1081_141),
	.V2C_18 (V2C_1126_141),
	.V2C_19 (V2C_1292_141),
	.V2C_20 (V2C_1293_141),
	.C2V_1 (C2V_141_32),
	.C2V_2 (C2V_141_59),
	.C2V_3 (C2V_141_124),
	.C2V_4 (C2V_141_158),
	.C2V_5 (C2V_141_224),
	.C2V_6 (C2V_141_243),
	.C2V_7 (C2V_141_340),
	.C2V_8 (C2V_141_395),
	.C2V_9 (C2V_141_554),
	.C2V_10 (C2V_141_611),
	.C2V_11 (C2V_141_639),
	.C2V_12 (C2V_141_743),
	.C2V_13 (C2V_141_874),
	.C2V_14 (C2V_141_918),
	.C2V_15 (C2V_141_991),
	.C2V_16 (C2V_141_1051),
	.C2V_17 (C2V_141_1081),
	.C2V_18 (C2V_141_1126),
	.C2V_19 (C2V_141_1292),
	.C2V_20 (C2V_141_1293),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU142 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_3_142),
	.V2C_2 (V2C_62_142),
	.V2C_3 (V2C_101_142),
	.V2C_4 (V2C_157_142),
	.V2C_5 (V2C_222_142),
	.V2C_6 (V2C_276_142),
	.V2C_7 (V2C_452_142),
	.V2C_8 (V2C_492_142),
	.V2C_9 (V2C_576_142),
	.V2C_10 (V2C_590_142),
	.V2C_11 (V2C_663_142),
	.V2C_12 (V2C_709_142),
	.V2C_13 (V2C_878_142),
	.V2C_14 (V2C_950_142),
	.V2C_15 (V2C_986_142),
	.V2C_16 (V2C_1016_142),
	.V2C_17 (V2C_1091_142),
	.V2C_18 (V2C_1107_142),
	.V2C_19 (V2C_1293_142),
	.V2C_20 (V2C_1294_142),
	.C2V_1 (C2V_142_3),
	.C2V_2 (C2V_142_62),
	.C2V_3 (C2V_142_101),
	.C2V_4 (C2V_142_157),
	.C2V_5 (C2V_142_222),
	.C2V_6 (C2V_142_276),
	.C2V_7 (C2V_142_452),
	.C2V_8 (C2V_142_492),
	.C2V_9 (C2V_142_576),
	.C2V_10 (C2V_142_590),
	.C2V_11 (C2V_142_663),
	.C2V_12 (C2V_142_709),
	.C2V_13 (C2V_142_878),
	.C2V_14 (C2V_142_950),
	.C2V_15 (C2V_142_986),
	.C2V_16 (C2V_142_1016),
	.C2V_17 (C2V_142_1091),
	.C2V_18 (C2V_142_1107),
	.C2V_19 (C2V_142_1293),
	.C2V_20 (C2V_142_1294),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU143 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_22_143),
	.V2C_2 (V2C_80_143),
	.V2C_3 (V2C_115_143),
	.V2C_4 (V2C_186_143),
	.V2C_5 (V2C_202_143),
	.V2C_6 (V2C_268_143),
	.V2C_7 (V2C_317_143),
	.V2C_8 (V2C_384_143),
	.V2C_9 (V2C_463_143),
	.V2C_10 (V2C_697_143),
	.V2C_11 (V2C_761_143),
	.V2C_12 (V2C_815_143),
	.V2C_13 (V2C_893_143),
	.V2C_14 (V2C_941_143),
	.V2C_15 (V2C_984_143),
	.V2C_16 (V2C_1036_143),
	.V2C_17 (V2C_1085_143),
	.V2C_18 (V2C_1133_143),
	.V2C_19 (V2C_1294_143),
	.V2C_20 (V2C_1295_143),
	.C2V_1 (C2V_143_22),
	.C2V_2 (C2V_143_80),
	.C2V_3 (C2V_143_115),
	.C2V_4 (C2V_143_186),
	.C2V_5 (C2V_143_202),
	.C2V_6 (C2V_143_268),
	.C2V_7 (C2V_143_317),
	.C2V_8 (C2V_143_384),
	.C2V_9 (C2V_143_463),
	.C2V_10 (C2V_143_697),
	.C2V_11 (C2V_143_761),
	.C2V_12 (C2V_143_815),
	.C2V_13 (C2V_143_893),
	.C2V_14 (C2V_143_941),
	.C2V_15 (C2V_143_984),
	.C2V_16 (C2V_143_1036),
	.C2V_17 (C2V_143_1085),
	.C2V_18 (C2V_143_1133),
	.C2V_19 (C2V_143_1294),
	.C2V_20 (C2V_143_1295),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU144 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_5_144),
	.V2C_2 (V2C_77_144),
	.V2C_3 (V2C_117_144),
	.V2C_4 (V2C_185_144),
	.V2C_5 (V2C_219_144),
	.V2C_6 (V2C_250_144),
	.V2C_7 (V2C_303_144),
	.V2C_8 (V2C_455_144),
	.V2C_9 (V2C_552_144),
	.V2C_10 (V2C_585_144),
	.V2C_11 (V2C_789_144),
	.V2C_12 (V2C_817_144),
	.V2C_13 (V2C_898_144),
	.V2C_14 (V2C_960_144),
	.V2C_15 (V2C_995_144),
	.V2C_16 (V2C_1014_144),
	.V2C_17 (V2C_1078_144),
	.V2C_18 (V2C_1128_144),
	.V2C_19 (V2C_1295_144),
	.V2C_20 (V2C_1296_144),
	.C2V_1 (C2V_144_5),
	.C2V_2 (C2V_144_77),
	.C2V_3 (C2V_144_117),
	.C2V_4 (C2V_144_185),
	.C2V_5 (C2V_144_219),
	.C2V_6 (C2V_144_250),
	.C2V_7 (C2V_144_303),
	.C2V_8 (C2V_144_455),
	.C2V_9 (C2V_144_552),
	.C2V_10 (C2V_144_585),
	.C2V_11 (C2V_144_789),
	.C2V_12 (C2V_144_817),
	.C2V_13 (C2V_144_898),
	.C2V_14 (C2V_144_960),
	.C2V_15 (C2V_144_995),
	.C2V_16 (C2V_144_1014),
	.C2V_17 (C2V_144_1078),
	.C2V_18 (C2V_144_1128),
	.C2V_19 (C2V_144_1295),
	.C2V_20 (C2V_144_1296),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU145 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_29_145),
	.V2C_2 (V2C_65_145),
	.V2C_3 (V2C_133_145),
	.V2C_4 (V2C_146_145),
	.V2C_5 (V2C_208_145),
	.V2C_6 (V2C_251_145),
	.V2C_7 (V2C_351_145),
	.V2C_8 (V2C_405_145),
	.V2C_9 (V2C_502_145),
	.V2C_10 (V2C_738_145),
	.V2C_11 (V2C_786_145),
	.V2C_12 (V2C_834_145),
	.V2C_13 (V2C_875_145),
	.V2C_14 (V2C_916_145),
	.V2C_15 (V2C_998_145),
	.V2C_16 (V2C_1037_145),
	.V2C_17 (V2C_1063_145),
	.V2C_18 (V2C_1122_145),
	.V2C_19 (V2C_1296_145),
	.V2C_20 (V2C_1297_145),
	.C2V_1 (C2V_145_29),
	.C2V_2 (C2V_145_65),
	.C2V_3 (C2V_145_133),
	.C2V_4 (C2V_145_146),
	.C2V_5 (C2V_145_208),
	.C2V_6 (C2V_145_251),
	.C2V_7 (C2V_145_351),
	.C2V_8 (C2V_145_405),
	.C2V_9 (C2V_145_502),
	.C2V_10 (C2V_145_738),
	.C2V_11 (C2V_145_786),
	.C2V_12 (C2V_145_834),
	.C2V_13 (C2V_145_875),
	.C2V_14 (C2V_145_916),
	.C2V_15 (C2V_145_998),
	.C2V_16 (C2V_145_1037),
	.C2V_17 (C2V_145_1063),
	.C2V_18 (C2V_145_1122),
	.C2V_19 (C2V_145_1296),
	.C2V_20 (C2V_145_1297),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU146 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_38_146),
	.V2C_2 (V2C_87_146),
	.V2C_3 (V2C_143_146),
	.V2C_4 (V2C_191_146),
	.V2C_5 (V2C_220_146),
	.V2C_6 (V2C_241_146),
	.V2C_7 (V2C_292_146),
	.V2C_8 (V2C_399_146),
	.V2C_9 (V2C_488_146),
	.V2C_10 (V2C_648_146),
	.V2C_11 (V2C_709_146),
	.V2C_12 (V2C_829_146),
	.V2C_13 (V2C_871_146),
	.V2C_14 (V2C_934_146),
	.V2C_15 (V2C_965_146),
	.V2C_16 (V2C_1045_146),
	.V2C_17 (V2C_1064_146),
	.V2C_18 (V2C_1143_146),
	.V2C_19 (V2C_1297_146),
	.V2C_20 (V2C_1298_146),
	.C2V_1 (C2V_146_38),
	.C2V_2 (C2V_146_87),
	.C2V_3 (C2V_146_143),
	.C2V_4 (C2V_146_191),
	.C2V_5 (C2V_146_220),
	.C2V_6 (C2V_146_241),
	.C2V_7 (C2V_146_292),
	.C2V_8 (C2V_146_399),
	.C2V_9 (C2V_146_488),
	.C2V_10 (C2V_146_648),
	.C2V_11 (C2V_146_709),
	.C2V_12 (C2V_146_829),
	.C2V_13 (C2V_146_871),
	.C2V_14 (C2V_146_934),
	.C2V_15 (C2V_146_965),
	.C2V_16 (C2V_146_1045),
	.C2V_17 (C2V_146_1064),
	.C2V_18 (C2V_146_1143),
	.C2V_19 (C2V_146_1297),
	.C2V_20 (C2V_146_1298),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU147 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_33_147),
	.V2C_2 (V2C_60_147),
	.V2C_3 (V2C_125_147),
	.V2C_4 (V2C_159_147),
	.V2C_5 (V2C_225_147),
	.V2C_6 (V2C_244_147),
	.V2C_7 (V2C_341_147),
	.V2C_8 (V2C_396_147),
	.V2C_9 (V2C_555_147),
	.V2C_10 (V2C_612_147),
	.V2C_11 (V2C_640_147),
	.V2C_12 (V2C_744_147),
	.V2C_13 (V2C_875_147),
	.V2C_14 (V2C_919_147),
	.V2C_15 (V2C_992_147),
	.V2C_16 (V2C_1052_147),
	.V2C_17 (V2C_1082_147),
	.V2C_18 (V2C_1127_147),
	.V2C_19 (V2C_1298_147),
	.V2C_20 (V2C_1299_147),
	.C2V_1 (C2V_147_33),
	.C2V_2 (C2V_147_60),
	.C2V_3 (C2V_147_125),
	.C2V_4 (C2V_147_159),
	.C2V_5 (C2V_147_225),
	.C2V_6 (C2V_147_244),
	.C2V_7 (C2V_147_341),
	.C2V_8 (C2V_147_396),
	.C2V_9 (C2V_147_555),
	.C2V_10 (C2V_147_612),
	.C2V_11 (C2V_147_640),
	.C2V_12 (C2V_147_744),
	.C2V_13 (C2V_147_875),
	.C2V_14 (C2V_147_919),
	.C2V_15 (C2V_147_992),
	.C2V_16 (C2V_147_1052),
	.C2V_17 (C2V_147_1082),
	.C2V_18 (C2V_147_1127),
	.C2V_19 (C2V_147_1298),
	.C2V_20 (C2V_147_1299),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU148 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_4_148),
	.V2C_2 (V2C_63_148),
	.V2C_3 (V2C_102_148),
	.V2C_4 (V2C_158_148),
	.V2C_5 (V2C_223_148),
	.V2C_6 (V2C_277_148),
	.V2C_7 (V2C_453_148),
	.V2C_8 (V2C_493_148),
	.V2C_9 (V2C_529_148),
	.V2C_10 (V2C_591_148),
	.V2C_11 (V2C_664_148),
	.V2C_12 (V2C_710_148),
	.V2C_13 (V2C_879_148),
	.V2C_14 (V2C_951_148),
	.V2C_15 (V2C_987_148),
	.V2C_16 (V2C_1017_148),
	.V2C_17 (V2C_1092_148),
	.V2C_18 (V2C_1108_148),
	.V2C_19 (V2C_1299_148),
	.V2C_20 (V2C_1300_148),
	.C2V_1 (C2V_148_4),
	.C2V_2 (C2V_148_63),
	.C2V_3 (C2V_148_102),
	.C2V_4 (C2V_148_158),
	.C2V_5 (C2V_148_223),
	.C2V_6 (C2V_148_277),
	.C2V_7 (C2V_148_453),
	.C2V_8 (C2V_148_493),
	.C2V_9 (C2V_148_529),
	.C2V_10 (C2V_148_591),
	.C2V_11 (C2V_148_664),
	.C2V_12 (C2V_148_710),
	.C2V_13 (C2V_148_879),
	.C2V_14 (C2V_148_951),
	.C2V_15 (C2V_148_987),
	.C2V_16 (C2V_148_1017),
	.C2V_17 (C2V_148_1092),
	.C2V_18 (C2V_148_1108),
	.C2V_19 (C2V_148_1299),
	.C2V_20 (C2V_148_1300),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU149 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_23_149),
	.V2C_2 (V2C_81_149),
	.V2C_3 (V2C_116_149),
	.V2C_4 (V2C_187_149),
	.V2C_5 (V2C_203_149),
	.V2C_6 (V2C_269_149),
	.V2C_7 (V2C_318_149),
	.V2C_8 (V2C_337_149),
	.V2C_9 (V2C_464_149),
	.V2C_10 (V2C_698_149),
	.V2C_11 (V2C_762_149),
	.V2C_12 (V2C_816_149),
	.V2C_13 (V2C_894_149),
	.V2C_14 (V2C_942_149),
	.V2C_15 (V2C_985_149),
	.V2C_16 (V2C_1037_149),
	.V2C_17 (V2C_1086_149),
	.V2C_18 (V2C_1134_149),
	.V2C_19 (V2C_1300_149),
	.V2C_20 (V2C_1301_149),
	.C2V_1 (C2V_149_23),
	.C2V_2 (C2V_149_81),
	.C2V_3 (C2V_149_116),
	.C2V_4 (C2V_149_187),
	.C2V_5 (C2V_149_203),
	.C2V_6 (C2V_149_269),
	.C2V_7 (C2V_149_318),
	.C2V_8 (C2V_149_337),
	.C2V_9 (C2V_149_464),
	.C2V_10 (C2V_149_698),
	.C2V_11 (C2V_149_762),
	.C2V_12 (C2V_149_816),
	.C2V_13 (C2V_149_894),
	.C2V_14 (C2V_149_942),
	.C2V_15 (C2V_149_985),
	.C2V_16 (C2V_149_1037),
	.C2V_17 (C2V_149_1086),
	.C2V_18 (C2V_149_1134),
	.C2V_19 (C2V_149_1300),
	.C2V_20 (C2V_149_1301),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU150 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_6_150),
	.V2C_2 (V2C_78_150),
	.V2C_3 (V2C_118_150),
	.V2C_4 (V2C_186_150),
	.V2C_5 (V2C_220_150),
	.V2C_6 (V2C_251_150),
	.V2C_7 (V2C_304_150),
	.V2C_8 (V2C_456_150),
	.V2C_9 (V2C_553_150),
	.V2C_10 (V2C_586_150),
	.V2C_11 (V2C_790_150),
	.V2C_12 (V2C_818_150),
	.V2C_13 (V2C_899_150),
	.V2C_14 (V2C_913_150),
	.V2C_15 (V2C_996_150),
	.V2C_16 (V2C_1015_150),
	.V2C_17 (V2C_1079_150),
	.V2C_18 (V2C_1129_150),
	.V2C_19 (V2C_1301_150),
	.V2C_20 (V2C_1302_150),
	.C2V_1 (C2V_150_6),
	.C2V_2 (C2V_150_78),
	.C2V_3 (C2V_150_118),
	.C2V_4 (C2V_150_186),
	.C2V_5 (C2V_150_220),
	.C2V_6 (C2V_150_251),
	.C2V_7 (C2V_150_304),
	.C2V_8 (C2V_150_456),
	.C2V_9 (C2V_150_553),
	.C2V_10 (C2V_150_586),
	.C2V_11 (C2V_150_790),
	.C2V_12 (C2V_150_818),
	.C2V_13 (C2V_150_899),
	.C2V_14 (C2V_150_913),
	.C2V_15 (C2V_150_996),
	.C2V_16 (C2V_150_1015),
	.C2V_17 (C2V_150_1079),
	.C2V_18 (C2V_150_1129),
	.C2V_19 (C2V_150_1301),
	.C2V_20 (C2V_150_1302),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU151 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_30_151),
	.V2C_2 (V2C_66_151),
	.V2C_3 (V2C_134_151),
	.V2C_4 (V2C_147_151),
	.V2C_5 (V2C_209_151),
	.V2C_6 (V2C_252_151),
	.V2C_7 (V2C_352_151),
	.V2C_8 (V2C_406_151),
	.V2C_9 (V2C_503_151),
	.V2C_10 (V2C_739_151),
	.V2C_11 (V2C_787_151),
	.V2C_12 (V2C_835_151),
	.V2C_13 (V2C_876_151),
	.V2C_14 (V2C_917_151),
	.V2C_15 (V2C_999_151),
	.V2C_16 (V2C_1038_151),
	.V2C_17 (V2C_1064_151),
	.V2C_18 (V2C_1123_151),
	.V2C_19 (V2C_1302_151),
	.V2C_20 (V2C_1303_151),
	.C2V_1 (C2V_151_30),
	.C2V_2 (C2V_151_66),
	.C2V_3 (C2V_151_134),
	.C2V_4 (C2V_151_147),
	.C2V_5 (C2V_151_209),
	.C2V_6 (C2V_151_252),
	.C2V_7 (C2V_151_352),
	.C2V_8 (C2V_151_406),
	.C2V_9 (C2V_151_503),
	.C2V_10 (C2V_151_739),
	.C2V_11 (C2V_151_787),
	.C2V_12 (C2V_151_835),
	.C2V_13 (C2V_151_876),
	.C2V_14 (C2V_151_917),
	.C2V_15 (C2V_151_999),
	.C2V_16 (C2V_151_1038),
	.C2V_17 (C2V_151_1064),
	.C2V_18 (C2V_151_1123),
	.C2V_19 (C2V_151_1302),
	.C2V_20 (C2V_151_1303),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU152 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_39_152),
	.V2C_2 (V2C_88_152),
	.V2C_3 (V2C_144_152),
	.V2C_4 (V2C_192_152),
	.V2C_5 (V2C_221_152),
	.V2C_6 (V2C_242_152),
	.V2C_7 (V2C_293_152),
	.V2C_8 (V2C_400_152),
	.V2C_9 (V2C_489_152),
	.V2C_10 (V2C_649_152),
	.V2C_11 (V2C_710_152),
	.V2C_12 (V2C_830_152),
	.V2C_13 (V2C_872_152),
	.V2C_14 (V2C_935_152),
	.V2C_15 (V2C_966_152),
	.V2C_16 (V2C_1046_152),
	.V2C_17 (V2C_1065_152),
	.V2C_18 (V2C_1144_152),
	.V2C_19 (V2C_1303_152),
	.V2C_20 (V2C_1304_152),
	.C2V_1 (C2V_152_39),
	.C2V_2 (C2V_152_88),
	.C2V_3 (C2V_152_144),
	.C2V_4 (C2V_152_192),
	.C2V_5 (C2V_152_221),
	.C2V_6 (C2V_152_242),
	.C2V_7 (C2V_152_293),
	.C2V_8 (C2V_152_400),
	.C2V_9 (C2V_152_489),
	.C2V_10 (C2V_152_649),
	.C2V_11 (C2V_152_710),
	.C2V_12 (C2V_152_830),
	.C2V_13 (C2V_152_872),
	.C2V_14 (C2V_152_935),
	.C2V_15 (C2V_152_966),
	.C2V_16 (C2V_152_1046),
	.C2V_17 (C2V_152_1065),
	.C2V_18 (C2V_152_1144),
	.C2V_19 (C2V_152_1303),
	.C2V_20 (C2V_152_1304),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU153 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_34_153),
	.V2C_2 (V2C_61_153),
	.V2C_3 (V2C_126_153),
	.V2C_4 (V2C_160_153),
	.V2C_5 (V2C_226_153),
	.V2C_6 (V2C_245_153),
	.V2C_7 (V2C_342_153),
	.V2C_8 (V2C_397_153),
	.V2C_9 (V2C_556_153),
	.V2C_10 (V2C_613_153),
	.V2C_11 (V2C_641_153),
	.V2C_12 (V2C_745_153),
	.V2C_13 (V2C_876_153),
	.V2C_14 (V2C_920_153),
	.V2C_15 (V2C_993_153),
	.V2C_16 (V2C_1053_153),
	.V2C_17 (V2C_1083_153),
	.V2C_18 (V2C_1128_153),
	.V2C_19 (V2C_1304_153),
	.V2C_20 (V2C_1305_153),
	.C2V_1 (C2V_153_34),
	.C2V_2 (C2V_153_61),
	.C2V_3 (C2V_153_126),
	.C2V_4 (C2V_153_160),
	.C2V_5 (C2V_153_226),
	.C2V_6 (C2V_153_245),
	.C2V_7 (C2V_153_342),
	.C2V_8 (C2V_153_397),
	.C2V_9 (C2V_153_556),
	.C2V_10 (C2V_153_613),
	.C2V_11 (C2V_153_641),
	.C2V_12 (C2V_153_745),
	.C2V_13 (C2V_153_876),
	.C2V_14 (C2V_153_920),
	.C2V_15 (C2V_153_993),
	.C2V_16 (C2V_153_1053),
	.C2V_17 (C2V_153_1083),
	.C2V_18 (C2V_153_1128),
	.C2V_19 (C2V_153_1304),
	.C2V_20 (C2V_153_1305),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU154 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_5_154),
	.V2C_2 (V2C_64_154),
	.V2C_3 (V2C_103_154),
	.V2C_4 (V2C_159_154),
	.V2C_5 (V2C_224_154),
	.V2C_6 (V2C_278_154),
	.V2C_7 (V2C_454_154),
	.V2C_8 (V2C_494_154),
	.V2C_9 (V2C_530_154),
	.V2C_10 (V2C_592_154),
	.V2C_11 (V2C_665_154),
	.V2C_12 (V2C_711_154),
	.V2C_13 (V2C_880_154),
	.V2C_14 (V2C_952_154),
	.V2C_15 (V2C_988_154),
	.V2C_16 (V2C_1018_154),
	.V2C_17 (V2C_1093_154),
	.V2C_18 (V2C_1109_154),
	.V2C_19 (V2C_1305_154),
	.V2C_20 (V2C_1306_154),
	.C2V_1 (C2V_154_5),
	.C2V_2 (C2V_154_64),
	.C2V_3 (C2V_154_103),
	.C2V_4 (C2V_154_159),
	.C2V_5 (C2V_154_224),
	.C2V_6 (C2V_154_278),
	.C2V_7 (C2V_154_454),
	.C2V_8 (C2V_154_494),
	.C2V_9 (C2V_154_530),
	.C2V_10 (C2V_154_592),
	.C2V_11 (C2V_154_665),
	.C2V_12 (C2V_154_711),
	.C2V_13 (C2V_154_880),
	.C2V_14 (C2V_154_952),
	.C2V_15 (C2V_154_988),
	.C2V_16 (C2V_154_1018),
	.C2V_17 (C2V_154_1093),
	.C2V_18 (C2V_154_1109),
	.C2V_19 (C2V_154_1305),
	.C2V_20 (C2V_154_1306),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU155 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_24_155),
	.V2C_2 (V2C_82_155),
	.V2C_3 (V2C_117_155),
	.V2C_4 (V2C_188_155),
	.V2C_5 (V2C_204_155),
	.V2C_6 (V2C_270_155),
	.V2C_7 (V2C_319_155),
	.V2C_8 (V2C_338_155),
	.V2C_9 (V2C_465_155),
	.V2C_10 (V2C_699_155),
	.V2C_11 (V2C_763_155),
	.V2C_12 (V2C_769_155),
	.V2C_13 (V2C_895_155),
	.V2C_14 (V2C_943_155),
	.V2C_15 (V2C_986_155),
	.V2C_16 (V2C_1038_155),
	.V2C_17 (V2C_1087_155),
	.V2C_18 (V2C_1135_155),
	.V2C_19 (V2C_1306_155),
	.V2C_20 (V2C_1307_155),
	.C2V_1 (C2V_155_24),
	.C2V_2 (C2V_155_82),
	.C2V_3 (C2V_155_117),
	.C2V_4 (C2V_155_188),
	.C2V_5 (C2V_155_204),
	.C2V_6 (C2V_155_270),
	.C2V_7 (C2V_155_319),
	.C2V_8 (C2V_155_338),
	.C2V_9 (C2V_155_465),
	.C2V_10 (C2V_155_699),
	.C2V_11 (C2V_155_763),
	.C2V_12 (C2V_155_769),
	.C2V_13 (C2V_155_895),
	.C2V_14 (C2V_155_943),
	.C2V_15 (C2V_155_986),
	.C2V_16 (C2V_155_1038),
	.C2V_17 (C2V_155_1087),
	.C2V_18 (C2V_155_1135),
	.C2V_19 (C2V_155_1306),
	.C2V_20 (C2V_155_1307),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU156 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_7_156),
	.V2C_2 (V2C_79_156),
	.V2C_3 (V2C_119_156),
	.V2C_4 (V2C_187_156),
	.V2C_5 (V2C_221_156),
	.V2C_6 (V2C_252_156),
	.V2C_7 (V2C_305_156),
	.V2C_8 (V2C_457_156),
	.V2C_9 (V2C_554_156),
	.V2C_10 (V2C_587_156),
	.V2C_11 (V2C_791_156),
	.V2C_12 (V2C_819_156),
	.V2C_13 (V2C_900_156),
	.V2C_14 (V2C_914_156),
	.V2C_15 (V2C_997_156),
	.V2C_16 (V2C_1016_156),
	.V2C_17 (V2C_1080_156),
	.V2C_18 (V2C_1130_156),
	.V2C_19 (V2C_1307_156),
	.V2C_20 (V2C_1308_156),
	.C2V_1 (C2V_156_7),
	.C2V_2 (C2V_156_79),
	.C2V_3 (C2V_156_119),
	.C2V_4 (C2V_156_187),
	.C2V_5 (C2V_156_221),
	.C2V_6 (C2V_156_252),
	.C2V_7 (C2V_156_305),
	.C2V_8 (C2V_156_457),
	.C2V_9 (C2V_156_554),
	.C2V_10 (C2V_156_587),
	.C2V_11 (C2V_156_791),
	.C2V_12 (C2V_156_819),
	.C2V_13 (C2V_156_900),
	.C2V_14 (C2V_156_914),
	.C2V_15 (C2V_156_997),
	.C2V_16 (C2V_156_1016),
	.C2V_17 (C2V_156_1080),
	.C2V_18 (C2V_156_1130),
	.C2V_19 (C2V_156_1307),
	.C2V_20 (C2V_156_1308),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU157 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_31_157),
	.V2C_2 (V2C_67_157),
	.V2C_3 (V2C_135_157),
	.V2C_4 (V2C_148_157),
	.V2C_5 (V2C_210_157),
	.V2C_6 (V2C_253_157),
	.V2C_7 (V2C_353_157),
	.V2C_8 (V2C_407_157),
	.V2C_9 (V2C_504_157),
	.V2C_10 (V2C_740_157),
	.V2C_11 (V2C_788_157),
	.V2C_12 (V2C_836_157),
	.V2C_13 (V2C_877_157),
	.V2C_14 (V2C_918_157),
	.V2C_15 (V2C_1000_157),
	.V2C_16 (V2C_1039_157),
	.V2C_17 (V2C_1065_157),
	.V2C_18 (V2C_1124_157),
	.V2C_19 (V2C_1308_157),
	.V2C_20 (V2C_1309_157),
	.C2V_1 (C2V_157_31),
	.C2V_2 (C2V_157_67),
	.C2V_3 (C2V_157_135),
	.C2V_4 (C2V_157_148),
	.C2V_5 (C2V_157_210),
	.C2V_6 (C2V_157_253),
	.C2V_7 (C2V_157_353),
	.C2V_8 (C2V_157_407),
	.C2V_9 (C2V_157_504),
	.C2V_10 (C2V_157_740),
	.C2V_11 (C2V_157_788),
	.C2V_12 (C2V_157_836),
	.C2V_13 (C2V_157_877),
	.C2V_14 (C2V_157_918),
	.C2V_15 (C2V_157_1000),
	.C2V_16 (C2V_157_1039),
	.C2V_17 (C2V_157_1065),
	.C2V_18 (C2V_157_1124),
	.C2V_19 (C2V_157_1308),
	.C2V_20 (C2V_157_1309),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU158 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_40_158),
	.V2C_2 (V2C_89_158),
	.V2C_3 (V2C_97_158),
	.V2C_4 (V2C_145_158),
	.V2C_5 (V2C_222_158),
	.V2C_6 (V2C_243_158),
	.V2C_7 (V2C_294_158),
	.V2C_8 (V2C_401_158),
	.V2C_9 (V2C_490_158),
	.V2C_10 (V2C_650_158),
	.V2C_11 (V2C_711_158),
	.V2C_12 (V2C_831_158),
	.V2C_13 (V2C_873_158),
	.V2C_14 (V2C_936_158),
	.V2C_15 (V2C_967_158),
	.V2C_16 (V2C_1047_158),
	.V2C_17 (V2C_1066_158),
	.V2C_18 (V2C_1145_158),
	.V2C_19 (V2C_1309_158),
	.V2C_20 (V2C_1310_158),
	.C2V_1 (C2V_158_40),
	.C2V_2 (C2V_158_89),
	.C2V_3 (C2V_158_97),
	.C2V_4 (C2V_158_145),
	.C2V_5 (C2V_158_222),
	.C2V_6 (C2V_158_243),
	.C2V_7 (C2V_158_294),
	.C2V_8 (C2V_158_401),
	.C2V_9 (C2V_158_490),
	.C2V_10 (C2V_158_650),
	.C2V_11 (C2V_158_711),
	.C2V_12 (C2V_158_831),
	.C2V_13 (C2V_158_873),
	.C2V_14 (C2V_158_936),
	.C2V_15 (C2V_158_967),
	.C2V_16 (C2V_158_1047),
	.C2V_17 (C2V_158_1066),
	.C2V_18 (C2V_158_1145),
	.C2V_19 (C2V_158_1309),
	.C2V_20 (C2V_158_1310),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU159 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_35_159),
	.V2C_2 (V2C_62_159),
	.V2C_3 (V2C_127_159),
	.V2C_4 (V2C_161_159),
	.V2C_5 (V2C_227_159),
	.V2C_6 (V2C_246_159),
	.V2C_7 (V2C_343_159),
	.V2C_8 (V2C_398_159),
	.V2C_9 (V2C_557_159),
	.V2C_10 (V2C_614_159),
	.V2C_11 (V2C_642_159),
	.V2C_12 (V2C_746_159),
	.V2C_13 (V2C_877_159),
	.V2C_14 (V2C_921_159),
	.V2C_15 (V2C_994_159),
	.V2C_16 (V2C_1054_159),
	.V2C_17 (V2C_1084_159),
	.V2C_18 (V2C_1129_159),
	.V2C_19 (V2C_1310_159),
	.V2C_20 (V2C_1311_159),
	.C2V_1 (C2V_159_35),
	.C2V_2 (C2V_159_62),
	.C2V_3 (C2V_159_127),
	.C2V_4 (C2V_159_161),
	.C2V_5 (C2V_159_227),
	.C2V_6 (C2V_159_246),
	.C2V_7 (C2V_159_343),
	.C2V_8 (C2V_159_398),
	.C2V_9 (C2V_159_557),
	.C2V_10 (C2V_159_614),
	.C2V_11 (C2V_159_642),
	.C2V_12 (C2V_159_746),
	.C2V_13 (C2V_159_877),
	.C2V_14 (C2V_159_921),
	.C2V_15 (C2V_159_994),
	.C2V_16 (C2V_159_1054),
	.C2V_17 (C2V_159_1084),
	.C2V_18 (C2V_159_1129),
	.C2V_19 (C2V_159_1310),
	.C2V_20 (C2V_159_1311),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU160 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_6_160),
	.V2C_2 (V2C_65_160),
	.V2C_3 (V2C_104_160),
	.V2C_4 (V2C_160_160),
	.V2C_5 (V2C_225_160),
	.V2C_6 (V2C_279_160),
	.V2C_7 (V2C_455_160),
	.V2C_8 (V2C_495_160),
	.V2C_9 (V2C_531_160),
	.V2C_10 (V2C_593_160),
	.V2C_11 (V2C_666_160),
	.V2C_12 (V2C_712_160),
	.V2C_13 (V2C_881_160),
	.V2C_14 (V2C_953_160),
	.V2C_15 (V2C_989_160),
	.V2C_16 (V2C_1019_160),
	.V2C_17 (V2C_1094_160),
	.V2C_18 (V2C_1110_160),
	.V2C_19 (V2C_1311_160),
	.V2C_20 (V2C_1312_160),
	.C2V_1 (C2V_160_6),
	.C2V_2 (C2V_160_65),
	.C2V_3 (C2V_160_104),
	.C2V_4 (C2V_160_160),
	.C2V_5 (C2V_160_225),
	.C2V_6 (C2V_160_279),
	.C2V_7 (C2V_160_455),
	.C2V_8 (C2V_160_495),
	.C2V_9 (C2V_160_531),
	.C2V_10 (C2V_160_593),
	.C2V_11 (C2V_160_666),
	.C2V_12 (C2V_160_712),
	.C2V_13 (C2V_160_881),
	.C2V_14 (C2V_160_953),
	.C2V_15 (C2V_160_989),
	.C2V_16 (C2V_160_1019),
	.C2V_17 (C2V_160_1094),
	.C2V_18 (C2V_160_1110),
	.C2V_19 (C2V_160_1311),
	.C2V_20 (C2V_160_1312),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU161 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_25_161),
	.V2C_2 (V2C_83_161),
	.V2C_3 (V2C_118_161),
	.V2C_4 (V2C_189_161),
	.V2C_5 (V2C_205_161),
	.V2C_6 (V2C_271_161),
	.V2C_7 (V2C_320_161),
	.V2C_8 (V2C_339_161),
	.V2C_9 (V2C_466_161),
	.V2C_10 (V2C_700_161),
	.V2C_11 (V2C_764_161),
	.V2C_12 (V2C_770_161),
	.V2C_13 (V2C_896_161),
	.V2C_14 (V2C_944_161),
	.V2C_15 (V2C_987_161),
	.V2C_16 (V2C_1039_161),
	.V2C_17 (V2C_1088_161),
	.V2C_18 (V2C_1136_161),
	.V2C_19 (V2C_1312_161),
	.V2C_20 (V2C_1313_161),
	.C2V_1 (C2V_161_25),
	.C2V_2 (C2V_161_83),
	.C2V_3 (C2V_161_118),
	.C2V_4 (C2V_161_189),
	.C2V_5 (C2V_161_205),
	.C2V_6 (C2V_161_271),
	.C2V_7 (C2V_161_320),
	.C2V_8 (C2V_161_339),
	.C2V_9 (C2V_161_466),
	.C2V_10 (C2V_161_700),
	.C2V_11 (C2V_161_764),
	.C2V_12 (C2V_161_770),
	.C2V_13 (C2V_161_896),
	.C2V_14 (C2V_161_944),
	.C2V_15 (C2V_161_987),
	.C2V_16 (C2V_161_1039),
	.C2V_17 (C2V_161_1088),
	.C2V_18 (C2V_161_1136),
	.C2V_19 (C2V_161_1312),
	.C2V_20 (C2V_161_1313),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU162 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_8_162),
	.V2C_2 (V2C_80_162),
	.V2C_3 (V2C_120_162),
	.V2C_4 (V2C_188_162),
	.V2C_5 (V2C_222_162),
	.V2C_6 (V2C_253_162),
	.V2C_7 (V2C_306_162),
	.V2C_8 (V2C_458_162),
	.V2C_9 (V2C_555_162),
	.V2C_10 (V2C_588_162),
	.V2C_11 (V2C_792_162),
	.V2C_12 (V2C_820_162),
	.V2C_13 (V2C_901_162),
	.V2C_14 (V2C_915_162),
	.V2C_15 (V2C_998_162),
	.V2C_16 (V2C_1017_162),
	.V2C_17 (V2C_1081_162),
	.V2C_18 (V2C_1131_162),
	.V2C_19 (V2C_1313_162),
	.V2C_20 (V2C_1314_162),
	.C2V_1 (C2V_162_8),
	.C2V_2 (C2V_162_80),
	.C2V_3 (C2V_162_120),
	.C2V_4 (C2V_162_188),
	.C2V_5 (C2V_162_222),
	.C2V_6 (C2V_162_253),
	.C2V_7 (C2V_162_306),
	.C2V_8 (C2V_162_458),
	.C2V_9 (C2V_162_555),
	.C2V_10 (C2V_162_588),
	.C2V_11 (C2V_162_792),
	.C2V_12 (C2V_162_820),
	.C2V_13 (C2V_162_901),
	.C2V_14 (C2V_162_915),
	.C2V_15 (C2V_162_998),
	.C2V_16 (C2V_162_1017),
	.C2V_17 (C2V_162_1081),
	.C2V_18 (C2V_162_1131),
	.C2V_19 (C2V_162_1313),
	.C2V_20 (C2V_162_1314),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU163 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_32_163),
	.V2C_2 (V2C_68_163),
	.V2C_3 (V2C_136_163),
	.V2C_4 (V2C_149_163),
	.V2C_5 (V2C_211_163),
	.V2C_6 (V2C_254_163),
	.V2C_7 (V2C_354_163),
	.V2C_8 (V2C_408_163),
	.V2C_9 (V2C_505_163),
	.V2C_10 (V2C_741_163),
	.V2C_11 (V2C_789_163),
	.V2C_12 (V2C_837_163),
	.V2C_13 (V2C_878_163),
	.V2C_14 (V2C_919_163),
	.V2C_15 (V2C_1001_163),
	.V2C_16 (V2C_1040_163),
	.V2C_17 (V2C_1066_163),
	.V2C_18 (V2C_1125_163),
	.V2C_19 (V2C_1314_163),
	.V2C_20 (V2C_1315_163),
	.C2V_1 (C2V_163_32),
	.C2V_2 (C2V_163_68),
	.C2V_3 (C2V_163_136),
	.C2V_4 (C2V_163_149),
	.C2V_5 (C2V_163_211),
	.C2V_6 (C2V_163_254),
	.C2V_7 (C2V_163_354),
	.C2V_8 (C2V_163_408),
	.C2V_9 (C2V_163_505),
	.C2V_10 (C2V_163_741),
	.C2V_11 (C2V_163_789),
	.C2V_12 (C2V_163_837),
	.C2V_13 (C2V_163_878),
	.C2V_14 (C2V_163_919),
	.C2V_15 (C2V_163_1001),
	.C2V_16 (C2V_163_1040),
	.C2V_17 (C2V_163_1066),
	.C2V_18 (C2V_163_1125),
	.C2V_19 (C2V_163_1314),
	.C2V_20 (C2V_163_1315),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU164 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_41_164),
	.V2C_2 (V2C_90_164),
	.V2C_3 (V2C_98_164),
	.V2C_4 (V2C_146_164),
	.V2C_5 (V2C_223_164),
	.V2C_6 (V2C_244_164),
	.V2C_7 (V2C_295_164),
	.V2C_8 (V2C_402_164),
	.V2C_9 (V2C_491_164),
	.V2C_10 (V2C_651_164),
	.V2C_11 (V2C_712_164),
	.V2C_12 (V2C_832_164),
	.V2C_13 (V2C_874_164),
	.V2C_14 (V2C_937_164),
	.V2C_15 (V2C_968_164),
	.V2C_16 (V2C_1048_164),
	.V2C_17 (V2C_1067_164),
	.V2C_18 (V2C_1146_164),
	.V2C_19 (V2C_1315_164),
	.V2C_20 (V2C_1316_164),
	.C2V_1 (C2V_164_41),
	.C2V_2 (C2V_164_90),
	.C2V_3 (C2V_164_98),
	.C2V_4 (C2V_164_146),
	.C2V_5 (C2V_164_223),
	.C2V_6 (C2V_164_244),
	.C2V_7 (C2V_164_295),
	.C2V_8 (C2V_164_402),
	.C2V_9 (C2V_164_491),
	.C2V_10 (C2V_164_651),
	.C2V_11 (C2V_164_712),
	.C2V_12 (C2V_164_832),
	.C2V_13 (C2V_164_874),
	.C2V_14 (C2V_164_937),
	.C2V_15 (C2V_164_968),
	.C2V_16 (C2V_164_1048),
	.C2V_17 (C2V_164_1067),
	.C2V_18 (C2V_164_1146),
	.C2V_19 (C2V_164_1315),
	.C2V_20 (C2V_164_1316),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU165 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_36_165),
	.V2C_2 (V2C_63_165),
	.V2C_3 (V2C_128_165),
	.V2C_4 (V2C_162_165),
	.V2C_5 (V2C_228_165),
	.V2C_6 (V2C_247_165),
	.V2C_7 (V2C_344_165),
	.V2C_8 (V2C_399_165),
	.V2C_9 (V2C_558_165),
	.V2C_10 (V2C_615_165),
	.V2C_11 (V2C_643_165),
	.V2C_12 (V2C_747_165),
	.V2C_13 (V2C_878_165),
	.V2C_14 (V2C_922_165),
	.V2C_15 (V2C_995_165),
	.V2C_16 (V2C_1055_165),
	.V2C_17 (V2C_1085_165),
	.V2C_18 (V2C_1130_165),
	.V2C_19 (V2C_1316_165),
	.V2C_20 (V2C_1317_165),
	.C2V_1 (C2V_165_36),
	.C2V_2 (C2V_165_63),
	.C2V_3 (C2V_165_128),
	.C2V_4 (C2V_165_162),
	.C2V_5 (C2V_165_228),
	.C2V_6 (C2V_165_247),
	.C2V_7 (C2V_165_344),
	.C2V_8 (C2V_165_399),
	.C2V_9 (C2V_165_558),
	.C2V_10 (C2V_165_615),
	.C2V_11 (C2V_165_643),
	.C2V_12 (C2V_165_747),
	.C2V_13 (C2V_165_878),
	.C2V_14 (C2V_165_922),
	.C2V_15 (C2V_165_995),
	.C2V_16 (C2V_165_1055),
	.C2V_17 (C2V_165_1085),
	.C2V_18 (C2V_165_1130),
	.C2V_19 (C2V_165_1316),
	.C2V_20 (C2V_165_1317),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU166 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_7_166),
	.V2C_2 (V2C_66_166),
	.V2C_3 (V2C_105_166),
	.V2C_4 (V2C_161_166),
	.V2C_5 (V2C_226_166),
	.V2C_6 (V2C_280_166),
	.V2C_7 (V2C_456_166),
	.V2C_8 (V2C_496_166),
	.V2C_9 (V2C_532_166),
	.V2C_10 (V2C_594_166),
	.V2C_11 (V2C_667_166),
	.V2C_12 (V2C_713_166),
	.V2C_13 (V2C_882_166),
	.V2C_14 (V2C_954_166),
	.V2C_15 (V2C_990_166),
	.V2C_16 (V2C_1020_166),
	.V2C_17 (V2C_1095_166),
	.V2C_18 (V2C_1111_166),
	.V2C_19 (V2C_1317_166),
	.V2C_20 (V2C_1318_166),
	.C2V_1 (C2V_166_7),
	.C2V_2 (C2V_166_66),
	.C2V_3 (C2V_166_105),
	.C2V_4 (C2V_166_161),
	.C2V_5 (C2V_166_226),
	.C2V_6 (C2V_166_280),
	.C2V_7 (C2V_166_456),
	.C2V_8 (C2V_166_496),
	.C2V_9 (C2V_166_532),
	.C2V_10 (C2V_166_594),
	.C2V_11 (C2V_166_667),
	.C2V_12 (C2V_166_713),
	.C2V_13 (C2V_166_882),
	.C2V_14 (C2V_166_954),
	.C2V_15 (C2V_166_990),
	.C2V_16 (C2V_166_1020),
	.C2V_17 (C2V_166_1095),
	.C2V_18 (C2V_166_1111),
	.C2V_19 (C2V_166_1317),
	.C2V_20 (C2V_166_1318),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU167 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_26_167),
	.V2C_2 (V2C_84_167),
	.V2C_3 (V2C_119_167),
	.V2C_4 (V2C_190_167),
	.V2C_5 (V2C_206_167),
	.V2C_6 (V2C_272_167),
	.V2C_7 (V2C_321_167),
	.V2C_8 (V2C_340_167),
	.V2C_9 (V2C_467_167),
	.V2C_10 (V2C_701_167),
	.V2C_11 (V2C_765_167),
	.V2C_12 (V2C_771_167),
	.V2C_13 (V2C_897_167),
	.V2C_14 (V2C_945_167),
	.V2C_15 (V2C_988_167),
	.V2C_16 (V2C_1040_167),
	.V2C_17 (V2C_1089_167),
	.V2C_18 (V2C_1137_167),
	.V2C_19 (V2C_1318_167),
	.V2C_20 (V2C_1319_167),
	.C2V_1 (C2V_167_26),
	.C2V_2 (C2V_167_84),
	.C2V_3 (C2V_167_119),
	.C2V_4 (C2V_167_190),
	.C2V_5 (C2V_167_206),
	.C2V_6 (C2V_167_272),
	.C2V_7 (C2V_167_321),
	.C2V_8 (C2V_167_340),
	.C2V_9 (C2V_167_467),
	.C2V_10 (C2V_167_701),
	.C2V_11 (C2V_167_765),
	.C2V_12 (C2V_167_771),
	.C2V_13 (C2V_167_897),
	.C2V_14 (C2V_167_945),
	.C2V_15 (C2V_167_988),
	.C2V_16 (C2V_167_1040),
	.C2V_17 (C2V_167_1089),
	.C2V_18 (C2V_167_1137),
	.C2V_19 (C2V_167_1318),
	.C2V_20 (C2V_167_1319),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU168 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_9_168),
	.V2C_2 (V2C_81_168),
	.V2C_3 (V2C_121_168),
	.V2C_4 (V2C_189_168),
	.V2C_5 (V2C_223_168),
	.V2C_6 (V2C_254_168),
	.V2C_7 (V2C_307_168),
	.V2C_8 (V2C_459_168),
	.V2C_9 (V2C_556_168),
	.V2C_10 (V2C_589_168),
	.V2C_11 (V2C_793_168),
	.V2C_12 (V2C_821_168),
	.V2C_13 (V2C_902_168),
	.V2C_14 (V2C_916_168),
	.V2C_15 (V2C_999_168),
	.V2C_16 (V2C_1018_168),
	.V2C_17 (V2C_1082_168),
	.V2C_18 (V2C_1132_168),
	.V2C_19 (V2C_1319_168),
	.V2C_20 (V2C_1320_168),
	.C2V_1 (C2V_168_9),
	.C2V_2 (C2V_168_81),
	.C2V_3 (C2V_168_121),
	.C2V_4 (C2V_168_189),
	.C2V_5 (C2V_168_223),
	.C2V_6 (C2V_168_254),
	.C2V_7 (C2V_168_307),
	.C2V_8 (C2V_168_459),
	.C2V_9 (C2V_168_556),
	.C2V_10 (C2V_168_589),
	.C2V_11 (C2V_168_793),
	.C2V_12 (C2V_168_821),
	.C2V_13 (C2V_168_902),
	.C2V_14 (C2V_168_916),
	.C2V_15 (C2V_168_999),
	.C2V_16 (C2V_168_1018),
	.C2V_17 (C2V_168_1082),
	.C2V_18 (C2V_168_1132),
	.C2V_19 (C2V_168_1319),
	.C2V_20 (C2V_168_1320),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU169 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_33_169),
	.V2C_2 (V2C_69_169),
	.V2C_3 (V2C_137_169),
	.V2C_4 (V2C_150_169),
	.V2C_5 (V2C_212_169),
	.V2C_6 (V2C_255_169),
	.V2C_7 (V2C_355_169),
	.V2C_8 (V2C_409_169),
	.V2C_9 (V2C_506_169),
	.V2C_10 (V2C_742_169),
	.V2C_11 (V2C_790_169),
	.V2C_12 (V2C_838_169),
	.V2C_13 (V2C_879_169),
	.V2C_14 (V2C_920_169),
	.V2C_15 (V2C_1002_169),
	.V2C_16 (V2C_1041_169),
	.V2C_17 (V2C_1067_169),
	.V2C_18 (V2C_1126_169),
	.V2C_19 (V2C_1320_169),
	.V2C_20 (V2C_1321_169),
	.C2V_1 (C2V_169_33),
	.C2V_2 (C2V_169_69),
	.C2V_3 (C2V_169_137),
	.C2V_4 (C2V_169_150),
	.C2V_5 (C2V_169_212),
	.C2V_6 (C2V_169_255),
	.C2V_7 (C2V_169_355),
	.C2V_8 (C2V_169_409),
	.C2V_9 (C2V_169_506),
	.C2V_10 (C2V_169_742),
	.C2V_11 (C2V_169_790),
	.C2V_12 (C2V_169_838),
	.C2V_13 (C2V_169_879),
	.C2V_14 (C2V_169_920),
	.C2V_15 (C2V_169_1002),
	.C2V_16 (C2V_169_1041),
	.C2V_17 (C2V_169_1067),
	.C2V_18 (C2V_169_1126),
	.C2V_19 (C2V_169_1320),
	.C2V_20 (C2V_169_1321),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU170 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_42_170),
	.V2C_2 (V2C_91_170),
	.V2C_3 (V2C_99_170),
	.V2C_4 (V2C_147_170),
	.V2C_5 (V2C_224_170),
	.V2C_6 (V2C_245_170),
	.V2C_7 (V2C_296_170),
	.V2C_8 (V2C_403_170),
	.V2C_9 (V2C_492_170),
	.V2C_10 (V2C_652_170),
	.V2C_11 (V2C_713_170),
	.V2C_12 (V2C_833_170),
	.V2C_13 (V2C_875_170),
	.V2C_14 (V2C_938_170),
	.V2C_15 (V2C_969_170),
	.V2C_16 (V2C_1049_170),
	.V2C_17 (V2C_1068_170),
	.V2C_18 (V2C_1147_170),
	.V2C_19 (V2C_1321_170),
	.V2C_20 (V2C_1322_170),
	.C2V_1 (C2V_170_42),
	.C2V_2 (C2V_170_91),
	.C2V_3 (C2V_170_99),
	.C2V_4 (C2V_170_147),
	.C2V_5 (C2V_170_224),
	.C2V_6 (C2V_170_245),
	.C2V_7 (C2V_170_296),
	.C2V_8 (C2V_170_403),
	.C2V_9 (C2V_170_492),
	.C2V_10 (C2V_170_652),
	.C2V_11 (C2V_170_713),
	.C2V_12 (C2V_170_833),
	.C2V_13 (C2V_170_875),
	.C2V_14 (C2V_170_938),
	.C2V_15 (C2V_170_969),
	.C2V_16 (C2V_170_1049),
	.C2V_17 (C2V_170_1068),
	.C2V_18 (C2V_170_1147),
	.C2V_19 (C2V_170_1321),
	.C2V_20 (C2V_170_1322),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU171 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_37_171),
	.V2C_2 (V2C_64_171),
	.V2C_3 (V2C_129_171),
	.V2C_4 (V2C_163_171),
	.V2C_5 (V2C_229_171),
	.V2C_6 (V2C_248_171),
	.V2C_7 (V2C_345_171),
	.V2C_8 (V2C_400_171),
	.V2C_9 (V2C_559_171),
	.V2C_10 (V2C_616_171),
	.V2C_11 (V2C_644_171),
	.V2C_12 (V2C_748_171),
	.V2C_13 (V2C_879_171),
	.V2C_14 (V2C_923_171),
	.V2C_15 (V2C_996_171),
	.V2C_16 (V2C_1056_171),
	.V2C_17 (V2C_1086_171),
	.V2C_18 (V2C_1131_171),
	.V2C_19 (V2C_1322_171),
	.V2C_20 (V2C_1323_171),
	.C2V_1 (C2V_171_37),
	.C2V_2 (C2V_171_64),
	.C2V_3 (C2V_171_129),
	.C2V_4 (C2V_171_163),
	.C2V_5 (C2V_171_229),
	.C2V_6 (C2V_171_248),
	.C2V_7 (C2V_171_345),
	.C2V_8 (C2V_171_400),
	.C2V_9 (C2V_171_559),
	.C2V_10 (C2V_171_616),
	.C2V_11 (C2V_171_644),
	.C2V_12 (C2V_171_748),
	.C2V_13 (C2V_171_879),
	.C2V_14 (C2V_171_923),
	.C2V_15 (C2V_171_996),
	.C2V_16 (C2V_171_1056),
	.C2V_17 (C2V_171_1086),
	.C2V_18 (C2V_171_1131),
	.C2V_19 (C2V_171_1322),
	.C2V_20 (C2V_171_1323),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU172 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_8_172),
	.V2C_2 (V2C_67_172),
	.V2C_3 (V2C_106_172),
	.V2C_4 (V2C_162_172),
	.V2C_5 (V2C_227_172),
	.V2C_6 (V2C_281_172),
	.V2C_7 (V2C_457_172),
	.V2C_8 (V2C_497_172),
	.V2C_9 (V2C_533_172),
	.V2C_10 (V2C_595_172),
	.V2C_11 (V2C_668_172),
	.V2C_12 (V2C_714_172),
	.V2C_13 (V2C_883_172),
	.V2C_14 (V2C_955_172),
	.V2C_15 (V2C_991_172),
	.V2C_16 (V2C_1021_172),
	.V2C_17 (V2C_1096_172),
	.V2C_18 (V2C_1112_172),
	.V2C_19 (V2C_1323_172),
	.V2C_20 (V2C_1324_172),
	.C2V_1 (C2V_172_8),
	.C2V_2 (C2V_172_67),
	.C2V_3 (C2V_172_106),
	.C2V_4 (C2V_172_162),
	.C2V_5 (C2V_172_227),
	.C2V_6 (C2V_172_281),
	.C2V_7 (C2V_172_457),
	.C2V_8 (C2V_172_497),
	.C2V_9 (C2V_172_533),
	.C2V_10 (C2V_172_595),
	.C2V_11 (C2V_172_668),
	.C2V_12 (C2V_172_714),
	.C2V_13 (C2V_172_883),
	.C2V_14 (C2V_172_955),
	.C2V_15 (C2V_172_991),
	.C2V_16 (C2V_172_1021),
	.C2V_17 (C2V_172_1096),
	.C2V_18 (C2V_172_1112),
	.C2V_19 (C2V_172_1323),
	.C2V_20 (C2V_172_1324),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU173 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_27_173),
	.V2C_2 (V2C_85_173),
	.V2C_3 (V2C_120_173),
	.V2C_4 (V2C_191_173),
	.V2C_5 (V2C_207_173),
	.V2C_6 (V2C_273_173),
	.V2C_7 (V2C_322_173),
	.V2C_8 (V2C_341_173),
	.V2C_9 (V2C_468_173),
	.V2C_10 (V2C_702_173),
	.V2C_11 (V2C_766_173),
	.V2C_12 (V2C_772_173),
	.V2C_13 (V2C_898_173),
	.V2C_14 (V2C_946_173),
	.V2C_15 (V2C_989_173),
	.V2C_16 (V2C_1041_173),
	.V2C_17 (V2C_1090_173),
	.V2C_18 (V2C_1138_173),
	.V2C_19 (V2C_1324_173),
	.V2C_20 (V2C_1325_173),
	.C2V_1 (C2V_173_27),
	.C2V_2 (C2V_173_85),
	.C2V_3 (C2V_173_120),
	.C2V_4 (C2V_173_191),
	.C2V_5 (C2V_173_207),
	.C2V_6 (C2V_173_273),
	.C2V_7 (C2V_173_322),
	.C2V_8 (C2V_173_341),
	.C2V_9 (C2V_173_468),
	.C2V_10 (C2V_173_702),
	.C2V_11 (C2V_173_766),
	.C2V_12 (C2V_173_772),
	.C2V_13 (C2V_173_898),
	.C2V_14 (C2V_173_946),
	.C2V_15 (C2V_173_989),
	.C2V_16 (C2V_173_1041),
	.C2V_17 (C2V_173_1090),
	.C2V_18 (C2V_173_1138),
	.C2V_19 (C2V_173_1324),
	.C2V_20 (C2V_173_1325),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU174 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_10_174),
	.V2C_2 (V2C_82_174),
	.V2C_3 (V2C_122_174),
	.V2C_4 (V2C_190_174),
	.V2C_5 (V2C_224_174),
	.V2C_6 (V2C_255_174),
	.V2C_7 (V2C_308_174),
	.V2C_8 (V2C_460_174),
	.V2C_9 (V2C_557_174),
	.V2C_10 (V2C_590_174),
	.V2C_11 (V2C_794_174),
	.V2C_12 (V2C_822_174),
	.V2C_13 (V2C_903_174),
	.V2C_14 (V2C_917_174),
	.V2C_15 (V2C_1000_174),
	.V2C_16 (V2C_1019_174),
	.V2C_17 (V2C_1083_174),
	.V2C_18 (V2C_1133_174),
	.V2C_19 (V2C_1325_174),
	.V2C_20 (V2C_1326_174),
	.C2V_1 (C2V_174_10),
	.C2V_2 (C2V_174_82),
	.C2V_3 (C2V_174_122),
	.C2V_4 (C2V_174_190),
	.C2V_5 (C2V_174_224),
	.C2V_6 (C2V_174_255),
	.C2V_7 (C2V_174_308),
	.C2V_8 (C2V_174_460),
	.C2V_9 (C2V_174_557),
	.C2V_10 (C2V_174_590),
	.C2V_11 (C2V_174_794),
	.C2V_12 (C2V_174_822),
	.C2V_13 (C2V_174_903),
	.C2V_14 (C2V_174_917),
	.C2V_15 (C2V_174_1000),
	.C2V_16 (C2V_174_1019),
	.C2V_17 (C2V_174_1083),
	.C2V_18 (C2V_174_1133),
	.C2V_19 (C2V_174_1325),
	.C2V_20 (C2V_174_1326),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU175 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_34_175),
	.V2C_2 (V2C_70_175),
	.V2C_3 (V2C_138_175),
	.V2C_4 (V2C_151_175),
	.V2C_5 (V2C_213_175),
	.V2C_6 (V2C_256_175),
	.V2C_7 (V2C_356_175),
	.V2C_8 (V2C_410_175),
	.V2C_9 (V2C_507_175),
	.V2C_10 (V2C_743_175),
	.V2C_11 (V2C_791_175),
	.V2C_12 (V2C_839_175),
	.V2C_13 (V2C_880_175),
	.V2C_14 (V2C_921_175),
	.V2C_15 (V2C_1003_175),
	.V2C_16 (V2C_1042_175),
	.V2C_17 (V2C_1068_175),
	.V2C_18 (V2C_1127_175),
	.V2C_19 (V2C_1326_175),
	.V2C_20 (V2C_1327_175),
	.C2V_1 (C2V_175_34),
	.C2V_2 (C2V_175_70),
	.C2V_3 (C2V_175_138),
	.C2V_4 (C2V_175_151),
	.C2V_5 (C2V_175_213),
	.C2V_6 (C2V_175_256),
	.C2V_7 (C2V_175_356),
	.C2V_8 (C2V_175_410),
	.C2V_9 (C2V_175_507),
	.C2V_10 (C2V_175_743),
	.C2V_11 (C2V_175_791),
	.C2V_12 (C2V_175_839),
	.C2V_13 (C2V_175_880),
	.C2V_14 (C2V_175_921),
	.C2V_15 (C2V_175_1003),
	.C2V_16 (C2V_175_1042),
	.C2V_17 (C2V_175_1068),
	.C2V_18 (C2V_175_1127),
	.C2V_19 (C2V_175_1326),
	.C2V_20 (C2V_175_1327),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU176 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_43_176),
	.V2C_2 (V2C_92_176),
	.V2C_3 (V2C_100_176),
	.V2C_4 (V2C_148_176),
	.V2C_5 (V2C_225_176),
	.V2C_6 (V2C_246_176),
	.V2C_7 (V2C_297_176),
	.V2C_8 (V2C_404_176),
	.V2C_9 (V2C_493_176),
	.V2C_10 (V2C_653_176),
	.V2C_11 (V2C_714_176),
	.V2C_12 (V2C_834_176),
	.V2C_13 (V2C_876_176),
	.V2C_14 (V2C_939_176),
	.V2C_15 (V2C_970_176),
	.V2C_16 (V2C_1050_176),
	.V2C_17 (V2C_1069_176),
	.V2C_18 (V2C_1148_176),
	.V2C_19 (V2C_1327_176),
	.V2C_20 (V2C_1328_176),
	.C2V_1 (C2V_176_43),
	.C2V_2 (C2V_176_92),
	.C2V_3 (C2V_176_100),
	.C2V_4 (C2V_176_148),
	.C2V_5 (C2V_176_225),
	.C2V_6 (C2V_176_246),
	.C2V_7 (C2V_176_297),
	.C2V_8 (C2V_176_404),
	.C2V_9 (C2V_176_493),
	.C2V_10 (C2V_176_653),
	.C2V_11 (C2V_176_714),
	.C2V_12 (C2V_176_834),
	.C2V_13 (C2V_176_876),
	.C2V_14 (C2V_176_939),
	.C2V_15 (C2V_176_970),
	.C2V_16 (C2V_176_1050),
	.C2V_17 (C2V_176_1069),
	.C2V_18 (C2V_176_1148),
	.C2V_19 (C2V_176_1327),
	.C2V_20 (C2V_176_1328),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU177 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_38_177),
	.V2C_2 (V2C_65_177),
	.V2C_3 (V2C_130_177),
	.V2C_4 (V2C_164_177),
	.V2C_5 (V2C_230_177),
	.V2C_6 (V2C_249_177),
	.V2C_7 (V2C_346_177),
	.V2C_8 (V2C_401_177),
	.V2C_9 (V2C_560_177),
	.V2C_10 (V2C_617_177),
	.V2C_11 (V2C_645_177),
	.V2C_12 (V2C_749_177),
	.V2C_13 (V2C_880_177),
	.V2C_14 (V2C_924_177),
	.V2C_15 (V2C_997_177),
	.V2C_16 (V2C_1009_177),
	.V2C_17 (V2C_1087_177),
	.V2C_18 (V2C_1132_177),
	.V2C_19 (V2C_1328_177),
	.V2C_20 (V2C_1329_177),
	.C2V_1 (C2V_177_38),
	.C2V_2 (C2V_177_65),
	.C2V_3 (C2V_177_130),
	.C2V_4 (C2V_177_164),
	.C2V_5 (C2V_177_230),
	.C2V_6 (C2V_177_249),
	.C2V_7 (C2V_177_346),
	.C2V_8 (C2V_177_401),
	.C2V_9 (C2V_177_560),
	.C2V_10 (C2V_177_617),
	.C2V_11 (C2V_177_645),
	.C2V_12 (C2V_177_749),
	.C2V_13 (C2V_177_880),
	.C2V_14 (C2V_177_924),
	.C2V_15 (C2V_177_997),
	.C2V_16 (C2V_177_1009),
	.C2V_17 (C2V_177_1087),
	.C2V_18 (C2V_177_1132),
	.C2V_19 (C2V_177_1328),
	.C2V_20 (C2V_177_1329),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU178 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_9_178),
	.V2C_2 (V2C_68_178),
	.V2C_3 (V2C_107_178),
	.V2C_4 (V2C_163_178),
	.V2C_5 (V2C_228_178),
	.V2C_6 (V2C_282_178),
	.V2C_7 (V2C_458_178),
	.V2C_8 (V2C_498_178),
	.V2C_9 (V2C_534_178),
	.V2C_10 (V2C_596_178),
	.V2C_11 (V2C_669_178),
	.V2C_12 (V2C_715_178),
	.V2C_13 (V2C_884_178),
	.V2C_14 (V2C_956_178),
	.V2C_15 (V2C_992_178),
	.V2C_16 (V2C_1022_178),
	.V2C_17 (V2C_1097_178),
	.V2C_18 (V2C_1113_178),
	.V2C_19 (V2C_1329_178),
	.V2C_20 (V2C_1330_178),
	.C2V_1 (C2V_178_9),
	.C2V_2 (C2V_178_68),
	.C2V_3 (C2V_178_107),
	.C2V_4 (C2V_178_163),
	.C2V_5 (C2V_178_228),
	.C2V_6 (C2V_178_282),
	.C2V_7 (C2V_178_458),
	.C2V_8 (C2V_178_498),
	.C2V_9 (C2V_178_534),
	.C2V_10 (C2V_178_596),
	.C2V_11 (C2V_178_669),
	.C2V_12 (C2V_178_715),
	.C2V_13 (C2V_178_884),
	.C2V_14 (C2V_178_956),
	.C2V_15 (C2V_178_992),
	.C2V_16 (C2V_178_1022),
	.C2V_17 (C2V_178_1097),
	.C2V_18 (C2V_178_1113),
	.C2V_19 (C2V_178_1329),
	.C2V_20 (C2V_178_1330),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU179 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_28_179),
	.V2C_2 (V2C_86_179),
	.V2C_3 (V2C_121_179),
	.V2C_4 (V2C_192_179),
	.V2C_5 (V2C_208_179),
	.V2C_6 (V2C_274_179),
	.V2C_7 (V2C_323_179),
	.V2C_8 (V2C_342_179),
	.V2C_9 (V2C_469_179),
	.V2C_10 (V2C_703_179),
	.V2C_11 (V2C_767_179),
	.V2C_12 (V2C_773_179),
	.V2C_13 (V2C_899_179),
	.V2C_14 (V2C_947_179),
	.V2C_15 (V2C_990_179),
	.V2C_16 (V2C_1042_179),
	.V2C_17 (V2C_1091_179),
	.V2C_18 (V2C_1139_179),
	.V2C_19 (V2C_1330_179),
	.V2C_20 (V2C_1331_179),
	.C2V_1 (C2V_179_28),
	.C2V_2 (C2V_179_86),
	.C2V_3 (C2V_179_121),
	.C2V_4 (C2V_179_192),
	.C2V_5 (C2V_179_208),
	.C2V_6 (C2V_179_274),
	.C2V_7 (C2V_179_323),
	.C2V_8 (C2V_179_342),
	.C2V_9 (C2V_179_469),
	.C2V_10 (C2V_179_703),
	.C2V_11 (C2V_179_767),
	.C2V_12 (C2V_179_773),
	.C2V_13 (C2V_179_899),
	.C2V_14 (C2V_179_947),
	.C2V_15 (C2V_179_990),
	.C2V_16 (C2V_179_1042),
	.C2V_17 (C2V_179_1091),
	.C2V_18 (C2V_179_1139),
	.C2V_19 (C2V_179_1330),
	.C2V_20 (C2V_179_1331),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU180 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_11_180),
	.V2C_2 (V2C_83_180),
	.V2C_3 (V2C_123_180),
	.V2C_4 (V2C_191_180),
	.V2C_5 (V2C_225_180),
	.V2C_6 (V2C_256_180),
	.V2C_7 (V2C_309_180),
	.V2C_8 (V2C_461_180),
	.V2C_9 (V2C_558_180),
	.V2C_10 (V2C_591_180),
	.V2C_11 (V2C_795_180),
	.V2C_12 (V2C_823_180),
	.V2C_13 (V2C_904_180),
	.V2C_14 (V2C_918_180),
	.V2C_15 (V2C_1001_180),
	.V2C_16 (V2C_1020_180),
	.V2C_17 (V2C_1084_180),
	.V2C_18 (V2C_1134_180),
	.V2C_19 (V2C_1331_180),
	.V2C_20 (V2C_1332_180),
	.C2V_1 (C2V_180_11),
	.C2V_2 (C2V_180_83),
	.C2V_3 (C2V_180_123),
	.C2V_4 (C2V_180_191),
	.C2V_5 (C2V_180_225),
	.C2V_6 (C2V_180_256),
	.C2V_7 (C2V_180_309),
	.C2V_8 (C2V_180_461),
	.C2V_9 (C2V_180_558),
	.C2V_10 (C2V_180_591),
	.C2V_11 (C2V_180_795),
	.C2V_12 (C2V_180_823),
	.C2V_13 (C2V_180_904),
	.C2V_14 (C2V_180_918),
	.C2V_15 (C2V_180_1001),
	.C2V_16 (C2V_180_1020),
	.C2V_17 (C2V_180_1084),
	.C2V_18 (C2V_180_1134),
	.C2V_19 (C2V_180_1331),
	.C2V_20 (C2V_180_1332),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU181 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_35_181),
	.V2C_2 (V2C_71_181),
	.V2C_3 (V2C_139_181),
	.V2C_4 (V2C_152_181),
	.V2C_5 (V2C_214_181),
	.V2C_6 (V2C_257_181),
	.V2C_7 (V2C_357_181),
	.V2C_8 (V2C_411_181),
	.V2C_9 (V2C_508_181),
	.V2C_10 (V2C_744_181),
	.V2C_11 (V2C_792_181),
	.V2C_12 (V2C_840_181),
	.V2C_13 (V2C_881_181),
	.V2C_14 (V2C_922_181),
	.V2C_15 (V2C_1004_181),
	.V2C_16 (V2C_1043_181),
	.V2C_17 (V2C_1069_181),
	.V2C_18 (V2C_1128_181),
	.V2C_19 (V2C_1332_181),
	.V2C_20 (V2C_1333_181),
	.C2V_1 (C2V_181_35),
	.C2V_2 (C2V_181_71),
	.C2V_3 (C2V_181_139),
	.C2V_4 (C2V_181_152),
	.C2V_5 (C2V_181_214),
	.C2V_6 (C2V_181_257),
	.C2V_7 (C2V_181_357),
	.C2V_8 (C2V_181_411),
	.C2V_9 (C2V_181_508),
	.C2V_10 (C2V_181_744),
	.C2V_11 (C2V_181_792),
	.C2V_12 (C2V_181_840),
	.C2V_13 (C2V_181_881),
	.C2V_14 (C2V_181_922),
	.C2V_15 (C2V_181_1004),
	.C2V_16 (C2V_181_1043),
	.C2V_17 (C2V_181_1069),
	.C2V_18 (C2V_181_1128),
	.C2V_19 (C2V_181_1332),
	.C2V_20 (C2V_181_1333),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU182 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_44_182),
	.V2C_2 (V2C_93_182),
	.V2C_3 (V2C_101_182),
	.V2C_4 (V2C_149_182),
	.V2C_5 (V2C_226_182),
	.V2C_6 (V2C_247_182),
	.V2C_7 (V2C_298_182),
	.V2C_8 (V2C_405_182),
	.V2C_9 (V2C_494_182),
	.V2C_10 (V2C_654_182),
	.V2C_11 (V2C_715_182),
	.V2C_12 (V2C_835_182),
	.V2C_13 (V2C_877_182),
	.V2C_14 (V2C_940_182),
	.V2C_15 (V2C_971_182),
	.V2C_16 (V2C_1051_182),
	.V2C_17 (V2C_1070_182),
	.V2C_18 (V2C_1149_182),
	.V2C_19 (V2C_1333_182),
	.V2C_20 (V2C_1334_182),
	.C2V_1 (C2V_182_44),
	.C2V_2 (C2V_182_93),
	.C2V_3 (C2V_182_101),
	.C2V_4 (C2V_182_149),
	.C2V_5 (C2V_182_226),
	.C2V_6 (C2V_182_247),
	.C2V_7 (C2V_182_298),
	.C2V_8 (C2V_182_405),
	.C2V_9 (C2V_182_494),
	.C2V_10 (C2V_182_654),
	.C2V_11 (C2V_182_715),
	.C2V_12 (C2V_182_835),
	.C2V_13 (C2V_182_877),
	.C2V_14 (C2V_182_940),
	.C2V_15 (C2V_182_971),
	.C2V_16 (C2V_182_1051),
	.C2V_17 (C2V_182_1070),
	.C2V_18 (C2V_182_1149),
	.C2V_19 (C2V_182_1333),
	.C2V_20 (C2V_182_1334),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU183 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_39_183),
	.V2C_2 (V2C_66_183),
	.V2C_3 (V2C_131_183),
	.V2C_4 (V2C_165_183),
	.V2C_5 (V2C_231_183),
	.V2C_6 (V2C_250_183),
	.V2C_7 (V2C_347_183),
	.V2C_8 (V2C_402_183),
	.V2C_9 (V2C_561_183),
	.V2C_10 (V2C_618_183),
	.V2C_11 (V2C_646_183),
	.V2C_12 (V2C_750_183),
	.V2C_13 (V2C_881_183),
	.V2C_14 (V2C_925_183),
	.V2C_15 (V2C_998_183),
	.V2C_16 (V2C_1010_183),
	.V2C_17 (V2C_1088_183),
	.V2C_18 (V2C_1133_183),
	.V2C_19 (V2C_1334_183),
	.V2C_20 (V2C_1335_183),
	.C2V_1 (C2V_183_39),
	.C2V_2 (C2V_183_66),
	.C2V_3 (C2V_183_131),
	.C2V_4 (C2V_183_165),
	.C2V_5 (C2V_183_231),
	.C2V_6 (C2V_183_250),
	.C2V_7 (C2V_183_347),
	.C2V_8 (C2V_183_402),
	.C2V_9 (C2V_183_561),
	.C2V_10 (C2V_183_618),
	.C2V_11 (C2V_183_646),
	.C2V_12 (C2V_183_750),
	.C2V_13 (C2V_183_881),
	.C2V_14 (C2V_183_925),
	.C2V_15 (C2V_183_998),
	.C2V_16 (C2V_183_1010),
	.C2V_17 (C2V_183_1088),
	.C2V_18 (C2V_183_1133),
	.C2V_19 (C2V_183_1334),
	.C2V_20 (C2V_183_1335),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU184 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_10_184),
	.V2C_2 (V2C_69_184),
	.V2C_3 (V2C_108_184),
	.V2C_4 (V2C_164_184),
	.V2C_5 (V2C_229_184),
	.V2C_6 (V2C_283_184),
	.V2C_7 (V2C_459_184),
	.V2C_8 (V2C_499_184),
	.V2C_9 (V2C_535_184),
	.V2C_10 (V2C_597_184),
	.V2C_11 (V2C_670_184),
	.V2C_12 (V2C_716_184),
	.V2C_13 (V2C_885_184),
	.V2C_14 (V2C_957_184),
	.V2C_15 (V2C_993_184),
	.V2C_16 (V2C_1023_184),
	.V2C_17 (V2C_1098_184),
	.V2C_18 (V2C_1114_184),
	.V2C_19 (V2C_1335_184),
	.V2C_20 (V2C_1336_184),
	.C2V_1 (C2V_184_10),
	.C2V_2 (C2V_184_69),
	.C2V_3 (C2V_184_108),
	.C2V_4 (C2V_184_164),
	.C2V_5 (C2V_184_229),
	.C2V_6 (C2V_184_283),
	.C2V_7 (C2V_184_459),
	.C2V_8 (C2V_184_499),
	.C2V_9 (C2V_184_535),
	.C2V_10 (C2V_184_597),
	.C2V_11 (C2V_184_670),
	.C2V_12 (C2V_184_716),
	.C2V_13 (C2V_184_885),
	.C2V_14 (C2V_184_957),
	.C2V_15 (C2V_184_993),
	.C2V_16 (C2V_184_1023),
	.C2V_17 (C2V_184_1098),
	.C2V_18 (C2V_184_1114),
	.C2V_19 (C2V_184_1335),
	.C2V_20 (C2V_184_1336),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU185 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_29_185),
	.V2C_2 (V2C_87_185),
	.V2C_3 (V2C_122_185),
	.V2C_4 (V2C_145_185),
	.V2C_5 (V2C_209_185),
	.V2C_6 (V2C_275_185),
	.V2C_7 (V2C_324_185),
	.V2C_8 (V2C_343_185),
	.V2C_9 (V2C_470_185),
	.V2C_10 (V2C_704_185),
	.V2C_11 (V2C_768_185),
	.V2C_12 (V2C_774_185),
	.V2C_13 (V2C_900_185),
	.V2C_14 (V2C_948_185),
	.V2C_15 (V2C_991_185),
	.V2C_16 (V2C_1043_185),
	.V2C_17 (V2C_1092_185),
	.V2C_18 (V2C_1140_185),
	.V2C_19 (V2C_1336_185),
	.V2C_20 (V2C_1337_185),
	.C2V_1 (C2V_185_29),
	.C2V_2 (C2V_185_87),
	.C2V_3 (C2V_185_122),
	.C2V_4 (C2V_185_145),
	.C2V_5 (C2V_185_209),
	.C2V_6 (C2V_185_275),
	.C2V_7 (C2V_185_324),
	.C2V_8 (C2V_185_343),
	.C2V_9 (C2V_185_470),
	.C2V_10 (C2V_185_704),
	.C2V_11 (C2V_185_768),
	.C2V_12 (C2V_185_774),
	.C2V_13 (C2V_185_900),
	.C2V_14 (C2V_185_948),
	.C2V_15 (C2V_185_991),
	.C2V_16 (C2V_185_1043),
	.C2V_17 (C2V_185_1092),
	.C2V_18 (C2V_185_1140),
	.C2V_19 (C2V_185_1336),
	.C2V_20 (C2V_185_1337),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU186 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_12_186),
	.V2C_2 (V2C_84_186),
	.V2C_3 (V2C_124_186),
	.V2C_4 (V2C_192_186),
	.V2C_5 (V2C_226_186),
	.V2C_6 (V2C_257_186),
	.V2C_7 (V2C_310_186),
	.V2C_8 (V2C_462_186),
	.V2C_9 (V2C_559_186),
	.V2C_10 (V2C_592_186),
	.V2C_11 (V2C_796_186),
	.V2C_12 (V2C_824_186),
	.V2C_13 (V2C_905_186),
	.V2C_14 (V2C_919_186),
	.V2C_15 (V2C_1002_186),
	.V2C_16 (V2C_1021_186),
	.V2C_17 (V2C_1085_186),
	.V2C_18 (V2C_1135_186),
	.V2C_19 (V2C_1337_186),
	.V2C_20 (V2C_1338_186),
	.C2V_1 (C2V_186_12),
	.C2V_2 (C2V_186_84),
	.C2V_3 (C2V_186_124),
	.C2V_4 (C2V_186_192),
	.C2V_5 (C2V_186_226),
	.C2V_6 (C2V_186_257),
	.C2V_7 (C2V_186_310),
	.C2V_8 (C2V_186_462),
	.C2V_9 (C2V_186_559),
	.C2V_10 (C2V_186_592),
	.C2V_11 (C2V_186_796),
	.C2V_12 (C2V_186_824),
	.C2V_13 (C2V_186_905),
	.C2V_14 (C2V_186_919),
	.C2V_15 (C2V_186_1002),
	.C2V_16 (C2V_186_1021),
	.C2V_17 (C2V_186_1085),
	.C2V_18 (C2V_186_1135),
	.C2V_19 (C2V_186_1337),
	.C2V_20 (C2V_186_1338),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU187 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_36_187),
	.V2C_2 (V2C_72_187),
	.V2C_3 (V2C_140_187),
	.V2C_4 (V2C_153_187),
	.V2C_5 (V2C_215_187),
	.V2C_6 (V2C_258_187),
	.V2C_7 (V2C_358_187),
	.V2C_8 (V2C_412_187),
	.V2C_9 (V2C_509_187),
	.V2C_10 (V2C_745_187),
	.V2C_11 (V2C_793_187),
	.V2C_12 (V2C_841_187),
	.V2C_13 (V2C_882_187),
	.V2C_14 (V2C_923_187),
	.V2C_15 (V2C_1005_187),
	.V2C_16 (V2C_1044_187),
	.V2C_17 (V2C_1070_187),
	.V2C_18 (V2C_1129_187),
	.V2C_19 (V2C_1338_187),
	.V2C_20 (V2C_1339_187),
	.C2V_1 (C2V_187_36),
	.C2V_2 (C2V_187_72),
	.C2V_3 (C2V_187_140),
	.C2V_4 (C2V_187_153),
	.C2V_5 (C2V_187_215),
	.C2V_6 (C2V_187_258),
	.C2V_7 (C2V_187_358),
	.C2V_8 (C2V_187_412),
	.C2V_9 (C2V_187_509),
	.C2V_10 (C2V_187_745),
	.C2V_11 (C2V_187_793),
	.C2V_12 (C2V_187_841),
	.C2V_13 (C2V_187_882),
	.C2V_14 (C2V_187_923),
	.C2V_15 (C2V_187_1005),
	.C2V_16 (C2V_187_1044),
	.C2V_17 (C2V_187_1070),
	.C2V_18 (C2V_187_1129),
	.C2V_19 (C2V_187_1338),
	.C2V_20 (C2V_187_1339),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU188 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_45_188),
	.V2C_2 (V2C_94_188),
	.V2C_3 (V2C_102_188),
	.V2C_4 (V2C_150_188),
	.V2C_5 (V2C_227_188),
	.V2C_6 (V2C_248_188),
	.V2C_7 (V2C_299_188),
	.V2C_8 (V2C_406_188),
	.V2C_9 (V2C_495_188),
	.V2C_10 (V2C_655_188),
	.V2C_11 (V2C_716_188),
	.V2C_12 (V2C_836_188),
	.V2C_13 (V2C_878_188),
	.V2C_14 (V2C_941_188),
	.V2C_15 (V2C_972_188),
	.V2C_16 (V2C_1052_188),
	.V2C_17 (V2C_1071_188),
	.V2C_18 (V2C_1150_188),
	.V2C_19 (V2C_1339_188),
	.V2C_20 (V2C_1340_188),
	.C2V_1 (C2V_188_45),
	.C2V_2 (C2V_188_94),
	.C2V_3 (C2V_188_102),
	.C2V_4 (C2V_188_150),
	.C2V_5 (C2V_188_227),
	.C2V_6 (C2V_188_248),
	.C2V_7 (C2V_188_299),
	.C2V_8 (C2V_188_406),
	.C2V_9 (C2V_188_495),
	.C2V_10 (C2V_188_655),
	.C2V_11 (C2V_188_716),
	.C2V_12 (C2V_188_836),
	.C2V_13 (C2V_188_878),
	.C2V_14 (C2V_188_941),
	.C2V_15 (C2V_188_972),
	.C2V_16 (C2V_188_1052),
	.C2V_17 (C2V_188_1071),
	.C2V_18 (C2V_188_1150),
	.C2V_19 (C2V_188_1339),
	.C2V_20 (C2V_188_1340),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU189 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_40_189),
	.V2C_2 (V2C_67_189),
	.V2C_3 (V2C_132_189),
	.V2C_4 (V2C_166_189),
	.V2C_5 (V2C_232_189),
	.V2C_6 (V2C_251_189),
	.V2C_7 (V2C_348_189),
	.V2C_8 (V2C_403_189),
	.V2C_9 (V2C_562_189),
	.V2C_10 (V2C_619_189),
	.V2C_11 (V2C_647_189),
	.V2C_12 (V2C_751_189),
	.V2C_13 (V2C_882_189),
	.V2C_14 (V2C_926_189),
	.V2C_15 (V2C_999_189),
	.V2C_16 (V2C_1011_189),
	.V2C_17 (V2C_1089_189),
	.V2C_18 (V2C_1134_189),
	.V2C_19 (V2C_1340_189),
	.V2C_20 (V2C_1341_189),
	.C2V_1 (C2V_189_40),
	.C2V_2 (C2V_189_67),
	.C2V_3 (C2V_189_132),
	.C2V_4 (C2V_189_166),
	.C2V_5 (C2V_189_232),
	.C2V_6 (C2V_189_251),
	.C2V_7 (C2V_189_348),
	.C2V_8 (C2V_189_403),
	.C2V_9 (C2V_189_562),
	.C2V_10 (C2V_189_619),
	.C2V_11 (C2V_189_647),
	.C2V_12 (C2V_189_751),
	.C2V_13 (C2V_189_882),
	.C2V_14 (C2V_189_926),
	.C2V_15 (C2V_189_999),
	.C2V_16 (C2V_189_1011),
	.C2V_17 (C2V_189_1089),
	.C2V_18 (C2V_189_1134),
	.C2V_19 (C2V_189_1340),
	.C2V_20 (C2V_189_1341),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU190 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_11_190),
	.V2C_2 (V2C_70_190),
	.V2C_3 (V2C_109_190),
	.V2C_4 (V2C_165_190),
	.V2C_5 (V2C_230_190),
	.V2C_6 (V2C_284_190),
	.V2C_7 (V2C_460_190),
	.V2C_8 (V2C_500_190),
	.V2C_9 (V2C_536_190),
	.V2C_10 (V2C_598_190),
	.V2C_11 (V2C_671_190),
	.V2C_12 (V2C_717_190),
	.V2C_13 (V2C_886_190),
	.V2C_14 (V2C_958_190),
	.V2C_15 (V2C_994_190),
	.V2C_16 (V2C_1024_190),
	.V2C_17 (V2C_1099_190),
	.V2C_18 (V2C_1115_190),
	.V2C_19 (V2C_1341_190),
	.V2C_20 (V2C_1342_190),
	.C2V_1 (C2V_190_11),
	.C2V_2 (C2V_190_70),
	.C2V_3 (C2V_190_109),
	.C2V_4 (C2V_190_165),
	.C2V_5 (C2V_190_230),
	.C2V_6 (C2V_190_284),
	.C2V_7 (C2V_190_460),
	.C2V_8 (C2V_190_500),
	.C2V_9 (C2V_190_536),
	.C2V_10 (C2V_190_598),
	.C2V_11 (C2V_190_671),
	.C2V_12 (C2V_190_717),
	.C2V_13 (C2V_190_886),
	.C2V_14 (C2V_190_958),
	.C2V_15 (C2V_190_994),
	.C2V_16 (C2V_190_1024),
	.C2V_17 (C2V_190_1099),
	.C2V_18 (C2V_190_1115),
	.C2V_19 (C2V_190_1341),
	.C2V_20 (C2V_190_1342),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU191 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_30_191),
	.V2C_2 (V2C_88_191),
	.V2C_3 (V2C_123_191),
	.V2C_4 (V2C_146_191),
	.V2C_5 (V2C_210_191),
	.V2C_6 (V2C_276_191),
	.V2C_7 (V2C_325_191),
	.V2C_8 (V2C_344_191),
	.V2C_9 (V2C_471_191),
	.V2C_10 (V2C_705_191),
	.V2C_11 (V2C_721_191),
	.V2C_12 (V2C_775_191),
	.V2C_13 (V2C_901_191),
	.V2C_14 (V2C_949_191),
	.V2C_15 (V2C_992_191),
	.V2C_16 (V2C_1044_191),
	.V2C_17 (V2C_1093_191),
	.V2C_18 (V2C_1141_191),
	.V2C_19 (V2C_1342_191),
	.V2C_20 (V2C_1343_191),
	.C2V_1 (C2V_191_30),
	.C2V_2 (C2V_191_88),
	.C2V_3 (C2V_191_123),
	.C2V_4 (C2V_191_146),
	.C2V_5 (C2V_191_210),
	.C2V_6 (C2V_191_276),
	.C2V_7 (C2V_191_325),
	.C2V_8 (C2V_191_344),
	.C2V_9 (C2V_191_471),
	.C2V_10 (C2V_191_705),
	.C2V_11 (C2V_191_721),
	.C2V_12 (C2V_191_775),
	.C2V_13 (C2V_191_901),
	.C2V_14 (C2V_191_949),
	.C2V_15 (C2V_191_992),
	.C2V_16 (C2V_191_1044),
	.C2V_17 (C2V_191_1093),
	.C2V_18 (C2V_191_1141),
	.C2V_19 (C2V_191_1342),
	.C2V_20 (C2V_191_1343),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU192 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_13_192),
	.V2C_2 (V2C_85_192),
	.V2C_3 (V2C_125_192),
	.V2C_4 (V2C_145_192),
	.V2C_5 (V2C_227_192),
	.V2C_6 (V2C_258_192),
	.V2C_7 (V2C_311_192),
	.V2C_8 (V2C_463_192),
	.V2C_9 (V2C_560_192),
	.V2C_10 (V2C_593_192),
	.V2C_11 (V2C_797_192),
	.V2C_12 (V2C_825_192),
	.V2C_13 (V2C_906_192),
	.V2C_14 (V2C_920_192),
	.V2C_15 (V2C_1003_192),
	.V2C_16 (V2C_1022_192),
	.V2C_17 (V2C_1086_192),
	.V2C_18 (V2C_1136_192),
	.V2C_19 (V2C_1343_192),
	.V2C_20 (V2C_1344_192),
	.C2V_1 (C2V_192_13),
	.C2V_2 (C2V_192_85),
	.C2V_3 (C2V_192_125),
	.C2V_4 (C2V_192_145),
	.C2V_5 (C2V_192_227),
	.C2V_6 (C2V_192_258),
	.C2V_7 (C2V_192_311),
	.C2V_8 (C2V_192_463),
	.C2V_9 (C2V_192_560),
	.C2V_10 (C2V_192_593),
	.C2V_11 (C2V_192_797),
	.C2V_12 (C2V_192_825),
	.C2V_13 (C2V_192_906),
	.C2V_14 (C2V_192_920),
	.C2V_15 (C2V_192_1003),
	.C2V_16 (C2V_192_1022),
	.C2V_17 (C2V_192_1086),
	.C2V_18 (C2V_192_1136),
	.C2V_19 (C2V_192_1343),
	.C2V_20 (C2V_192_1344),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU193 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_37_193),
	.V2C_2 (V2C_73_193),
	.V2C_3 (V2C_141_193),
	.V2C_4 (V2C_154_193),
	.V2C_5 (V2C_216_193),
	.V2C_6 (V2C_259_193),
	.V2C_7 (V2C_359_193),
	.V2C_8 (V2C_413_193),
	.V2C_9 (V2C_510_193),
	.V2C_10 (V2C_746_193),
	.V2C_11 (V2C_794_193),
	.V2C_12 (V2C_842_193),
	.V2C_13 (V2C_883_193),
	.V2C_14 (V2C_924_193),
	.V2C_15 (V2C_1006_193),
	.V2C_16 (V2C_1045_193),
	.V2C_17 (V2C_1071_193),
	.V2C_18 (V2C_1130_193),
	.V2C_19 (V2C_1344_193),
	.V2C_20 (V2C_1345_193),
	.C2V_1 (C2V_193_37),
	.C2V_2 (C2V_193_73),
	.C2V_3 (C2V_193_141),
	.C2V_4 (C2V_193_154),
	.C2V_5 (C2V_193_216),
	.C2V_6 (C2V_193_259),
	.C2V_7 (C2V_193_359),
	.C2V_8 (C2V_193_413),
	.C2V_9 (C2V_193_510),
	.C2V_10 (C2V_193_746),
	.C2V_11 (C2V_193_794),
	.C2V_12 (C2V_193_842),
	.C2V_13 (C2V_193_883),
	.C2V_14 (C2V_193_924),
	.C2V_15 (C2V_193_1006),
	.C2V_16 (C2V_193_1045),
	.C2V_17 (C2V_193_1071),
	.C2V_18 (C2V_193_1130),
	.C2V_19 (C2V_193_1344),
	.C2V_20 (C2V_193_1345),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU194 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_46_194),
	.V2C_2 (V2C_95_194),
	.V2C_3 (V2C_103_194),
	.V2C_4 (V2C_151_194),
	.V2C_5 (V2C_228_194),
	.V2C_6 (V2C_249_194),
	.V2C_7 (V2C_300_194),
	.V2C_8 (V2C_407_194),
	.V2C_9 (V2C_496_194),
	.V2C_10 (V2C_656_194),
	.V2C_11 (V2C_717_194),
	.V2C_12 (V2C_837_194),
	.V2C_13 (V2C_879_194),
	.V2C_14 (V2C_942_194),
	.V2C_15 (V2C_973_194),
	.V2C_16 (V2C_1053_194),
	.V2C_17 (V2C_1072_194),
	.V2C_18 (V2C_1151_194),
	.V2C_19 (V2C_1345_194),
	.V2C_20 (V2C_1346_194),
	.C2V_1 (C2V_194_46),
	.C2V_2 (C2V_194_95),
	.C2V_3 (C2V_194_103),
	.C2V_4 (C2V_194_151),
	.C2V_5 (C2V_194_228),
	.C2V_6 (C2V_194_249),
	.C2V_7 (C2V_194_300),
	.C2V_8 (C2V_194_407),
	.C2V_9 (C2V_194_496),
	.C2V_10 (C2V_194_656),
	.C2V_11 (C2V_194_717),
	.C2V_12 (C2V_194_837),
	.C2V_13 (C2V_194_879),
	.C2V_14 (C2V_194_942),
	.C2V_15 (C2V_194_973),
	.C2V_16 (C2V_194_1053),
	.C2V_17 (C2V_194_1072),
	.C2V_18 (C2V_194_1151),
	.C2V_19 (C2V_194_1345),
	.C2V_20 (C2V_194_1346),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU195 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_41_195),
	.V2C_2 (V2C_68_195),
	.V2C_3 (V2C_133_195),
	.V2C_4 (V2C_167_195),
	.V2C_5 (V2C_233_195),
	.V2C_6 (V2C_252_195),
	.V2C_7 (V2C_349_195),
	.V2C_8 (V2C_404_195),
	.V2C_9 (V2C_563_195),
	.V2C_10 (V2C_620_195),
	.V2C_11 (V2C_648_195),
	.V2C_12 (V2C_752_195),
	.V2C_13 (V2C_883_195),
	.V2C_14 (V2C_927_195),
	.V2C_15 (V2C_1000_195),
	.V2C_16 (V2C_1012_195),
	.V2C_17 (V2C_1090_195),
	.V2C_18 (V2C_1135_195),
	.V2C_19 (V2C_1346_195),
	.V2C_20 (V2C_1347_195),
	.C2V_1 (C2V_195_41),
	.C2V_2 (C2V_195_68),
	.C2V_3 (C2V_195_133),
	.C2V_4 (C2V_195_167),
	.C2V_5 (C2V_195_233),
	.C2V_6 (C2V_195_252),
	.C2V_7 (C2V_195_349),
	.C2V_8 (C2V_195_404),
	.C2V_9 (C2V_195_563),
	.C2V_10 (C2V_195_620),
	.C2V_11 (C2V_195_648),
	.C2V_12 (C2V_195_752),
	.C2V_13 (C2V_195_883),
	.C2V_14 (C2V_195_927),
	.C2V_15 (C2V_195_1000),
	.C2V_16 (C2V_195_1012),
	.C2V_17 (C2V_195_1090),
	.C2V_18 (C2V_195_1135),
	.C2V_19 (C2V_195_1346),
	.C2V_20 (C2V_195_1347),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU196 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_12_196),
	.V2C_2 (V2C_71_196),
	.V2C_3 (V2C_110_196),
	.V2C_4 (V2C_166_196),
	.V2C_5 (V2C_231_196),
	.V2C_6 (V2C_285_196),
	.V2C_7 (V2C_461_196),
	.V2C_8 (V2C_501_196),
	.V2C_9 (V2C_537_196),
	.V2C_10 (V2C_599_196),
	.V2C_11 (V2C_672_196),
	.V2C_12 (V2C_718_196),
	.V2C_13 (V2C_887_196),
	.V2C_14 (V2C_959_196),
	.V2C_15 (V2C_995_196),
	.V2C_16 (V2C_1025_196),
	.V2C_17 (V2C_1100_196),
	.V2C_18 (V2C_1116_196),
	.V2C_19 (V2C_1347_196),
	.V2C_20 (V2C_1348_196),
	.C2V_1 (C2V_196_12),
	.C2V_2 (C2V_196_71),
	.C2V_3 (C2V_196_110),
	.C2V_4 (C2V_196_166),
	.C2V_5 (C2V_196_231),
	.C2V_6 (C2V_196_285),
	.C2V_7 (C2V_196_461),
	.C2V_8 (C2V_196_501),
	.C2V_9 (C2V_196_537),
	.C2V_10 (C2V_196_599),
	.C2V_11 (C2V_196_672),
	.C2V_12 (C2V_196_718),
	.C2V_13 (C2V_196_887),
	.C2V_14 (C2V_196_959),
	.C2V_15 (C2V_196_995),
	.C2V_16 (C2V_196_1025),
	.C2V_17 (C2V_196_1100),
	.C2V_18 (C2V_196_1116),
	.C2V_19 (C2V_196_1347),
	.C2V_20 (C2V_196_1348),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU197 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_31_197),
	.V2C_2 (V2C_89_197),
	.V2C_3 (V2C_124_197),
	.V2C_4 (V2C_147_197),
	.V2C_5 (V2C_211_197),
	.V2C_6 (V2C_277_197),
	.V2C_7 (V2C_326_197),
	.V2C_8 (V2C_345_197),
	.V2C_9 (V2C_472_197),
	.V2C_10 (V2C_706_197),
	.V2C_11 (V2C_722_197),
	.V2C_12 (V2C_776_197),
	.V2C_13 (V2C_902_197),
	.V2C_14 (V2C_950_197),
	.V2C_15 (V2C_993_197),
	.V2C_16 (V2C_1045_197),
	.V2C_17 (V2C_1094_197),
	.V2C_18 (V2C_1142_197),
	.V2C_19 (V2C_1348_197),
	.V2C_20 (V2C_1349_197),
	.C2V_1 (C2V_197_31),
	.C2V_2 (C2V_197_89),
	.C2V_3 (C2V_197_124),
	.C2V_4 (C2V_197_147),
	.C2V_5 (C2V_197_211),
	.C2V_6 (C2V_197_277),
	.C2V_7 (C2V_197_326),
	.C2V_8 (C2V_197_345),
	.C2V_9 (C2V_197_472),
	.C2V_10 (C2V_197_706),
	.C2V_11 (C2V_197_722),
	.C2V_12 (C2V_197_776),
	.C2V_13 (C2V_197_902),
	.C2V_14 (C2V_197_950),
	.C2V_15 (C2V_197_993),
	.C2V_16 (C2V_197_1045),
	.C2V_17 (C2V_197_1094),
	.C2V_18 (C2V_197_1142),
	.C2V_19 (C2V_197_1348),
	.C2V_20 (C2V_197_1349),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU198 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_14_198),
	.V2C_2 (V2C_86_198),
	.V2C_3 (V2C_126_198),
	.V2C_4 (V2C_146_198),
	.V2C_5 (V2C_228_198),
	.V2C_6 (V2C_259_198),
	.V2C_7 (V2C_312_198),
	.V2C_8 (V2C_464_198),
	.V2C_9 (V2C_561_198),
	.V2C_10 (V2C_594_198),
	.V2C_11 (V2C_798_198),
	.V2C_12 (V2C_826_198),
	.V2C_13 (V2C_907_198),
	.V2C_14 (V2C_921_198),
	.V2C_15 (V2C_1004_198),
	.V2C_16 (V2C_1023_198),
	.V2C_17 (V2C_1087_198),
	.V2C_18 (V2C_1137_198),
	.V2C_19 (V2C_1349_198),
	.V2C_20 (V2C_1350_198),
	.C2V_1 (C2V_198_14),
	.C2V_2 (C2V_198_86),
	.C2V_3 (C2V_198_126),
	.C2V_4 (C2V_198_146),
	.C2V_5 (C2V_198_228),
	.C2V_6 (C2V_198_259),
	.C2V_7 (C2V_198_312),
	.C2V_8 (C2V_198_464),
	.C2V_9 (C2V_198_561),
	.C2V_10 (C2V_198_594),
	.C2V_11 (C2V_198_798),
	.C2V_12 (C2V_198_826),
	.C2V_13 (C2V_198_907),
	.C2V_14 (C2V_198_921),
	.C2V_15 (C2V_198_1004),
	.C2V_16 (C2V_198_1023),
	.C2V_17 (C2V_198_1087),
	.C2V_18 (C2V_198_1137),
	.C2V_19 (C2V_198_1349),
	.C2V_20 (C2V_198_1350),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU199 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_38_199),
	.V2C_2 (V2C_74_199),
	.V2C_3 (V2C_142_199),
	.V2C_4 (V2C_155_199),
	.V2C_5 (V2C_217_199),
	.V2C_6 (V2C_260_199),
	.V2C_7 (V2C_360_199),
	.V2C_8 (V2C_414_199),
	.V2C_9 (V2C_511_199),
	.V2C_10 (V2C_747_199),
	.V2C_11 (V2C_795_199),
	.V2C_12 (V2C_843_199),
	.V2C_13 (V2C_884_199),
	.V2C_14 (V2C_925_199),
	.V2C_15 (V2C_1007_199),
	.V2C_16 (V2C_1046_199),
	.V2C_17 (V2C_1072_199),
	.V2C_18 (V2C_1131_199),
	.V2C_19 (V2C_1350_199),
	.V2C_20 (V2C_1351_199),
	.C2V_1 (C2V_199_38),
	.C2V_2 (C2V_199_74),
	.C2V_3 (C2V_199_142),
	.C2V_4 (C2V_199_155),
	.C2V_5 (C2V_199_217),
	.C2V_6 (C2V_199_260),
	.C2V_7 (C2V_199_360),
	.C2V_8 (C2V_199_414),
	.C2V_9 (C2V_199_511),
	.C2V_10 (C2V_199_747),
	.C2V_11 (C2V_199_795),
	.C2V_12 (C2V_199_843),
	.C2V_13 (C2V_199_884),
	.C2V_14 (C2V_199_925),
	.C2V_15 (C2V_199_1007),
	.C2V_16 (C2V_199_1046),
	.C2V_17 (C2V_199_1072),
	.C2V_18 (C2V_199_1131),
	.C2V_19 (C2V_199_1350),
	.C2V_20 (C2V_199_1351),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU200 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_47_200),
	.V2C_2 (V2C_96_200),
	.V2C_3 (V2C_104_200),
	.V2C_4 (V2C_152_200),
	.V2C_5 (V2C_229_200),
	.V2C_6 (V2C_250_200),
	.V2C_7 (V2C_301_200),
	.V2C_8 (V2C_408_200),
	.V2C_9 (V2C_497_200),
	.V2C_10 (V2C_657_200),
	.V2C_11 (V2C_718_200),
	.V2C_12 (V2C_838_200),
	.V2C_13 (V2C_880_200),
	.V2C_14 (V2C_943_200),
	.V2C_15 (V2C_974_200),
	.V2C_16 (V2C_1054_200),
	.V2C_17 (V2C_1073_200),
	.V2C_18 (V2C_1152_200),
	.V2C_19 (V2C_1351_200),
	.V2C_20 (V2C_1352_200),
	.C2V_1 (C2V_200_47),
	.C2V_2 (C2V_200_96),
	.C2V_3 (C2V_200_104),
	.C2V_4 (C2V_200_152),
	.C2V_5 (C2V_200_229),
	.C2V_6 (C2V_200_250),
	.C2V_7 (C2V_200_301),
	.C2V_8 (C2V_200_408),
	.C2V_9 (C2V_200_497),
	.C2V_10 (C2V_200_657),
	.C2V_11 (C2V_200_718),
	.C2V_12 (C2V_200_838),
	.C2V_13 (C2V_200_880),
	.C2V_14 (C2V_200_943),
	.C2V_15 (C2V_200_974),
	.C2V_16 (C2V_200_1054),
	.C2V_17 (C2V_200_1073),
	.C2V_18 (C2V_200_1152),
	.C2V_19 (C2V_200_1351),
	.C2V_20 (C2V_200_1352),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU201 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_42_201),
	.V2C_2 (V2C_69_201),
	.V2C_3 (V2C_134_201),
	.V2C_4 (V2C_168_201),
	.V2C_5 (V2C_234_201),
	.V2C_6 (V2C_253_201),
	.V2C_7 (V2C_350_201),
	.V2C_8 (V2C_405_201),
	.V2C_9 (V2C_564_201),
	.V2C_10 (V2C_621_201),
	.V2C_11 (V2C_649_201),
	.V2C_12 (V2C_753_201),
	.V2C_13 (V2C_884_201),
	.V2C_14 (V2C_928_201),
	.V2C_15 (V2C_1001_201),
	.V2C_16 (V2C_1013_201),
	.V2C_17 (V2C_1091_201),
	.V2C_18 (V2C_1136_201),
	.V2C_19 (V2C_1352_201),
	.V2C_20 (V2C_1353_201),
	.C2V_1 (C2V_201_42),
	.C2V_2 (C2V_201_69),
	.C2V_3 (C2V_201_134),
	.C2V_4 (C2V_201_168),
	.C2V_5 (C2V_201_234),
	.C2V_6 (C2V_201_253),
	.C2V_7 (C2V_201_350),
	.C2V_8 (C2V_201_405),
	.C2V_9 (C2V_201_564),
	.C2V_10 (C2V_201_621),
	.C2V_11 (C2V_201_649),
	.C2V_12 (C2V_201_753),
	.C2V_13 (C2V_201_884),
	.C2V_14 (C2V_201_928),
	.C2V_15 (C2V_201_1001),
	.C2V_16 (C2V_201_1013),
	.C2V_17 (C2V_201_1091),
	.C2V_18 (C2V_201_1136),
	.C2V_19 (C2V_201_1352),
	.C2V_20 (C2V_201_1353),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU202 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_13_202),
	.V2C_2 (V2C_72_202),
	.V2C_3 (V2C_111_202),
	.V2C_4 (V2C_167_202),
	.V2C_5 (V2C_232_202),
	.V2C_6 (V2C_286_202),
	.V2C_7 (V2C_462_202),
	.V2C_8 (V2C_502_202),
	.V2C_9 (V2C_538_202),
	.V2C_10 (V2C_600_202),
	.V2C_11 (V2C_625_202),
	.V2C_12 (V2C_719_202),
	.V2C_13 (V2C_888_202),
	.V2C_14 (V2C_960_202),
	.V2C_15 (V2C_996_202),
	.V2C_16 (V2C_1026_202),
	.V2C_17 (V2C_1101_202),
	.V2C_18 (V2C_1117_202),
	.V2C_19 (V2C_1353_202),
	.V2C_20 (V2C_1354_202),
	.C2V_1 (C2V_202_13),
	.C2V_2 (C2V_202_72),
	.C2V_3 (C2V_202_111),
	.C2V_4 (C2V_202_167),
	.C2V_5 (C2V_202_232),
	.C2V_6 (C2V_202_286),
	.C2V_7 (C2V_202_462),
	.C2V_8 (C2V_202_502),
	.C2V_9 (C2V_202_538),
	.C2V_10 (C2V_202_600),
	.C2V_11 (C2V_202_625),
	.C2V_12 (C2V_202_719),
	.C2V_13 (C2V_202_888),
	.C2V_14 (C2V_202_960),
	.C2V_15 (C2V_202_996),
	.C2V_16 (C2V_202_1026),
	.C2V_17 (C2V_202_1101),
	.C2V_18 (C2V_202_1117),
	.C2V_19 (C2V_202_1353),
	.C2V_20 (C2V_202_1354),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU203 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_32_203),
	.V2C_2 (V2C_90_203),
	.V2C_3 (V2C_125_203),
	.V2C_4 (V2C_148_203),
	.V2C_5 (V2C_212_203),
	.V2C_6 (V2C_278_203),
	.V2C_7 (V2C_327_203),
	.V2C_8 (V2C_346_203),
	.V2C_9 (V2C_473_203),
	.V2C_10 (V2C_707_203),
	.V2C_11 (V2C_723_203),
	.V2C_12 (V2C_777_203),
	.V2C_13 (V2C_903_203),
	.V2C_14 (V2C_951_203),
	.V2C_15 (V2C_994_203),
	.V2C_16 (V2C_1046_203),
	.V2C_17 (V2C_1095_203),
	.V2C_18 (V2C_1143_203),
	.V2C_19 (V2C_1354_203),
	.V2C_20 (V2C_1355_203),
	.C2V_1 (C2V_203_32),
	.C2V_2 (C2V_203_90),
	.C2V_3 (C2V_203_125),
	.C2V_4 (C2V_203_148),
	.C2V_5 (C2V_203_212),
	.C2V_6 (C2V_203_278),
	.C2V_7 (C2V_203_327),
	.C2V_8 (C2V_203_346),
	.C2V_9 (C2V_203_473),
	.C2V_10 (C2V_203_707),
	.C2V_11 (C2V_203_723),
	.C2V_12 (C2V_203_777),
	.C2V_13 (C2V_203_903),
	.C2V_14 (C2V_203_951),
	.C2V_15 (C2V_203_994),
	.C2V_16 (C2V_203_1046),
	.C2V_17 (C2V_203_1095),
	.C2V_18 (C2V_203_1143),
	.C2V_19 (C2V_203_1354),
	.C2V_20 (C2V_203_1355),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU204 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_15_204),
	.V2C_2 (V2C_87_204),
	.V2C_3 (V2C_127_204),
	.V2C_4 (V2C_147_204),
	.V2C_5 (V2C_229_204),
	.V2C_6 (V2C_260_204),
	.V2C_7 (V2C_313_204),
	.V2C_8 (V2C_465_204),
	.V2C_9 (V2C_562_204),
	.V2C_10 (V2C_595_204),
	.V2C_11 (V2C_799_204),
	.V2C_12 (V2C_827_204),
	.V2C_13 (V2C_908_204),
	.V2C_14 (V2C_922_204),
	.V2C_15 (V2C_1005_204),
	.V2C_16 (V2C_1024_204),
	.V2C_17 (V2C_1088_204),
	.V2C_18 (V2C_1138_204),
	.V2C_19 (V2C_1355_204),
	.V2C_20 (V2C_1356_204),
	.C2V_1 (C2V_204_15),
	.C2V_2 (C2V_204_87),
	.C2V_3 (C2V_204_127),
	.C2V_4 (C2V_204_147),
	.C2V_5 (C2V_204_229),
	.C2V_6 (C2V_204_260),
	.C2V_7 (C2V_204_313),
	.C2V_8 (C2V_204_465),
	.C2V_9 (C2V_204_562),
	.C2V_10 (C2V_204_595),
	.C2V_11 (C2V_204_799),
	.C2V_12 (C2V_204_827),
	.C2V_13 (C2V_204_908),
	.C2V_14 (C2V_204_922),
	.C2V_15 (C2V_204_1005),
	.C2V_16 (C2V_204_1024),
	.C2V_17 (C2V_204_1088),
	.C2V_18 (C2V_204_1138),
	.C2V_19 (C2V_204_1355),
	.C2V_20 (C2V_204_1356),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU205 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_39_205),
	.V2C_2 (V2C_75_205),
	.V2C_3 (V2C_143_205),
	.V2C_4 (V2C_156_205),
	.V2C_5 (V2C_218_205),
	.V2C_6 (V2C_261_205),
	.V2C_7 (V2C_361_205),
	.V2C_8 (V2C_415_205),
	.V2C_9 (V2C_512_205),
	.V2C_10 (V2C_748_205),
	.V2C_11 (V2C_796_205),
	.V2C_12 (V2C_844_205),
	.V2C_13 (V2C_885_205),
	.V2C_14 (V2C_926_205),
	.V2C_15 (V2C_1008_205),
	.V2C_16 (V2C_1047_205),
	.V2C_17 (V2C_1073_205),
	.V2C_18 (V2C_1132_205),
	.V2C_19 (V2C_1356_205),
	.V2C_20 (V2C_1357_205),
	.C2V_1 (C2V_205_39),
	.C2V_2 (C2V_205_75),
	.C2V_3 (C2V_205_143),
	.C2V_4 (C2V_205_156),
	.C2V_5 (C2V_205_218),
	.C2V_6 (C2V_205_261),
	.C2V_7 (C2V_205_361),
	.C2V_8 (C2V_205_415),
	.C2V_9 (C2V_205_512),
	.C2V_10 (C2V_205_748),
	.C2V_11 (C2V_205_796),
	.C2V_12 (C2V_205_844),
	.C2V_13 (C2V_205_885),
	.C2V_14 (C2V_205_926),
	.C2V_15 (C2V_205_1008),
	.C2V_16 (C2V_205_1047),
	.C2V_17 (C2V_205_1073),
	.C2V_18 (C2V_205_1132),
	.C2V_19 (C2V_205_1356),
	.C2V_20 (C2V_205_1357),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU206 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_48_206),
	.V2C_2 (V2C_49_206),
	.V2C_3 (V2C_105_206),
	.V2C_4 (V2C_153_206),
	.V2C_5 (V2C_230_206),
	.V2C_6 (V2C_251_206),
	.V2C_7 (V2C_302_206),
	.V2C_8 (V2C_409_206),
	.V2C_9 (V2C_498_206),
	.V2C_10 (V2C_658_206),
	.V2C_11 (V2C_719_206),
	.V2C_12 (V2C_839_206),
	.V2C_13 (V2C_881_206),
	.V2C_14 (V2C_944_206),
	.V2C_15 (V2C_975_206),
	.V2C_16 (V2C_1055_206),
	.V2C_17 (V2C_1074_206),
	.V2C_18 (V2C_1105_206),
	.V2C_19 (V2C_1357_206),
	.V2C_20 (V2C_1358_206),
	.C2V_1 (C2V_206_48),
	.C2V_2 (C2V_206_49),
	.C2V_3 (C2V_206_105),
	.C2V_4 (C2V_206_153),
	.C2V_5 (C2V_206_230),
	.C2V_6 (C2V_206_251),
	.C2V_7 (C2V_206_302),
	.C2V_8 (C2V_206_409),
	.C2V_9 (C2V_206_498),
	.C2V_10 (C2V_206_658),
	.C2V_11 (C2V_206_719),
	.C2V_12 (C2V_206_839),
	.C2V_13 (C2V_206_881),
	.C2V_14 (C2V_206_944),
	.C2V_15 (C2V_206_975),
	.C2V_16 (C2V_206_1055),
	.C2V_17 (C2V_206_1074),
	.C2V_18 (C2V_206_1105),
	.C2V_19 (C2V_206_1357),
	.C2V_20 (C2V_206_1358),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU207 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_43_207),
	.V2C_2 (V2C_70_207),
	.V2C_3 (V2C_135_207),
	.V2C_4 (V2C_169_207),
	.V2C_5 (V2C_235_207),
	.V2C_6 (V2C_254_207),
	.V2C_7 (V2C_351_207),
	.V2C_8 (V2C_406_207),
	.V2C_9 (V2C_565_207),
	.V2C_10 (V2C_622_207),
	.V2C_11 (V2C_650_207),
	.V2C_12 (V2C_754_207),
	.V2C_13 (V2C_885_207),
	.V2C_14 (V2C_929_207),
	.V2C_15 (V2C_1002_207),
	.V2C_16 (V2C_1014_207),
	.V2C_17 (V2C_1092_207),
	.V2C_18 (V2C_1137_207),
	.V2C_19 (V2C_1358_207),
	.V2C_20 (V2C_1359_207),
	.C2V_1 (C2V_207_43),
	.C2V_2 (C2V_207_70),
	.C2V_3 (C2V_207_135),
	.C2V_4 (C2V_207_169),
	.C2V_5 (C2V_207_235),
	.C2V_6 (C2V_207_254),
	.C2V_7 (C2V_207_351),
	.C2V_8 (C2V_207_406),
	.C2V_9 (C2V_207_565),
	.C2V_10 (C2V_207_622),
	.C2V_11 (C2V_207_650),
	.C2V_12 (C2V_207_754),
	.C2V_13 (C2V_207_885),
	.C2V_14 (C2V_207_929),
	.C2V_15 (C2V_207_1002),
	.C2V_16 (C2V_207_1014),
	.C2V_17 (C2V_207_1092),
	.C2V_18 (C2V_207_1137),
	.C2V_19 (C2V_207_1358),
	.C2V_20 (C2V_207_1359),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU208 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_14_208),
	.V2C_2 (V2C_73_208),
	.V2C_3 (V2C_112_208),
	.V2C_4 (V2C_168_208),
	.V2C_5 (V2C_233_208),
	.V2C_6 (V2C_287_208),
	.V2C_7 (V2C_463_208),
	.V2C_8 (V2C_503_208),
	.V2C_9 (V2C_539_208),
	.V2C_10 (V2C_601_208),
	.V2C_11 (V2C_626_208),
	.V2C_12 (V2C_720_208),
	.V2C_13 (V2C_889_208),
	.V2C_14 (V2C_913_208),
	.V2C_15 (V2C_997_208),
	.V2C_16 (V2C_1027_208),
	.V2C_17 (V2C_1102_208),
	.V2C_18 (V2C_1118_208),
	.V2C_19 (V2C_1359_208),
	.V2C_20 (V2C_1360_208),
	.C2V_1 (C2V_208_14),
	.C2V_2 (C2V_208_73),
	.C2V_3 (C2V_208_112),
	.C2V_4 (C2V_208_168),
	.C2V_5 (C2V_208_233),
	.C2V_6 (C2V_208_287),
	.C2V_7 (C2V_208_463),
	.C2V_8 (C2V_208_503),
	.C2V_9 (C2V_208_539),
	.C2V_10 (C2V_208_601),
	.C2V_11 (C2V_208_626),
	.C2V_12 (C2V_208_720),
	.C2V_13 (C2V_208_889),
	.C2V_14 (C2V_208_913),
	.C2V_15 (C2V_208_997),
	.C2V_16 (C2V_208_1027),
	.C2V_17 (C2V_208_1102),
	.C2V_18 (C2V_208_1118),
	.C2V_19 (C2V_208_1359),
	.C2V_20 (C2V_208_1360),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU209 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_33_209),
	.V2C_2 (V2C_91_209),
	.V2C_3 (V2C_126_209),
	.V2C_4 (V2C_149_209),
	.V2C_5 (V2C_213_209),
	.V2C_6 (V2C_279_209),
	.V2C_7 (V2C_328_209),
	.V2C_8 (V2C_347_209),
	.V2C_9 (V2C_474_209),
	.V2C_10 (V2C_708_209),
	.V2C_11 (V2C_724_209),
	.V2C_12 (V2C_778_209),
	.V2C_13 (V2C_904_209),
	.V2C_14 (V2C_952_209),
	.V2C_15 (V2C_995_209),
	.V2C_16 (V2C_1047_209),
	.V2C_17 (V2C_1096_209),
	.V2C_18 (V2C_1144_209),
	.V2C_19 (V2C_1360_209),
	.V2C_20 (V2C_1361_209),
	.C2V_1 (C2V_209_33),
	.C2V_2 (C2V_209_91),
	.C2V_3 (C2V_209_126),
	.C2V_4 (C2V_209_149),
	.C2V_5 (C2V_209_213),
	.C2V_6 (C2V_209_279),
	.C2V_7 (C2V_209_328),
	.C2V_8 (C2V_209_347),
	.C2V_9 (C2V_209_474),
	.C2V_10 (C2V_209_708),
	.C2V_11 (C2V_209_724),
	.C2V_12 (C2V_209_778),
	.C2V_13 (C2V_209_904),
	.C2V_14 (C2V_209_952),
	.C2V_15 (C2V_209_995),
	.C2V_16 (C2V_209_1047),
	.C2V_17 (C2V_209_1096),
	.C2V_18 (C2V_209_1144),
	.C2V_19 (C2V_209_1360),
	.C2V_20 (C2V_209_1361),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU210 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_16_210),
	.V2C_2 (V2C_88_210),
	.V2C_3 (V2C_128_210),
	.V2C_4 (V2C_148_210),
	.V2C_5 (V2C_230_210),
	.V2C_6 (V2C_261_210),
	.V2C_7 (V2C_314_210),
	.V2C_8 (V2C_466_210),
	.V2C_9 (V2C_563_210),
	.V2C_10 (V2C_596_210),
	.V2C_11 (V2C_800_210),
	.V2C_12 (V2C_828_210),
	.V2C_13 (V2C_909_210),
	.V2C_14 (V2C_923_210),
	.V2C_15 (V2C_1006_210),
	.V2C_16 (V2C_1025_210),
	.V2C_17 (V2C_1089_210),
	.V2C_18 (V2C_1139_210),
	.V2C_19 (V2C_1361_210),
	.V2C_20 (V2C_1362_210),
	.C2V_1 (C2V_210_16),
	.C2V_2 (C2V_210_88),
	.C2V_3 (C2V_210_128),
	.C2V_4 (C2V_210_148),
	.C2V_5 (C2V_210_230),
	.C2V_6 (C2V_210_261),
	.C2V_7 (C2V_210_314),
	.C2V_8 (C2V_210_466),
	.C2V_9 (C2V_210_563),
	.C2V_10 (C2V_210_596),
	.C2V_11 (C2V_210_800),
	.C2V_12 (C2V_210_828),
	.C2V_13 (C2V_210_909),
	.C2V_14 (C2V_210_923),
	.C2V_15 (C2V_210_1006),
	.C2V_16 (C2V_210_1025),
	.C2V_17 (C2V_210_1089),
	.C2V_18 (C2V_210_1139),
	.C2V_19 (C2V_210_1361),
	.C2V_20 (C2V_210_1362),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU211 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_40_211),
	.V2C_2 (V2C_76_211),
	.V2C_3 (V2C_144_211),
	.V2C_4 (V2C_157_211),
	.V2C_5 (V2C_219_211),
	.V2C_6 (V2C_262_211),
	.V2C_7 (V2C_362_211),
	.V2C_8 (V2C_416_211),
	.V2C_9 (V2C_513_211),
	.V2C_10 (V2C_749_211),
	.V2C_11 (V2C_797_211),
	.V2C_12 (V2C_845_211),
	.V2C_13 (V2C_886_211),
	.V2C_14 (V2C_927_211),
	.V2C_15 (V2C_961_211),
	.V2C_16 (V2C_1048_211),
	.V2C_17 (V2C_1074_211),
	.V2C_18 (V2C_1133_211),
	.V2C_19 (V2C_1362_211),
	.V2C_20 (V2C_1363_211),
	.C2V_1 (C2V_211_40),
	.C2V_2 (C2V_211_76),
	.C2V_3 (C2V_211_144),
	.C2V_4 (C2V_211_157),
	.C2V_5 (C2V_211_219),
	.C2V_6 (C2V_211_262),
	.C2V_7 (C2V_211_362),
	.C2V_8 (C2V_211_416),
	.C2V_9 (C2V_211_513),
	.C2V_10 (C2V_211_749),
	.C2V_11 (C2V_211_797),
	.C2V_12 (C2V_211_845),
	.C2V_13 (C2V_211_886),
	.C2V_14 (C2V_211_927),
	.C2V_15 (C2V_211_961),
	.C2V_16 (C2V_211_1048),
	.C2V_17 (C2V_211_1074),
	.C2V_18 (C2V_211_1133),
	.C2V_19 (C2V_211_1362),
	.C2V_20 (C2V_211_1363),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU212 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_1_212),
	.V2C_2 (V2C_50_212),
	.V2C_3 (V2C_106_212),
	.V2C_4 (V2C_154_212),
	.V2C_5 (V2C_231_212),
	.V2C_6 (V2C_252_212),
	.V2C_7 (V2C_303_212),
	.V2C_8 (V2C_410_212),
	.V2C_9 (V2C_499_212),
	.V2C_10 (V2C_659_212),
	.V2C_11 (V2C_720_212),
	.V2C_12 (V2C_840_212),
	.V2C_13 (V2C_882_212),
	.V2C_14 (V2C_945_212),
	.V2C_15 (V2C_976_212),
	.V2C_16 (V2C_1056_212),
	.V2C_17 (V2C_1075_212),
	.V2C_18 (V2C_1106_212),
	.V2C_19 (V2C_1363_212),
	.V2C_20 (V2C_1364_212),
	.C2V_1 (C2V_212_1),
	.C2V_2 (C2V_212_50),
	.C2V_3 (C2V_212_106),
	.C2V_4 (C2V_212_154),
	.C2V_5 (C2V_212_231),
	.C2V_6 (C2V_212_252),
	.C2V_7 (C2V_212_303),
	.C2V_8 (C2V_212_410),
	.C2V_9 (C2V_212_499),
	.C2V_10 (C2V_212_659),
	.C2V_11 (C2V_212_720),
	.C2V_12 (C2V_212_840),
	.C2V_13 (C2V_212_882),
	.C2V_14 (C2V_212_945),
	.C2V_15 (C2V_212_976),
	.C2V_16 (C2V_212_1056),
	.C2V_17 (C2V_212_1075),
	.C2V_18 (C2V_212_1106),
	.C2V_19 (C2V_212_1363),
	.C2V_20 (C2V_212_1364),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU213 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_44_213),
	.V2C_2 (V2C_71_213),
	.V2C_3 (V2C_136_213),
	.V2C_4 (V2C_170_213),
	.V2C_5 (V2C_236_213),
	.V2C_6 (V2C_255_213),
	.V2C_7 (V2C_352_213),
	.V2C_8 (V2C_407_213),
	.V2C_9 (V2C_566_213),
	.V2C_10 (V2C_623_213),
	.V2C_11 (V2C_651_213),
	.V2C_12 (V2C_755_213),
	.V2C_13 (V2C_886_213),
	.V2C_14 (V2C_930_213),
	.V2C_15 (V2C_1003_213),
	.V2C_16 (V2C_1015_213),
	.V2C_17 (V2C_1093_213),
	.V2C_18 (V2C_1138_213),
	.V2C_19 (V2C_1364_213),
	.V2C_20 (V2C_1365_213),
	.C2V_1 (C2V_213_44),
	.C2V_2 (C2V_213_71),
	.C2V_3 (C2V_213_136),
	.C2V_4 (C2V_213_170),
	.C2V_5 (C2V_213_236),
	.C2V_6 (C2V_213_255),
	.C2V_7 (C2V_213_352),
	.C2V_8 (C2V_213_407),
	.C2V_9 (C2V_213_566),
	.C2V_10 (C2V_213_623),
	.C2V_11 (C2V_213_651),
	.C2V_12 (C2V_213_755),
	.C2V_13 (C2V_213_886),
	.C2V_14 (C2V_213_930),
	.C2V_15 (C2V_213_1003),
	.C2V_16 (C2V_213_1015),
	.C2V_17 (C2V_213_1093),
	.C2V_18 (C2V_213_1138),
	.C2V_19 (C2V_213_1364),
	.C2V_20 (C2V_213_1365),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU214 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_15_214),
	.V2C_2 (V2C_74_214),
	.V2C_3 (V2C_113_214),
	.V2C_4 (V2C_169_214),
	.V2C_5 (V2C_234_214),
	.V2C_6 (V2C_288_214),
	.V2C_7 (V2C_464_214),
	.V2C_8 (V2C_504_214),
	.V2C_9 (V2C_540_214),
	.V2C_10 (V2C_602_214),
	.V2C_11 (V2C_627_214),
	.V2C_12 (V2C_673_214),
	.V2C_13 (V2C_890_214),
	.V2C_14 (V2C_914_214),
	.V2C_15 (V2C_998_214),
	.V2C_16 (V2C_1028_214),
	.V2C_17 (V2C_1103_214),
	.V2C_18 (V2C_1119_214),
	.V2C_19 (V2C_1365_214),
	.V2C_20 (V2C_1366_214),
	.C2V_1 (C2V_214_15),
	.C2V_2 (C2V_214_74),
	.C2V_3 (C2V_214_113),
	.C2V_4 (C2V_214_169),
	.C2V_5 (C2V_214_234),
	.C2V_6 (C2V_214_288),
	.C2V_7 (C2V_214_464),
	.C2V_8 (C2V_214_504),
	.C2V_9 (C2V_214_540),
	.C2V_10 (C2V_214_602),
	.C2V_11 (C2V_214_627),
	.C2V_12 (C2V_214_673),
	.C2V_13 (C2V_214_890),
	.C2V_14 (C2V_214_914),
	.C2V_15 (C2V_214_998),
	.C2V_16 (C2V_214_1028),
	.C2V_17 (C2V_214_1103),
	.C2V_18 (C2V_214_1119),
	.C2V_19 (C2V_214_1365),
	.C2V_20 (C2V_214_1366),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU215 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_34_215),
	.V2C_2 (V2C_92_215),
	.V2C_3 (V2C_127_215),
	.V2C_4 (V2C_150_215),
	.V2C_5 (V2C_214_215),
	.V2C_6 (V2C_280_215),
	.V2C_7 (V2C_329_215),
	.V2C_8 (V2C_348_215),
	.V2C_9 (V2C_475_215),
	.V2C_10 (V2C_709_215),
	.V2C_11 (V2C_725_215),
	.V2C_12 (V2C_779_215),
	.V2C_13 (V2C_905_215),
	.V2C_14 (V2C_953_215),
	.V2C_15 (V2C_996_215),
	.V2C_16 (V2C_1048_215),
	.V2C_17 (V2C_1097_215),
	.V2C_18 (V2C_1145_215),
	.V2C_19 (V2C_1366_215),
	.V2C_20 (V2C_1367_215),
	.C2V_1 (C2V_215_34),
	.C2V_2 (C2V_215_92),
	.C2V_3 (C2V_215_127),
	.C2V_4 (C2V_215_150),
	.C2V_5 (C2V_215_214),
	.C2V_6 (C2V_215_280),
	.C2V_7 (C2V_215_329),
	.C2V_8 (C2V_215_348),
	.C2V_9 (C2V_215_475),
	.C2V_10 (C2V_215_709),
	.C2V_11 (C2V_215_725),
	.C2V_12 (C2V_215_779),
	.C2V_13 (C2V_215_905),
	.C2V_14 (C2V_215_953),
	.C2V_15 (C2V_215_996),
	.C2V_16 (C2V_215_1048),
	.C2V_17 (C2V_215_1097),
	.C2V_18 (C2V_215_1145),
	.C2V_19 (C2V_215_1366),
	.C2V_20 (C2V_215_1367),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU216 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_17_216),
	.V2C_2 (V2C_89_216),
	.V2C_3 (V2C_129_216),
	.V2C_4 (V2C_149_216),
	.V2C_5 (V2C_231_216),
	.V2C_6 (V2C_262_216),
	.V2C_7 (V2C_315_216),
	.V2C_8 (V2C_467_216),
	.V2C_9 (V2C_564_216),
	.V2C_10 (V2C_597_216),
	.V2C_11 (V2C_801_216),
	.V2C_12 (V2C_829_216),
	.V2C_13 (V2C_910_216),
	.V2C_14 (V2C_924_216),
	.V2C_15 (V2C_1007_216),
	.V2C_16 (V2C_1026_216),
	.V2C_17 (V2C_1090_216),
	.V2C_18 (V2C_1140_216),
	.V2C_19 (V2C_1367_216),
	.V2C_20 (V2C_1368_216),
	.C2V_1 (C2V_216_17),
	.C2V_2 (C2V_216_89),
	.C2V_3 (C2V_216_129),
	.C2V_4 (C2V_216_149),
	.C2V_5 (C2V_216_231),
	.C2V_6 (C2V_216_262),
	.C2V_7 (C2V_216_315),
	.C2V_8 (C2V_216_467),
	.C2V_9 (C2V_216_564),
	.C2V_10 (C2V_216_597),
	.C2V_11 (C2V_216_801),
	.C2V_12 (C2V_216_829),
	.C2V_13 (C2V_216_910),
	.C2V_14 (C2V_216_924),
	.C2V_15 (C2V_216_1007),
	.C2V_16 (C2V_216_1026),
	.C2V_17 (C2V_216_1090),
	.C2V_18 (C2V_216_1140),
	.C2V_19 (C2V_216_1367),
	.C2V_20 (C2V_216_1368),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU217 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_41_217),
	.V2C_2 (V2C_77_217),
	.V2C_3 (V2C_97_217),
	.V2C_4 (V2C_158_217),
	.V2C_5 (V2C_220_217),
	.V2C_6 (V2C_263_217),
	.V2C_7 (V2C_363_217),
	.V2C_8 (V2C_417_217),
	.V2C_9 (V2C_514_217),
	.V2C_10 (V2C_750_217),
	.V2C_11 (V2C_798_217),
	.V2C_12 (V2C_846_217),
	.V2C_13 (V2C_887_217),
	.V2C_14 (V2C_928_217),
	.V2C_15 (V2C_962_217),
	.V2C_16 (V2C_1049_217),
	.V2C_17 (V2C_1075_217),
	.V2C_18 (V2C_1134_217),
	.V2C_19 (V2C_1368_217),
	.V2C_20 (V2C_1369_217),
	.C2V_1 (C2V_217_41),
	.C2V_2 (C2V_217_77),
	.C2V_3 (C2V_217_97),
	.C2V_4 (C2V_217_158),
	.C2V_5 (C2V_217_220),
	.C2V_6 (C2V_217_263),
	.C2V_7 (C2V_217_363),
	.C2V_8 (C2V_217_417),
	.C2V_9 (C2V_217_514),
	.C2V_10 (C2V_217_750),
	.C2V_11 (C2V_217_798),
	.C2V_12 (C2V_217_846),
	.C2V_13 (C2V_217_887),
	.C2V_14 (C2V_217_928),
	.C2V_15 (C2V_217_962),
	.C2V_16 (C2V_217_1049),
	.C2V_17 (C2V_217_1075),
	.C2V_18 (C2V_217_1134),
	.C2V_19 (C2V_217_1368),
	.C2V_20 (C2V_217_1369),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU218 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_2_218),
	.V2C_2 (V2C_51_218),
	.V2C_3 (V2C_107_218),
	.V2C_4 (V2C_155_218),
	.V2C_5 (V2C_232_218),
	.V2C_6 (V2C_253_218),
	.V2C_7 (V2C_304_218),
	.V2C_8 (V2C_411_218),
	.V2C_9 (V2C_500_218),
	.V2C_10 (V2C_660_218),
	.V2C_11 (V2C_673_218),
	.V2C_12 (V2C_841_218),
	.V2C_13 (V2C_883_218),
	.V2C_14 (V2C_946_218),
	.V2C_15 (V2C_977_218),
	.V2C_16 (V2C_1009_218),
	.V2C_17 (V2C_1076_218),
	.V2C_18 (V2C_1107_218),
	.V2C_19 (V2C_1369_218),
	.V2C_20 (V2C_1370_218),
	.C2V_1 (C2V_218_2),
	.C2V_2 (C2V_218_51),
	.C2V_3 (C2V_218_107),
	.C2V_4 (C2V_218_155),
	.C2V_5 (C2V_218_232),
	.C2V_6 (C2V_218_253),
	.C2V_7 (C2V_218_304),
	.C2V_8 (C2V_218_411),
	.C2V_9 (C2V_218_500),
	.C2V_10 (C2V_218_660),
	.C2V_11 (C2V_218_673),
	.C2V_12 (C2V_218_841),
	.C2V_13 (C2V_218_883),
	.C2V_14 (C2V_218_946),
	.C2V_15 (C2V_218_977),
	.C2V_16 (C2V_218_1009),
	.C2V_17 (C2V_218_1076),
	.C2V_18 (C2V_218_1107),
	.C2V_19 (C2V_218_1369),
	.C2V_20 (C2V_218_1370),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU219 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_45_219),
	.V2C_2 (V2C_72_219),
	.V2C_3 (V2C_137_219),
	.V2C_4 (V2C_171_219),
	.V2C_5 (V2C_237_219),
	.V2C_6 (V2C_256_219),
	.V2C_7 (V2C_353_219),
	.V2C_8 (V2C_408_219),
	.V2C_9 (V2C_567_219),
	.V2C_10 (V2C_624_219),
	.V2C_11 (V2C_652_219),
	.V2C_12 (V2C_756_219),
	.V2C_13 (V2C_887_219),
	.V2C_14 (V2C_931_219),
	.V2C_15 (V2C_1004_219),
	.V2C_16 (V2C_1016_219),
	.V2C_17 (V2C_1094_219),
	.V2C_18 (V2C_1139_219),
	.V2C_19 (V2C_1370_219),
	.V2C_20 (V2C_1371_219),
	.C2V_1 (C2V_219_45),
	.C2V_2 (C2V_219_72),
	.C2V_3 (C2V_219_137),
	.C2V_4 (C2V_219_171),
	.C2V_5 (C2V_219_237),
	.C2V_6 (C2V_219_256),
	.C2V_7 (C2V_219_353),
	.C2V_8 (C2V_219_408),
	.C2V_9 (C2V_219_567),
	.C2V_10 (C2V_219_624),
	.C2V_11 (C2V_219_652),
	.C2V_12 (C2V_219_756),
	.C2V_13 (C2V_219_887),
	.C2V_14 (C2V_219_931),
	.C2V_15 (C2V_219_1004),
	.C2V_16 (C2V_219_1016),
	.C2V_17 (C2V_219_1094),
	.C2V_18 (C2V_219_1139),
	.C2V_19 (C2V_219_1370),
	.C2V_20 (C2V_219_1371),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU220 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_16_220),
	.V2C_2 (V2C_75_220),
	.V2C_3 (V2C_114_220),
	.V2C_4 (V2C_170_220),
	.V2C_5 (V2C_235_220),
	.V2C_6 (V2C_241_220),
	.V2C_7 (V2C_465_220),
	.V2C_8 (V2C_505_220),
	.V2C_9 (V2C_541_220),
	.V2C_10 (V2C_603_220),
	.V2C_11 (V2C_628_220),
	.V2C_12 (V2C_674_220),
	.V2C_13 (V2C_891_220),
	.V2C_14 (V2C_915_220),
	.V2C_15 (V2C_999_220),
	.V2C_16 (V2C_1029_220),
	.V2C_17 (V2C_1104_220),
	.V2C_18 (V2C_1120_220),
	.V2C_19 (V2C_1371_220),
	.V2C_20 (V2C_1372_220),
	.C2V_1 (C2V_220_16),
	.C2V_2 (C2V_220_75),
	.C2V_3 (C2V_220_114),
	.C2V_4 (C2V_220_170),
	.C2V_5 (C2V_220_235),
	.C2V_6 (C2V_220_241),
	.C2V_7 (C2V_220_465),
	.C2V_8 (C2V_220_505),
	.C2V_9 (C2V_220_541),
	.C2V_10 (C2V_220_603),
	.C2V_11 (C2V_220_628),
	.C2V_12 (C2V_220_674),
	.C2V_13 (C2V_220_891),
	.C2V_14 (C2V_220_915),
	.C2V_15 (C2V_220_999),
	.C2V_16 (C2V_220_1029),
	.C2V_17 (C2V_220_1104),
	.C2V_18 (C2V_220_1120),
	.C2V_19 (C2V_220_1371),
	.C2V_20 (C2V_220_1372),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU221 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_35_221),
	.V2C_2 (V2C_93_221),
	.V2C_3 (V2C_128_221),
	.V2C_4 (V2C_151_221),
	.V2C_5 (V2C_215_221),
	.V2C_6 (V2C_281_221),
	.V2C_7 (V2C_330_221),
	.V2C_8 (V2C_349_221),
	.V2C_9 (V2C_476_221),
	.V2C_10 (V2C_710_221),
	.V2C_11 (V2C_726_221),
	.V2C_12 (V2C_780_221),
	.V2C_13 (V2C_906_221),
	.V2C_14 (V2C_954_221),
	.V2C_15 (V2C_997_221),
	.V2C_16 (V2C_1049_221),
	.V2C_17 (V2C_1098_221),
	.V2C_18 (V2C_1146_221),
	.V2C_19 (V2C_1372_221),
	.V2C_20 (V2C_1373_221),
	.C2V_1 (C2V_221_35),
	.C2V_2 (C2V_221_93),
	.C2V_3 (C2V_221_128),
	.C2V_4 (C2V_221_151),
	.C2V_5 (C2V_221_215),
	.C2V_6 (C2V_221_281),
	.C2V_7 (C2V_221_330),
	.C2V_8 (C2V_221_349),
	.C2V_9 (C2V_221_476),
	.C2V_10 (C2V_221_710),
	.C2V_11 (C2V_221_726),
	.C2V_12 (C2V_221_780),
	.C2V_13 (C2V_221_906),
	.C2V_14 (C2V_221_954),
	.C2V_15 (C2V_221_997),
	.C2V_16 (C2V_221_1049),
	.C2V_17 (C2V_221_1098),
	.C2V_18 (C2V_221_1146),
	.C2V_19 (C2V_221_1372),
	.C2V_20 (C2V_221_1373),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU222 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_18_222),
	.V2C_2 (V2C_90_222),
	.V2C_3 (V2C_130_222),
	.V2C_4 (V2C_150_222),
	.V2C_5 (V2C_232_222),
	.V2C_6 (V2C_263_222),
	.V2C_7 (V2C_316_222),
	.V2C_8 (V2C_468_222),
	.V2C_9 (V2C_565_222),
	.V2C_10 (V2C_598_222),
	.V2C_11 (V2C_802_222),
	.V2C_12 (V2C_830_222),
	.V2C_13 (V2C_911_222),
	.V2C_14 (V2C_925_222),
	.V2C_15 (V2C_1008_222),
	.V2C_16 (V2C_1027_222),
	.V2C_17 (V2C_1091_222),
	.V2C_18 (V2C_1141_222),
	.V2C_19 (V2C_1373_222),
	.V2C_20 (V2C_1374_222),
	.C2V_1 (C2V_222_18),
	.C2V_2 (C2V_222_90),
	.C2V_3 (C2V_222_130),
	.C2V_4 (C2V_222_150),
	.C2V_5 (C2V_222_232),
	.C2V_6 (C2V_222_263),
	.C2V_7 (C2V_222_316),
	.C2V_8 (C2V_222_468),
	.C2V_9 (C2V_222_565),
	.C2V_10 (C2V_222_598),
	.C2V_11 (C2V_222_802),
	.C2V_12 (C2V_222_830),
	.C2V_13 (C2V_222_911),
	.C2V_14 (C2V_222_925),
	.C2V_15 (C2V_222_1008),
	.C2V_16 (C2V_222_1027),
	.C2V_17 (C2V_222_1091),
	.C2V_18 (C2V_222_1141),
	.C2V_19 (C2V_222_1373),
	.C2V_20 (C2V_222_1374),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU223 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_42_223),
	.V2C_2 (V2C_78_223),
	.V2C_3 (V2C_98_223),
	.V2C_4 (V2C_159_223),
	.V2C_5 (V2C_221_223),
	.V2C_6 (V2C_264_223),
	.V2C_7 (V2C_364_223),
	.V2C_8 (V2C_418_223),
	.V2C_9 (V2C_515_223),
	.V2C_10 (V2C_751_223),
	.V2C_11 (V2C_799_223),
	.V2C_12 (V2C_847_223),
	.V2C_13 (V2C_888_223),
	.V2C_14 (V2C_929_223),
	.V2C_15 (V2C_963_223),
	.V2C_16 (V2C_1050_223),
	.V2C_17 (V2C_1076_223),
	.V2C_18 (V2C_1135_223),
	.V2C_19 (V2C_1374_223),
	.V2C_20 (V2C_1375_223),
	.C2V_1 (C2V_223_42),
	.C2V_2 (C2V_223_78),
	.C2V_3 (C2V_223_98),
	.C2V_4 (C2V_223_159),
	.C2V_5 (C2V_223_221),
	.C2V_6 (C2V_223_264),
	.C2V_7 (C2V_223_364),
	.C2V_8 (C2V_223_418),
	.C2V_9 (C2V_223_515),
	.C2V_10 (C2V_223_751),
	.C2V_11 (C2V_223_799),
	.C2V_12 (C2V_223_847),
	.C2V_13 (C2V_223_888),
	.C2V_14 (C2V_223_929),
	.C2V_15 (C2V_223_963),
	.C2V_16 (C2V_223_1050),
	.C2V_17 (C2V_223_1076),
	.C2V_18 (C2V_223_1135),
	.C2V_19 (C2V_223_1374),
	.C2V_20 (C2V_223_1375),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU224 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_3_224),
	.V2C_2 (V2C_52_224),
	.V2C_3 (V2C_108_224),
	.V2C_4 (V2C_156_224),
	.V2C_5 (V2C_233_224),
	.V2C_6 (V2C_254_224),
	.V2C_7 (V2C_305_224),
	.V2C_8 (V2C_412_224),
	.V2C_9 (V2C_501_224),
	.V2C_10 (V2C_661_224),
	.V2C_11 (V2C_674_224),
	.V2C_12 (V2C_842_224),
	.V2C_13 (V2C_884_224),
	.V2C_14 (V2C_947_224),
	.V2C_15 (V2C_978_224),
	.V2C_16 (V2C_1010_224),
	.V2C_17 (V2C_1077_224),
	.V2C_18 (V2C_1108_224),
	.V2C_19 (V2C_1375_224),
	.V2C_20 (V2C_1376_224),
	.C2V_1 (C2V_224_3),
	.C2V_2 (C2V_224_52),
	.C2V_3 (C2V_224_108),
	.C2V_4 (C2V_224_156),
	.C2V_5 (C2V_224_233),
	.C2V_6 (C2V_224_254),
	.C2V_7 (C2V_224_305),
	.C2V_8 (C2V_224_412),
	.C2V_9 (C2V_224_501),
	.C2V_10 (C2V_224_661),
	.C2V_11 (C2V_224_674),
	.C2V_12 (C2V_224_842),
	.C2V_13 (C2V_224_884),
	.C2V_14 (C2V_224_947),
	.C2V_15 (C2V_224_978),
	.C2V_16 (C2V_224_1010),
	.C2V_17 (C2V_224_1077),
	.C2V_18 (C2V_224_1108),
	.C2V_19 (C2V_224_1375),
	.C2V_20 (C2V_224_1376),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU225 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_46_225),
	.V2C_2 (V2C_73_225),
	.V2C_3 (V2C_138_225),
	.V2C_4 (V2C_172_225),
	.V2C_5 (V2C_238_225),
	.V2C_6 (V2C_257_225),
	.V2C_7 (V2C_354_225),
	.V2C_8 (V2C_409_225),
	.V2C_9 (V2C_568_225),
	.V2C_10 (V2C_577_225),
	.V2C_11 (V2C_653_225),
	.V2C_12 (V2C_757_225),
	.V2C_13 (V2C_888_225),
	.V2C_14 (V2C_932_225),
	.V2C_15 (V2C_1005_225),
	.V2C_16 (V2C_1017_225),
	.V2C_17 (V2C_1095_225),
	.V2C_18 (V2C_1140_225),
	.V2C_19 (V2C_1376_225),
	.V2C_20 (V2C_1377_225),
	.C2V_1 (C2V_225_46),
	.C2V_2 (C2V_225_73),
	.C2V_3 (C2V_225_138),
	.C2V_4 (C2V_225_172),
	.C2V_5 (C2V_225_238),
	.C2V_6 (C2V_225_257),
	.C2V_7 (C2V_225_354),
	.C2V_8 (C2V_225_409),
	.C2V_9 (C2V_225_568),
	.C2V_10 (C2V_225_577),
	.C2V_11 (C2V_225_653),
	.C2V_12 (C2V_225_757),
	.C2V_13 (C2V_225_888),
	.C2V_14 (C2V_225_932),
	.C2V_15 (C2V_225_1005),
	.C2V_16 (C2V_225_1017),
	.C2V_17 (C2V_225_1095),
	.C2V_18 (C2V_225_1140),
	.C2V_19 (C2V_225_1376),
	.C2V_20 (C2V_225_1377),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU226 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_17_226),
	.V2C_2 (V2C_76_226),
	.V2C_3 (V2C_115_226),
	.V2C_4 (V2C_171_226),
	.V2C_5 (V2C_236_226),
	.V2C_6 (V2C_242_226),
	.V2C_7 (V2C_466_226),
	.V2C_8 (V2C_506_226),
	.V2C_9 (V2C_542_226),
	.V2C_10 (V2C_604_226),
	.V2C_11 (V2C_629_226),
	.V2C_12 (V2C_675_226),
	.V2C_13 (V2C_892_226),
	.V2C_14 (V2C_916_226),
	.V2C_15 (V2C_1000_226),
	.V2C_16 (V2C_1030_226),
	.V2C_17 (V2C_1057_226),
	.V2C_18 (V2C_1121_226),
	.V2C_19 (V2C_1377_226),
	.V2C_20 (V2C_1378_226),
	.C2V_1 (C2V_226_17),
	.C2V_2 (C2V_226_76),
	.C2V_3 (C2V_226_115),
	.C2V_4 (C2V_226_171),
	.C2V_5 (C2V_226_236),
	.C2V_6 (C2V_226_242),
	.C2V_7 (C2V_226_466),
	.C2V_8 (C2V_226_506),
	.C2V_9 (C2V_226_542),
	.C2V_10 (C2V_226_604),
	.C2V_11 (C2V_226_629),
	.C2V_12 (C2V_226_675),
	.C2V_13 (C2V_226_892),
	.C2V_14 (C2V_226_916),
	.C2V_15 (C2V_226_1000),
	.C2V_16 (C2V_226_1030),
	.C2V_17 (C2V_226_1057),
	.C2V_18 (C2V_226_1121),
	.C2V_19 (C2V_226_1377),
	.C2V_20 (C2V_226_1378),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU227 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_36_227),
	.V2C_2 (V2C_94_227),
	.V2C_3 (V2C_129_227),
	.V2C_4 (V2C_152_227),
	.V2C_5 (V2C_216_227),
	.V2C_6 (V2C_282_227),
	.V2C_7 (V2C_331_227),
	.V2C_8 (V2C_350_227),
	.V2C_9 (V2C_477_227),
	.V2C_10 (V2C_711_227),
	.V2C_11 (V2C_727_227),
	.V2C_12 (V2C_781_227),
	.V2C_13 (V2C_907_227),
	.V2C_14 (V2C_955_227),
	.V2C_15 (V2C_998_227),
	.V2C_16 (V2C_1050_227),
	.V2C_17 (V2C_1099_227),
	.V2C_18 (V2C_1147_227),
	.V2C_19 (V2C_1378_227),
	.V2C_20 (V2C_1379_227),
	.C2V_1 (C2V_227_36),
	.C2V_2 (C2V_227_94),
	.C2V_3 (C2V_227_129),
	.C2V_4 (C2V_227_152),
	.C2V_5 (C2V_227_216),
	.C2V_6 (C2V_227_282),
	.C2V_7 (C2V_227_331),
	.C2V_8 (C2V_227_350),
	.C2V_9 (C2V_227_477),
	.C2V_10 (C2V_227_711),
	.C2V_11 (C2V_227_727),
	.C2V_12 (C2V_227_781),
	.C2V_13 (C2V_227_907),
	.C2V_14 (C2V_227_955),
	.C2V_15 (C2V_227_998),
	.C2V_16 (C2V_227_1050),
	.C2V_17 (C2V_227_1099),
	.C2V_18 (C2V_227_1147),
	.C2V_19 (C2V_227_1378),
	.C2V_20 (C2V_227_1379),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU228 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_19_228),
	.V2C_2 (V2C_91_228),
	.V2C_3 (V2C_131_228),
	.V2C_4 (V2C_151_228),
	.V2C_5 (V2C_233_228),
	.V2C_6 (V2C_264_228),
	.V2C_7 (V2C_317_228),
	.V2C_8 (V2C_469_228),
	.V2C_9 (V2C_566_228),
	.V2C_10 (V2C_599_228),
	.V2C_11 (V2C_803_228),
	.V2C_12 (V2C_831_228),
	.V2C_13 (V2C_912_228),
	.V2C_14 (V2C_926_228),
	.V2C_15 (V2C_961_228),
	.V2C_16 (V2C_1028_228),
	.V2C_17 (V2C_1092_228),
	.V2C_18 (V2C_1142_228),
	.V2C_19 (V2C_1379_228),
	.V2C_20 (V2C_1380_228),
	.C2V_1 (C2V_228_19),
	.C2V_2 (C2V_228_91),
	.C2V_3 (C2V_228_131),
	.C2V_4 (C2V_228_151),
	.C2V_5 (C2V_228_233),
	.C2V_6 (C2V_228_264),
	.C2V_7 (C2V_228_317),
	.C2V_8 (C2V_228_469),
	.C2V_9 (C2V_228_566),
	.C2V_10 (C2V_228_599),
	.C2V_11 (C2V_228_803),
	.C2V_12 (C2V_228_831),
	.C2V_13 (C2V_228_912),
	.C2V_14 (C2V_228_926),
	.C2V_15 (C2V_228_961),
	.C2V_16 (C2V_228_1028),
	.C2V_17 (C2V_228_1092),
	.C2V_18 (C2V_228_1142),
	.C2V_19 (C2V_228_1379),
	.C2V_20 (C2V_228_1380),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU229 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_43_229),
	.V2C_2 (V2C_79_229),
	.V2C_3 (V2C_99_229),
	.V2C_4 (V2C_160_229),
	.V2C_5 (V2C_222_229),
	.V2C_6 (V2C_265_229),
	.V2C_7 (V2C_365_229),
	.V2C_8 (V2C_419_229),
	.V2C_9 (V2C_516_229),
	.V2C_10 (V2C_752_229),
	.V2C_11 (V2C_800_229),
	.V2C_12 (V2C_848_229),
	.V2C_13 (V2C_889_229),
	.V2C_14 (V2C_930_229),
	.V2C_15 (V2C_964_229),
	.V2C_16 (V2C_1051_229),
	.V2C_17 (V2C_1077_229),
	.V2C_18 (V2C_1136_229),
	.V2C_19 (V2C_1380_229),
	.V2C_20 (V2C_1381_229),
	.C2V_1 (C2V_229_43),
	.C2V_2 (C2V_229_79),
	.C2V_3 (C2V_229_99),
	.C2V_4 (C2V_229_160),
	.C2V_5 (C2V_229_222),
	.C2V_6 (C2V_229_265),
	.C2V_7 (C2V_229_365),
	.C2V_8 (C2V_229_419),
	.C2V_9 (C2V_229_516),
	.C2V_10 (C2V_229_752),
	.C2V_11 (C2V_229_800),
	.C2V_12 (C2V_229_848),
	.C2V_13 (C2V_229_889),
	.C2V_14 (C2V_229_930),
	.C2V_15 (C2V_229_964),
	.C2V_16 (C2V_229_1051),
	.C2V_17 (C2V_229_1077),
	.C2V_18 (C2V_229_1136),
	.C2V_19 (C2V_229_1380),
	.C2V_20 (C2V_229_1381),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU230 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_4_230),
	.V2C_2 (V2C_53_230),
	.V2C_3 (V2C_109_230),
	.V2C_4 (V2C_157_230),
	.V2C_5 (V2C_234_230),
	.V2C_6 (V2C_255_230),
	.V2C_7 (V2C_306_230),
	.V2C_8 (V2C_413_230),
	.V2C_9 (V2C_502_230),
	.V2C_10 (V2C_662_230),
	.V2C_11 (V2C_675_230),
	.V2C_12 (V2C_843_230),
	.V2C_13 (V2C_885_230),
	.V2C_14 (V2C_948_230),
	.V2C_15 (V2C_979_230),
	.V2C_16 (V2C_1011_230),
	.V2C_17 (V2C_1078_230),
	.V2C_18 (V2C_1109_230),
	.V2C_19 (V2C_1381_230),
	.V2C_20 (V2C_1382_230),
	.C2V_1 (C2V_230_4),
	.C2V_2 (C2V_230_53),
	.C2V_3 (C2V_230_109),
	.C2V_4 (C2V_230_157),
	.C2V_5 (C2V_230_234),
	.C2V_6 (C2V_230_255),
	.C2V_7 (C2V_230_306),
	.C2V_8 (C2V_230_413),
	.C2V_9 (C2V_230_502),
	.C2V_10 (C2V_230_662),
	.C2V_11 (C2V_230_675),
	.C2V_12 (C2V_230_843),
	.C2V_13 (C2V_230_885),
	.C2V_14 (C2V_230_948),
	.C2V_15 (C2V_230_979),
	.C2V_16 (C2V_230_1011),
	.C2V_17 (C2V_230_1078),
	.C2V_18 (C2V_230_1109),
	.C2V_19 (C2V_230_1381),
	.C2V_20 (C2V_230_1382),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU231 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_47_231),
	.V2C_2 (V2C_74_231),
	.V2C_3 (V2C_139_231),
	.V2C_4 (V2C_173_231),
	.V2C_5 (V2C_239_231),
	.V2C_6 (V2C_258_231),
	.V2C_7 (V2C_355_231),
	.V2C_8 (V2C_410_231),
	.V2C_9 (V2C_569_231),
	.V2C_10 (V2C_578_231),
	.V2C_11 (V2C_654_231),
	.V2C_12 (V2C_758_231),
	.V2C_13 (V2C_889_231),
	.V2C_14 (V2C_933_231),
	.V2C_15 (V2C_1006_231),
	.V2C_16 (V2C_1018_231),
	.V2C_17 (V2C_1096_231),
	.V2C_18 (V2C_1141_231),
	.V2C_19 (V2C_1382_231),
	.V2C_20 (V2C_1383_231),
	.C2V_1 (C2V_231_47),
	.C2V_2 (C2V_231_74),
	.C2V_3 (C2V_231_139),
	.C2V_4 (C2V_231_173),
	.C2V_5 (C2V_231_239),
	.C2V_6 (C2V_231_258),
	.C2V_7 (C2V_231_355),
	.C2V_8 (C2V_231_410),
	.C2V_9 (C2V_231_569),
	.C2V_10 (C2V_231_578),
	.C2V_11 (C2V_231_654),
	.C2V_12 (C2V_231_758),
	.C2V_13 (C2V_231_889),
	.C2V_14 (C2V_231_933),
	.C2V_15 (C2V_231_1006),
	.C2V_16 (C2V_231_1018),
	.C2V_17 (C2V_231_1096),
	.C2V_18 (C2V_231_1141),
	.C2V_19 (C2V_231_1382),
	.C2V_20 (C2V_231_1383),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU232 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_18_232),
	.V2C_2 (V2C_77_232),
	.V2C_3 (V2C_116_232),
	.V2C_4 (V2C_172_232),
	.V2C_5 (V2C_237_232),
	.V2C_6 (V2C_243_232),
	.V2C_7 (V2C_467_232),
	.V2C_8 (V2C_507_232),
	.V2C_9 (V2C_543_232),
	.V2C_10 (V2C_605_232),
	.V2C_11 (V2C_630_232),
	.V2C_12 (V2C_676_232),
	.V2C_13 (V2C_893_232),
	.V2C_14 (V2C_917_232),
	.V2C_15 (V2C_1001_232),
	.V2C_16 (V2C_1031_232),
	.V2C_17 (V2C_1058_232),
	.V2C_18 (V2C_1122_232),
	.V2C_19 (V2C_1383_232),
	.V2C_20 (V2C_1384_232),
	.C2V_1 (C2V_232_18),
	.C2V_2 (C2V_232_77),
	.C2V_3 (C2V_232_116),
	.C2V_4 (C2V_232_172),
	.C2V_5 (C2V_232_237),
	.C2V_6 (C2V_232_243),
	.C2V_7 (C2V_232_467),
	.C2V_8 (C2V_232_507),
	.C2V_9 (C2V_232_543),
	.C2V_10 (C2V_232_605),
	.C2V_11 (C2V_232_630),
	.C2V_12 (C2V_232_676),
	.C2V_13 (C2V_232_893),
	.C2V_14 (C2V_232_917),
	.C2V_15 (C2V_232_1001),
	.C2V_16 (C2V_232_1031),
	.C2V_17 (C2V_232_1058),
	.C2V_18 (C2V_232_1122),
	.C2V_19 (C2V_232_1383),
	.C2V_20 (C2V_232_1384),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU233 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_37_233),
	.V2C_2 (V2C_95_233),
	.V2C_3 (V2C_130_233),
	.V2C_4 (V2C_153_233),
	.V2C_5 (V2C_217_233),
	.V2C_6 (V2C_283_233),
	.V2C_7 (V2C_332_233),
	.V2C_8 (V2C_351_233),
	.V2C_9 (V2C_478_233),
	.V2C_10 (V2C_712_233),
	.V2C_11 (V2C_728_233),
	.V2C_12 (V2C_782_233),
	.V2C_13 (V2C_908_233),
	.V2C_14 (V2C_956_233),
	.V2C_15 (V2C_999_233),
	.V2C_16 (V2C_1051_233),
	.V2C_17 (V2C_1100_233),
	.V2C_18 (V2C_1148_233),
	.V2C_19 (V2C_1384_233),
	.V2C_20 (V2C_1385_233),
	.C2V_1 (C2V_233_37),
	.C2V_2 (C2V_233_95),
	.C2V_3 (C2V_233_130),
	.C2V_4 (C2V_233_153),
	.C2V_5 (C2V_233_217),
	.C2V_6 (C2V_233_283),
	.C2V_7 (C2V_233_332),
	.C2V_8 (C2V_233_351),
	.C2V_9 (C2V_233_478),
	.C2V_10 (C2V_233_712),
	.C2V_11 (C2V_233_728),
	.C2V_12 (C2V_233_782),
	.C2V_13 (C2V_233_908),
	.C2V_14 (C2V_233_956),
	.C2V_15 (C2V_233_999),
	.C2V_16 (C2V_233_1051),
	.C2V_17 (C2V_233_1100),
	.C2V_18 (C2V_233_1148),
	.C2V_19 (C2V_233_1384),
	.C2V_20 (C2V_233_1385),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU234 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_20_234),
	.V2C_2 (V2C_92_234),
	.V2C_3 (V2C_132_234),
	.V2C_4 (V2C_152_234),
	.V2C_5 (V2C_234_234),
	.V2C_6 (V2C_265_234),
	.V2C_7 (V2C_318_234),
	.V2C_8 (V2C_470_234),
	.V2C_9 (V2C_567_234),
	.V2C_10 (V2C_600_234),
	.V2C_11 (V2C_804_234),
	.V2C_12 (V2C_832_234),
	.V2C_13 (V2C_865_234),
	.V2C_14 (V2C_927_234),
	.V2C_15 (V2C_962_234),
	.V2C_16 (V2C_1029_234),
	.V2C_17 (V2C_1093_234),
	.V2C_18 (V2C_1143_234),
	.V2C_19 (V2C_1385_234),
	.V2C_20 (V2C_1386_234),
	.C2V_1 (C2V_234_20),
	.C2V_2 (C2V_234_92),
	.C2V_3 (C2V_234_132),
	.C2V_4 (C2V_234_152),
	.C2V_5 (C2V_234_234),
	.C2V_6 (C2V_234_265),
	.C2V_7 (C2V_234_318),
	.C2V_8 (C2V_234_470),
	.C2V_9 (C2V_234_567),
	.C2V_10 (C2V_234_600),
	.C2V_11 (C2V_234_804),
	.C2V_12 (C2V_234_832),
	.C2V_13 (C2V_234_865),
	.C2V_14 (C2V_234_927),
	.C2V_15 (C2V_234_962),
	.C2V_16 (C2V_234_1029),
	.C2V_17 (C2V_234_1093),
	.C2V_18 (C2V_234_1143),
	.C2V_19 (C2V_234_1385),
	.C2V_20 (C2V_234_1386),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU235 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_44_235),
	.V2C_2 (V2C_80_235),
	.V2C_3 (V2C_100_235),
	.V2C_4 (V2C_161_235),
	.V2C_5 (V2C_223_235),
	.V2C_6 (V2C_266_235),
	.V2C_7 (V2C_366_235),
	.V2C_8 (V2C_420_235),
	.V2C_9 (V2C_517_235),
	.V2C_10 (V2C_753_235),
	.V2C_11 (V2C_801_235),
	.V2C_12 (V2C_849_235),
	.V2C_13 (V2C_890_235),
	.V2C_14 (V2C_931_235),
	.V2C_15 (V2C_965_235),
	.V2C_16 (V2C_1052_235),
	.V2C_17 (V2C_1078_235),
	.V2C_18 (V2C_1137_235),
	.V2C_19 (V2C_1386_235),
	.V2C_20 (V2C_1387_235),
	.C2V_1 (C2V_235_44),
	.C2V_2 (C2V_235_80),
	.C2V_3 (C2V_235_100),
	.C2V_4 (C2V_235_161),
	.C2V_5 (C2V_235_223),
	.C2V_6 (C2V_235_266),
	.C2V_7 (C2V_235_366),
	.C2V_8 (C2V_235_420),
	.C2V_9 (C2V_235_517),
	.C2V_10 (C2V_235_753),
	.C2V_11 (C2V_235_801),
	.C2V_12 (C2V_235_849),
	.C2V_13 (C2V_235_890),
	.C2V_14 (C2V_235_931),
	.C2V_15 (C2V_235_965),
	.C2V_16 (C2V_235_1052),
	.C2V_17 (C2V_235_1078),
	.C2V_18 (C2V_235_1137),
	.C2V_19 (C2V_235_1386),
	.C2V_20 (C2V_235_1387),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU236 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_5_236),
	.V2C_2 (V2C_54_236),
	.V2C_3 (V2C_110_236),
	.V2C_4 (V2C_158_236),
	.V2C_5 (V2C_235_236),
	.V2C_6 (V2C_256_236),
	.V2C_7 (V2C_307_236),
	.V2C_8 (V2C_414_236),
	.V2C_9 (V2C_503_236),
	.V2C_10 (V2C_663_236),
	.V2C_11 (V2C_676_236),
	.V2C_12 (V2C_844_236),
	.V2C_13 (V2C_886_236),
	.V2C_14 (V2C_949_236),
	.V2C_15 (V2C_980_236),
	.V2C_16 (V2C_1012_236),
	.V2C_17 (V2C_1079_236),
	.V2C_18 (V2C_1110_236),
	.V2C_19 (V2C_1387_236),
	.V2C_20 (V2C_1388_236),
	.C2V_1 (C2V_236_5),
	.C2V_2 (C2V_236_54),
	.C2V_3 (C2V_236_110),
	.C2V_4 (C2V_236_158),
	.C2V_5 (C2V_236_235),
	.C2V_6 (C2V_236_256),
	.C2V_7 (C2V_236_307),
	.C2V_8 (C2V_236_414),
	.C2V_9 (C2V_236_503),
	.C2V_10 (C2V_236_663),
	.C2V_11 (C2V_236_676),
	.C2V_12 (C2V_236_844),
	.C2V_13 (C2V_236_886),
	.C2V_14 (C2V_236_949),
	.C2V_15 (C2V_236_980),
	.C2V_16 (C2V_236_1012),
	.C2V_17 (C2V_236_1079),
	.C2V_18 (C2V_236_1110),
	.C2V_19 (C2V_236_1387),
	.C2V_20 (C2V_236_1388),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU237 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_48_237),
	.V2C_2 (V2C_75_237),
	.V2C_3 (V2C_140_237),
	.V2C_4 (V2C_174_237),
	.V2C_5 (V2C_240_237),
	.V2C_6 (V2C_259_237),
	.V2C_7 (V2C_356_237),
	.V2C_8 (V2C_411_237),
	.V2C_9 (V2C_570_237),
	.V2C_10 (V2C_579_237),
	.V2C_11 (V2C_655_237),
	.V2C_12 (V2C_759_237),
	.V2C_13 (V2C_890_237),
	.V2C_14 (V2C_934_237),
	.V2C_15 (V2C_1007_237),
	.V2C_16 (V2C_1019_237),
	.V2C_17 (V2C_1097_237),
	.V2C_18 (V2C_1142_237),
	.V2C_19 (V2C_1388_237),
	.V2C_20 (V2C_1389_237),
	.C2V_1 (C2V_237_48),
	.C2V_2 (C2V_237_75),
	.C2V_3 (C2V_237_140),
	.C2V_4 (C2V_237_174),
	.C2V_5 (C2V_237_240),
	.C2V_6 (C2V_237_259),
	.C2V_7 (C2V_237_356),
	.C2V_8 (C2V_237_411),
	.C2V_9 (C2V_237_570),
	.C2V_10 (C2V_237_579),
	.C2V_11 (C2V_237_655),
	.C2V_12 (C2V_237_759),
	.C2V_13 (C2V_237_890),
	.C2V_14 (C2V_237_934),
	.C2V_15 (C2V_237_1007),
	.C2V_16 (C2V_237_1019),
	.C2V_17 (C2V_237_1097),
	.C2V_18 (C2V_237_1142),
	.C2V_19 (C2V_237_1388),
	.C2V_20 (C2V_237_1389),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU238 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_19_238),
	.V2C_2 (V2C_78_238),
	.V2C_3 (V2C_117_238),
	.V2C_4 (V2C_173_238),
	.V2C_5 (V2C_238_238),
	.V2C_6 (V2C_244_238),
	.V2C_7 (V2C_468_238),
	.V2C_8 (V2C_508_238),
	.V2C_9 (V2C_544_238),
	.V2C_10 (V2C_606_238),
	.V2C_11 (V2C_631_238),
	.V2C_12 (V2C_677_238),
	.V2C_13 (V2C_894_238),
	.V2C_14 (V2C_918_238),
	.V2C_15 (V2C_1002_238),
	.V2C_16 (V2C_1032_238),
	.V2C_17 (V2C_1059_238),
	.V2C_18 (V2C_1123_238),
	.V2C_19 (V2C_1389_238),
	.V2C_20 (V2C_1390_238),
	.C2V_1 (C2V_238_19),
	.C2V_2 (C2V_238_78),
	.C2V_3 (C2V_238_117),
	.C2V_4 (C2V_238_173),
	.C2V_5 (C2V_238_238),
	.C2V_6 (C2V_238_244),
	.C2V_7 (C2V_238_468),
	.C2V_8 (C2V_238_508),
	.C2V_9 (C2V_238_544),
	.C2V_10 (C2V_238_606),
	.C2V_11 (C2V_238_631),
	.C2V_12 (C2V_238_677),
	.C2V_13 (C2V_238_894),
	.C2V_14 (C2V_238_918),
	.C2V_15 (C2V_238_1002),
	.C2V_16 (C2V_238_1032),
	.C2V_17 (C2V_238_1059),
	.C2V_18 (C2V_238_1123),
	.C2V_19 (C2V_238_1389),
	.C2V_20 (C2V_238_1390),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU239 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_38_239),
	.V2C_2 (V2C_96_239),
	.V2C_3 (V2C_131_239),
	.V2C_4 (V2C_154_239),
	.V2C_5 (V2C_218_239),
	.V2C_6 (V2C_284_239),
	.V2C_7 (V2C_333_239),
	.V2C_8 (V2C_352_239),
	.V2C_9 (V2C_479_239),
	.V2C_10 (V2C_713_239),
	.V2C_11 (V2C_729_239),
	.V2C_12 (V2C_783_239),
	.V2C_13 (V2C_909_239),
	.V2C_14 (V2C_957_239),
	.V2C_15 (V2C_1000_239),
	.V2C_16 (V2C_1052_239),
	.V2C_17 (V2C_1101_239),
	.V2C_18 (V2C_1149_239),
	.V2C_19 (V2C_1390_239),
	.V2C_20 (V2C_1391_239),
	.C2V_1 (C2V_239_38),
	.C2V_2 (C2V_239_96),
	.C2V_3 (C2V_239_131),
	.C2V_4 (C2V_239_154),
	.C2V_5 (C2V_239_218),
	.C2V_6 (C2V_239_284),
	.C2V_7 (C2V_239_333),
	.C2V_8 (C2V_239_352),
	.C2V_9 (C2V_239_479),
	.C2V_10 (C2V_239_713),
	.C2V_11 (C2V_239_729),
	.C2V_12 (C2V_239_783),
	.C2V_13 (C2V_239_909),
	.C2V_14 (C2V_239_957),
	.C2V_15 (C2V_239_1000),
	.C2V_16 (C2V_239_1052),
	.C2V_17 (C2V_239_1101),
	.C2V_18 (C2V_239_1149),
	.C2V_19 (C2V_239_1390),
	.C2V_20 (C2V_239_1391),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU240 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_21_240),
	.V2C_2 (V2C_93_240),
	.V2C_3 (V2C_133_240),
	.V2C_4 (V2C_153_240),
	.V2C_5 (V2C_235_240),
	.V2C_6 (V2C_266_240),
	.V2C_7 (V2C_319_240),
	.V2C_8 (V2C_471_240),
	.V2C_9 (V2C_568_240),
	.V2C_10 (V2C_601_240),
	.V2C_11 (V2C_805_240),
	.V2C_12 (V2C_833_240),
	.V2C_13 (V2C_866_240),
	.V2C_14 (V2C_928_240),
	.V2C_15 (V2C_963_240),
	.V2C_16 (V2C_1030_240),
	.V2C_17 (V2C_1094_240),
	.V2C_18 (V2C_1144_240),
	.V2C_19 (V2C_1391_240),
	.V2C_20 (V2C_1392_240),
	.C2V_1 (C2V_240_21),
	.C2V_2 (C2V_240_93),
	.C2V_3 (C2V_240_133),
	.C2V_4 (C2V_240_153),
	.C2V_5 (C2V_240_235),
	.C2V_6 (C2V_240_266),
	.C2V_7 (C2V_240_319),
	.C2V_8 (C2V_240_471),
	.C2V_9 (C2V_240_568),
	.C2V_10 (C2V_240_601),
	.C2V_11 (C2V_240_805),
	.C2V_12 (C2V_240_833),
	.C2V_13 (C2V_240_866),
	.C2V_14 (C2V_240_928),
	.C2V_15 (C2V_240_963),
	.C2V_16 (C2V_240_1030),
	.C2V_17 (C2V_240_1094),
	.C2V_18 (C2V_240_1144),
	.C2V_19 (C2V_240_1391),
	.C2V_20 (C2V_240_1392),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU241 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_45_241),
	.V2C_2 (V2C_81_241),
	.V2C_3 (V2C_101_241),
	.V2C_4 (V2C_162_241),
	.V2C_5 (V2C_224_241),
	.V2C_6 (V2C_267_241),
	.V2C_7 (V2C_367_241),
	.V2C_8 (V2C_421_241),
	.V2C_9 (V2C_518_241),
	.V2C_10 (V2C_754_241),
	.V2C_11 (V2C_802_241),
	.V2C_12 (V2C_850_241),
	.V2C_13 (V2C_891_241),
	.V2C_14 (V2C_932_241),
	.V2C_15 (V2C_966_241),
	.V2C_16 (V2C_1053_241),
	.V2C_17 (V2C_1079_241),
	.V2C_18 (V2C_1138_241),
	.V2C_19 (V2C_1392_241),
	.V2C_20 (V2C_1393_241),
	.C2V_1 (C2V_241_45),
	.C2V_2 (C2V_241_81),
	.C2V_3 (C2V_241_101),
	.C2V_4 (C2V_241_162),
	.C2V_5 (C2V_241_224),
	.C2V_6 (C2V_241_267),
	.C2V_7 (C2V_241_367),
	.C2V_8 (C2V_241_421),
	.C2V_9 (C2V_241_518),
	.C2V_10 (C2V_241_754),
	.C2V_11 (C2V_241_802),
	.C2V_12 (C2V_241_850),
	.C2V_13 (C2V_241_891),
	.C2V_14 (C2V_241_932),
	.C2V_15 (C2V_241_966),
	.C2V_16 (C2V_241_1053),
	.C2V_17 (C2V_241_1079),
	.C2V_18 (C2V_241_1138),
	.C2V_19 (C2V_241_1392),
	.C2V_20 (C2V_241_1393),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU242 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_6_242),
	.V2C_2 (V2C_55_242),
	.V2C_3 (V2C_111_242),
	.V2C_4 (V2C_159_242),
	.V2C_5 (V2C_236_242),
	.V2C_6 (V2C_257_242),
	.V2C_7 (V2C_308_242),
	.V2C_8 (V2C_415_242),
	.V2C_9 (V2C_504_242),
	.V2C_10 (V2C_664_242),
	.V2C_11 (V2C_677_242),
	.V2C_12 (V2C_845_242),
	.V2C_13 (V2C_887_242),
	.V2C_14 (V2C_950_242),
	.V2C_15 (V2C_981_242),
	.V2C_16 (V2C_1013_242),
	.V2C_17 (V2C_1080_242),
	.V2C_18 (V2C_1111_242),
	.V2C_19 (V2C_1393_242),
	.V2C_20 (V2C_1394_242),
	.C2V_1 (C2V_242_6),
	.C2V_2 (C2V_242_55),
	.C2V_3 (C2V_242_111),
	.C2V_4 (C2V_242_159),
	.C2V_5 (C2V_242_236),
	.C2V_6 (C2V_242_257),
	.C2V_7 (C2V_242_308),
	.C2V_8 (C2V_242_415),
	.C2V_9 (C2V_242_504),
	.C2V_10 (C2V_242_664),
	.C2V_11 (C2V_242_677),
	.C2V_12 (C2V_242_845),
	.C2V_13 (C2V_242_887),
	.C2V_14 (C2V_242_950),
	.C2V_15 (C2V_242_981),
	.C2V_16 (C2V_242_1013),
	.C2V_17 (C2V_242_1080),
	.C2V_18 (C2V_242_1111),
	.C2V_19 (C2V_242_1393),
	.C2V_20 (C2V_242_1394),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU243 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_1_243),
	.V2C_2 (V2C_76_243),
	.V2C_3 (V2C_141_243),
	.V2C_4 (V2C_175_243),
	.V2C_5 (V2C_193_243),
	.V2C_6 (V2C_260_243),
	.V2C_7 (V2C_357_243),
	.V2C_8 (V2C_412_243),
	.V2C_9 (V2C_571_243),
	.V2C_10 (V2C_580_243),
	.V2C_11 (V2C_656_243),
	.V2C_12 (V2C_760_243),
	.V2C_13 (V2C_891_243),
	.V2C_14 (V2C_935_243),
	.V2C_15 (V2C_1008_243),
	.V2C_16 (V2C_1020_243),
	.V2C_17 (V2C_1098_243),
	.V2C_18 (V2C_1143_243),
	.V2C_19 (V2C_1394_243),
	.V2C_20 (V2C_1395_243),
	.C2V_1 (C2V_243_1),
	.C2V_2 (C2V_243_76),
	.C2V_3 (C2V_243_141),
	.C2V_4 (C2V_243_175),
	.C2V_5 (C2V_243_193),
	.C2V_6 (C2V_243_260),
	.C2V_7 (C2V_243_357),
	.C2V_8 (C2V_243_412),
	.C2V_9 (C2V_243_571),
	.C2V_10 (C2V_243_580),
	.C2V_11 (C2V_243_656),
	.C2V_12 (C2V_243_760),
	.C2V_13 (C2V_243_891),
	.C2V_14 (C2V_243_935),
	.C2V_15 (C2V_243_1008),
	.C2V_16 (C2V_243_1020),
	.C2V_17 (C2V_243_1098),
	.C2V_18 (C2V_243_1143),
	.C2V_19 (C2V_243_1394),
	.C2V_20 (C2V_243_1395),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU244 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_20_244),
	.V2C_2 (V2C_79_244),
	.V2C_3 (V2C_118_244),
	.V2C_4 (V2C_174_244),
	.V2C_5 (V2C_239_244),
	.V2C_6 (V2C_245_244),
	.V2C_7 (V2C_469_244),
	.V2C_8 (V2C_509_244),
	.V2C_9 (V2C_545_244),
	.V2C_10 (V2C_607_244),
	.V2C_11 (V2C_632_244),
	.V2C_12 (V2C_678_244),
	.V2C_13 (V2C_895_244),
	.V2C_14 (V2C_919_244),
	.V2C_15 (V2C_1003_244),
	.V2C_16 (V2C_1033_244),
	.V2C_17 (V2C_1060_244),
	.V2C_18 (V2C_1124_244),
	.V2C_19 (V2C_1395_244),
	.V2C_20 (V2C_1396_244),
	.C2V_1 (C2V_244_20),
	.C2V_2 (C2V_244_79),
	.C2V_3 (C2V_244_118),
	.C2V_4 (C2V_244_174),
	.C2V_5 (C2V_244_239),
	.C2V_6 (C2V_244_245),
	.C2V_7 (C2V_244_469),
	.C2V_8 (C2V_244_509),
	.C2V_9 (C2V_244_545),
	.C2V_10 (C2V_244_607),
	.C2V_11 (C2V_244_632),
	.C2V_12 (C2V_244_678),
	.C2V_13 (C2V_244_895),
	.C2V_14 (C2V_244_919),
	.C2V_15 (C2V_244_1003),
	.C2V_16 (C2V_244_1033),
	.C2V_17 (C2V_244_1060),
	.C2V_18 (C2V_244_1124),
	.C2V_19 (C2V_244_1395),
	.C2V_20 (C2V_244_1396),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU245 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_39_245),
	.V2C_2 (V2C_49_245),
	.V2C_3 (V2C_132_245),
	.V2C_4 (V2C_155_245),
	.V2C_5 (V2C_219_245),
	.V2C_6 (V2C_285_245),
	.V2C_7 (V2C_334_245),
	.V2C_8 (V2C_353_245),
	.V2C_9 (V2C_480_245),
	.V2C_10 (V2C_714_245),
	.V2C_11 (V2C_730_245),
	.V2C_12 (V2C_784_245),
	.V2C_13 (V2C_910_245),
	.V2C_14 (V2C_958_245),
	.V2C_15 (V2C_1001_245),
	.V2C_16 (V2C_1053_245),
	.V2C_17 (V2C_1102_245),
	.V2C_18 (V2C_1150_245),
	.V2C_19 (V2C_1396_245),
	.V2C_20 (V2C_1397_245),
	.C2V_1 (C2V_245_39),
	.C2V_2 (C2V_245_49),
	.C2V_3 (C2V_245_132),
	.C2V_4 (C2V_245_155),
	.C2V_5 (C2V_245_219),
	.C2V_6 (C2V_245_285),
	.C2V_7 (C2V_245_334),
	.C2V_8 (C2V_245_353),
	.C2V_9 (C2V_245_480),
	.C2V_10 (C2V_245_714),
	.C2V_11 (C2V_245_730),
	.C2V_12 (C2V_245_784),
	.C2V_13 (C2V_245_910),
	.C2V_14 (C2V_245_958),
	.C2V_15 (C2V_245_1001),
	.C2V_16 (C2V_245_1053),
	.C2V_17 (C2V_245_1102),
	.C2V_18 (C2V_245_1150),
	.C2V_19 (C2V_245_1396),
	.C2V_20 (C2V_245_1397),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU246 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_22_246),
	.V2C_2 (V2C_94_246),
	.V2C_3 (V2C_134_246),
	.V2C_4 (V2C_154_246),
	.V2C_5 (V2C_236_246),
	.V2C_6 (V2C_267_246),
	.V2C_7 (V2C_320_246),
	.V2C_8 (V2C_472_246),
	.V2C_9 (V2C_569_246),
	.V2C_10 (V2C_602_246),
	.V2C_11 (V2C_806_246),
	.V2C_12 (V2C_834_246),
	.V2C_13 (V2C_867_246),
	.V2C_14 (V2C_929_246),
	.V2C_15 (V2C_964_246),
	.V2C_16 (V2C_1031_246),
	.V2C_17 (V2C_1095_246),
	.V2C_18 (V2C_1145_246),
	.V2C_19 (V2C_1397_246),
	.V2C_20 (V2C_1398_246),
	.C2V_1 (C2V_246_22),
	.C2V_2 (C2V_246_94),
	.C2V_3 (C2V_246_134),
	.C2V_4 (C2V_246_154),
	.C2V_5 (C2V_246_236),
	.C2V_6 (C2V_246_267),
	.C2V_7 (C2V_246_320),
	.C2V_8 (C2V_246_472),
	.C2V_9 (C2V_246_569),
	.C2V_10 (C2V_246_602),
	.C2V_11 (C2V_246_806),
	.C2V_12 (C2V_246_834),
	.C2V_13 (C2V_246_867),
	.C2V_14 (C2V_246_929),
	.C2V_15 (C2V_246_964),
	.C2V_16 (C2V_246_1031),
	.C2V_17 (C2V_246_1095),
	.C2V_18 (C2V_246_1145),
	.C2V_19 (C2V_246_1397),
	.C2V_20 (C2V_246_1398),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU247 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_46_247),
	.V2C_2 (V2C_82_247),
	.V2C_3 (V2C_102_247),
	.V2C_4 (V2C_163_247),
	.V2C_5 (V2C_225_247),
	.V2C_6 (V2C_268_247),
	.V2C_7 (V2C_368_247),
	.V2C_8 (V2C_422_247),
	.V2C_9 (V2C_519_247),
	.V2C_10 (V2C_755_247),
	.V2C_11 (V2C_803_247),
	.V2C_12 (V2C_851_247),
	.V2C_13 (V2C_892_247),
	.V2C_14 (V2C_933_247),
	.V2C_15 (V2C_967_247),
	.V2C_16 (V2C_1054_247),
	.V2C_17 (V2C_1080_247),
	.V2C_18 (V2C_1139_247),
	.V2C_19 (V2C_1398_247),
	.V2C_20 (V2C_1399_247),
	.C2V_1 (C2V_247_46),
	.C2V_2 (C2V_247_82),
	.C2V_3 (C2V_247_102),
	.C2V_4 (C2V_247_163),
	.C2V_5 (C2V_247_225),
	.C2V_6 (C2V_247_268),
	.C2V_7 (C2V_247_368),
	.C2V_8 (C2V_247_422),
	.C2V_9 (C2V_247_519),
	.C2V_10 (C2V_247_755),
	.C2V_11 (C2V_247_803),
	.C2V_12 (C2V_247_851),
	.C2V_13 (C2V_247_892),
	.C2V_14 (C2V_247_933),
	.C2V_15 (C2V_247_967),
	.C2V_16 (C2V_247_1054),
	.C2V_17 (C2V_247_1080),
	.C2V_18 (C2V_247_1139),
	.C2V_19 (C2V_247_1398),
	.C2V_20 (C2V_247_1399),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU248 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_7_248),
	.V2C_2 (V2C_56_248),
	.V2C_3 (V2C_112_248),
	.V2C_4 (V2C_160_248),
	.V2C_5 (V2C_237_248),
	.V2C_6 (V2C_258_248),
	.V2C_7 (V2C_309_248),
	.V2C_8 (V2C_416_248),
	.V2C_9 (V2C_505_248),
	.V2C_10 (V2C_665_248),
	.V2C_11 (V2C_678_248),
	.V2C_12 (V2C_846_248),
	.V2C_13 (V2C_888_248),
	.V2C_14 (V2C_951_248),
	.V2C_15 (V2C_982_248),
	.V2C_16 (V2C_1014_248),
	.V2C_17 (V2C_1081_248),
	.V2C_18 (V2C_1112_248),
	.V2C_19 (V2C_1399_248),
	.V2C_20 (V2C_1400_248),
	.C2V_1 (C2V_248_7),
	.C2V_2 (C2V_248_56),
	.C2V_3 (C2V_248_112),
	.C2V_4 (C2V_248_160),
	.C2V_5 (C2V_248_237),
	.C2V_6 (C2V_248_258),
	.C2V_7 (C2V_248_309),
	.C2V_8 (C2V_248_416),
	.C2V_9 (C2V_248_505),
	.C2V_10 (C2V_248_665),
	.C2V_11 (C2V_248_678),
	.C2V_12 (C2V_248_846),
	.C2V_13 (C2V_248_888),
	.C2V_14 (C2V_248_951),
	.C2V_15 (C2V_248_982),
	.C2V_16 (C2V_248_1014),
	.C2V_17 (C2V_248_1081),
	.C2V_18 (C2V_248_1112),
	.C2V_19 (C2V_248_1399),
	.C2V_20 (C2V_248_1400),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU249 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_2_249),
	.V2C_2 (V2C_77_249),
	.V2C_3 (V2C_142_249),
	.V2C_4 (V2C_176_249),
	.V2C_5 (V2C_194_249),
	.V2C_6 (V2C_261_249),
	.V2C_7 (V2C_358_249),
	.V2C_8 (V2C_413_249),
	.V2C_9 (V2C_572_249),
	.V2C_10 (V2C_581_249),
	.V2C_11 (V2C_657_249),
	.V2C_12 (V2C_761_249),
	.V2C_13 (V2C_892_249),
	.V2C_14 (V2C_936_249),
	.V2C_15 (V2C_961_249),
	.V2C_16 (V2C_1021_249),
	.V2C_17 (V2C_1099_249),
	.V2C_18 (V2C_1144_249),
	.V2C_19 (V2C_1400_249),
	.V2C_20 (V2C_1401_249),
	.C2V_1 (C2V_249_2),
	.C2V_2 (C2V_249_77),
	.C2V_3 (C2V_249_142),
	.C2V_4 (C2V_249_176),
	.C2V_5 (C2V_249_194),
	.C2V_6 (C2V_249_261),
	.C2V_7 (C2V_249_358),
	.C2V_8 (C2V_249_413),
	.C2V_9 (C2V_249_572),
	.C2V_10 (C2V_249_581),
	.C2V_11 (C2V_249_657),
	.C2V_12 (C2V_249_761),
	.C2V_13 (C2V_249_892),
	.C2V_14 (C2V_249_936),
	.C2V_15 (C2V_249_961),
	.C2V_16 (C2V_249_1021),
	.C2V_17 (C2V_249_1099),
	.C2V_18 (C2V_249_1144),
	.C2V_19 (C2V_249_1400),
	.C2V_20 (C2V_249_1401),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU250 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_21_250),
	.V2C_2 (V2C_80_250),
	.V2C_3 (V2C_119_250),
	.V2C_4 (V2C_175_250),
	.V2C_5 (V2C_240_250),
	.V2C_6 (V2C_246_250),
	.V2C_7 (V2C_470_250),
	.V2C_8 (V2C_510_250),
	.V2C_9 (V2C_546_250),
	.V2C_10 (V2C_608_250),
	.V2C_11 (V2C_633_250),
	.V2C_12 (V2C_679_250),
	.V2C_13 (V2C_896_250),
	.V2C_14 (V2C_920_250),
	.V2C_15 (V2C_1004_250),
	.V2C_16 (V2C_1034_250),
	.V2C_17 (V2C_1061_250),
	.V2C_18 (V2C_1125_250),
	.V2C_19 (V2C_1401_250),
	.V2C_20 (V2C_1402_250),
	.C2V_1 (C2V_250_21),
	.C2V_2 (C2V_250_80),
	.C2V_3 (C2V_250_119),
	.C2V_4 (C2V_250_175),
	.C2V_5 (C2V_250_240),
	.C2V_6 (C2V_250_246),
	.C2V_7 (C2V_250_470),
	.C2V_8 (C2V_250_510),
	.C2V_9 (C2V_250_546),
	.C2V_10 (C2V_250_608),
	.C2V_11 (C2V_250_633),
	.C2V_12 (C2V_250_679),
	.C2V_13 (C2V_250_896),
	.C2V_14 (C2V_250_920),
	.C2V_15 (C2V_250_1004),
	.C2V_16 (C2V_250_1034),
	.C2V_17 (C2V_250_1061),
	.C2V_18 (C2V_250_1125),
	.C2V_19 (C2V_250_1401),
	.C2V_20 (C2V_250_1402),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU251 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_40_251),
	.V2C_2 (V2C_50_251),
	.V2C_3 (V2C_133_251),
	.V2C_4 (V2C_156_251),
	.V2C_5 (V2C_220_251),
	.V2C_6 (V2C_286_251),
	.V2C_7 (V2C_335_251),
	.V2C_8 (V2C_354_251),
	.V2C_9 (V2C_433_251),
	.V2C_10 (V2C_715_251),
	.V2C_11 (V2C_731_251),
	.V2C_12 (V2C_785_251),
	.V2C_13 (V2C_911_251),
	.V2C_14 (V2C_959_251),
	.V2C_15 (V2C_1002_251),
	.V2C_16 (V2C_1054_251),
	.V2C_17 (V2C_1103_251),
	.V2C_18 (V2C_1151_251),
	.V2C_19 (V2C_1402_251),
	.V2C_20 (V2C_1403_251),
	.C2V_1 (C2V_251_40),
	.C2V_2 (C2V_251_50),
	.C2V_3 (C2V_251_133),
	.C2V_4 (C2V_251_156),
	.C2V_5 (C2V_251_220),
	.C2V_6 (C2V_251_286),
	.C2V_7 (C2V_251_335),
	.C2V_8 (C2V_251_354),
	.C2V_9 (C2V_251_433),
	.C2V_10 (C2V_251_715),
	.C2V_11 (C2V_251_731),
	.C2V_12 (C2V_251_785),
	.C2V_13 (C2V_251_911),
	.C2V_14 (C2V_251_959),
	.C2V_15 (C2V_251_1002),
	.C2V_16 (C2V_251_1054),
	.C2V_17 (C2V_251_1103),
	.C2V_18 (C2V_251_1151),
	.C2V_19 (C2V_251_1402),
	.C2V_20 (C2V_251_1403),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU252 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_23_252),
	.V2C_2 (V2C_95_252),
	.V2C_3 (V2C_135_252),
	.V2C_4 (V2C_155_252),
	.V2C_5 (V2C_237_252),
	.V2C_6 (V2C_268_252),
	.V2C_7 (V2C_321_252),
	.V2C_8 (V2C_473_252),
	.V2C_9 (V2C_570_252),
	.V2C_10 (V2C_603_252),
	.V2C_11 (V2C_807_252),
	.V2C_12 (V2C_835_252),
	.V2C_13 (V2C_868_252),
	.V2C_14 (V2C_930_252),
	.V2C_15 (V2C_965_252),
	.V2C_16 (V2C_1032_252),
	.V2C_17 (V2C_1096_252),
	.V2C_18 (V2C_1146_252),
	.V2C_19 (V2C_1403_252),
	.V2C_20 (V2C_1404_252),
	.C2V_1 (C2V_252_23),
	.C2V_2 (C2V_252_95),
	.C2V_3 (C2V_252_135),
	.C2V_4 (C2V_252_155),
	.C2V_5 (C2V_252_237),
	.C2V_6 (C2V_252_268),
	.C2V_7 (C2V_252_321),
	.C2V_8 (C2V_252_473),
	.C2V_9 (C2V_252_570),
	.C2V_10 (C2V_252_603),
	.C2V_11 (C2V_252_807),
	.C2V_12 (C2V_252_835),
	.C2V_13 (C2V_252_868),
	.C2V_14 (C2V_252_930),
	.C2V_15 (C2V_252_965),
	.C2V_16 (C2V_252_1032),
	.C2V_17 (C2V_252_1096),
	.C2V_18 (C2V_252_1146),
	.C2V_19 (C2V_252_1403),
	.C2V_20 (C2V_252_1404),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU253 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_47_253),
	.V2C_2 (V2C_83_253),
	.V2C_3 (V2C_103_253),
	.V2C_4 (V2C_164_253),
	.V2C_5 (V2C_226_253),
	.V2C_6 (V2C_269_253),
	.V2C_7 (V2C_369_253),
	.V2C_8 (V2C_423_253),
	.V2C_9 (V2C_520_253),
	.V2C_10 (V2C_756_253),
	.V2C_11 (V2C_804_253),
	.V2C_12 (V2C_852_253),
	.V2C_13 (V2C_893_253),
	.V2C_14 (V2C_934_253),
	.V2C_15 (V2C_968_253),
	.V2C_16 (V2C_1055_253),
	.V2C_17 (V2C_1081_253),
	.V2C_18 (V2C_1140_253),
	.V2C_19 (V2C_1404_253),
	.V2C_20 (V2C_1405_253),
	.C2V_1 (C2V_253_47),
	.C2V_2 (C2V_253_83),
	.C2V_3 (C2V_253_103),
	.C2V_4 (C2V_253_164),
	.C2V_5 (C2V_253_226),
	.C2V_6 (C2V_253_269),
	.C2V_7 (C2V_253_369),
	.C2V_8 (C2V_253_423),
	.C2V_9 (C2V_253_520),
	.C2V_10 (C2V_253_756),
	.C2V_11 (C2V_253_804),
	.C2V_12 (C2V_253_852),
	.C2V_13 (C2V_253_893),
	.C2V_14 (C2V_253_934),
	.C2V_15 (C2V_253_968),
	.C2V_16 (C2V_253_1055),
	.C2V_17 (C2V_253_1081),
	.C2V_18 (C2V_253_1140),
	.C2V_19 (C2V_253_1404),
	.C2V_20 (C2V_253_1405),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU254 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_8_254),
	.V2C_2 (V2C_57_254),
	.V2C_3 (V2C_113_254),
	.V2C_4 (V2C_161_254),
	.V2C_5 (V2C_238_254),
	.V2C_6 (V2C_259_254),
	.V2C_7 (V2C_310_254),
	.V2C_8 (V2C_417_254),
	.V2C_9 (V2C_506_254),
	.V2C_10 (V2C_666_254),
	.V2C_11 (V2C_679_254),
	.V2C_12 (V2C_847_254),
	.V2C_13 (V2C_889_254),
	.V2C_14 (V2C_952_254),
	.V2C_15 (V2C_983_254),
	.V2C_16 (V2C_1015_254),
	.V2C_17 (V2C_1082_254),
	.V2C_18 (V2C_1113_254),
	.V2C_19 (V2C_1405_254),
	.V2C_20 (V2C_1406_254),
	.C2V_1 (C2V_254_8),
	.C2V_2 (C2V_254_57),
	.C2V_3 (C2V_254_113),
	.C2V_4 (C2V_254_161),
	.C2V_5 (C2V_254_238),
	.C2V_6 (C2V_254_259),
	.C2V_7 (C2V_254_310),
	.C2V_8 (C2V_254_417),
	.C2V_9 (C2V_254_506),
	.C2V_10 (C2V_254_666),
	.C2V_11 (C2V_254_679),
	.C2V_12 (C2V_254_847),
	.C2V_13 (C2V_254_889),
	.C2V_14 (C2V_254_952),
	.C2V_15 (C2V_254_983),
	.C2V_16 (C2V_254_1015),
	.C2V_17 (C2V_254_1082),
	.C2V_18 (C2V_254_1113),
	.C2V_19 (C2V_254_1405),
	.C2V_20 (C2V_254_1406),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU255 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_3_255),
	.V2C_2 (V2C_78_255),
	.V2C_3 (V2C_143_255),
	.V2C_4 (V2C_177_255),
	.V2C_5 (V2C_195_255),
	.V2C_6 (V2C_262_255),
	.V2C_7 (V2C_359_255),
	.V2C_8 (V2C_414_255),
	.V2C_9 (V2C_573_255),
	.V2C_10 (V2C_582_255),
	.V2C_11 (V2C_658_255),
	.V2C_12 (V2C_762_255),
	.V2C_13 (V2C_893_255),
	.V2C_14 (V2C_937_255),
	.V2C_15 (V2C_962_255),
	.V2C_16 (V2C_1022_255),
	.V2C_17 (V2C_1100_255),
	.V2C_18 (V2C_1145_255),
	.V2C_19 (V2C_1406_255),
	.V2C_20 (V2C_1407_255),
	.C2V_1 (C2V_255_3),
	.C2V_2 (C2V_255_78),
	.C2V_3 (C2V_255_143),
	.C2V_4 (C2V_255_177),
	.C2V_5 (C2V_255_195),
	.C2V_6 (C2V_255_262),
	.C2V_7 (C2V_255_359),
	.C2V_8 (C2V_255_414),
	.C2V_9 (C2V_255_573),
	.C2V_10 (C2V_255_582),
	.C2V_11 (C2V_255_658),
	.C2V_12 (C2V_255_762),
	.C2V_13 (C2V_255_893),
	.C2V_14 (C2V_255_937),
	.C2V_15 (C2V_255_962),
	.C2V_16 (C2V_255_1022),
	.C2V_17 (C2V_255_1100),
	.C2V_18 (C2V_255_1145),
	.C2V_19 (C2V_255_1406),
	.C2V_20 (C2V_255_1407),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU256 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_22_256),
	.V2C_2 (V2C_81_256),
	.V2C_3 (V2C_120_256),
	.V2C_4 (V2C_176_256),
	.V2C_5 (V2C_193_256),
	.V2C_6 (V2C_247_256),
	.V2C_7 (V2C_471_256),
	.V2C_8 (V2C_511_256),
	.V2C_9 (V2C_547_256),
	.V2C_10 (V2C_609_256),
	.V2C_11 (V2C_634_256),
	.V2C_12 (V2C_680_256),
	.V2C_13 (V2C_897_256),
	.V2C_14 (V2C_921_256),
	.V2C_15 (V2C_1005_256),
	.V2C_16 (V2C_1035_256),
	.V2C_17 (V2C_1062_256),
	.V2C_18 (V2C_1126_256),
	.V2C_19 (V2C_1407_256),
	.V2C_20 (V2C_1408_256),
	.C2V_1 (C2V_256_22),
	.C2V_2 (C2V_256_81),
	.C2V_3 (C2V_256_120),
	.C2V_4 (C2V_256_176),
	.C2V_5 (C2V_256_193),
	.C2V_6 (C2V_256_247),
	.C2V_7 (C2V_256_471),
	.C2V_8 (C2V_256_511),
	.C2V_9 (C2V_256_547),
	.C2V_10 (C2V_256_609),
	.C2V_11 (C2V_256_634),
	.C2V_12 (C2V_256_680),
	.C2V_13 (C2V_256_897),
	.C2V_14 (C2V_256_921),
	.C2V_15 (C2V_256_1005),
	.C2V_16 (C2V_256_1035),
	.C2V_17 (C2V_256_1062),
	.C2V_18 (C2V_256_1126),
	.C2V_19 (C2V_256_1407),
	.C2V_20 (C2V_256_1408),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU257 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_41_257),
	.V2C_2 (V2C_51_257),
	.V2C_3 (V2C_134_257),
	.V2C_4 (V2C_157_257),
	.V2C_5 (V2C_221_257),
	.V2C_6 (V2C_287_257),
	.V2C_7 (V2C_336_257),
	.V2C_8 (V2C_355_257),
	.V2C_9 (V2C_434_257),
	.V2C_10 (V2C_716_257),
	.V2C_11 (V2C_732_257),
	.V2C_12 (V2C_786_257),
	.V2C_13 (V2C_912_257),
	.V2C_14 (V2C_960_257),
	.V2C_15 (V2C_1003_257),
	.V2C_16 (V2C_1055_257),
	.V2C_17 (V2C_1104_257),
	.V2C_18 (V2C_1152_257),
	.V2C_19 (V2C_1408_257),
	.V2C_20 (V2C_1409_257),
	.C2V_1 (C2V_257_41),
	.C2V_2 (C2V_257_51),
	.C2V_3 (C2V_257_134),
	.C2V_4 (C2V_257_157),
	.C2V_5 (C2V_257_221),
	.C2V_6 (C2V_257_287),
	.C2V_7 (C2V_257_336),
	.C2V_8 (C2V_257_355),
	.C2V_9 (C2V_257_434),
	.C2V_10 (C2V_257_716),
	.C2V_11 (C2V_257_732),
	.C2V_12 (C2V_257_786),
	.C2V_13 (C2V_257_912),
	.C2V_14 (C2V_257_960),
	.C2V_15 (C2V_257_1003),
	.C2V_16 (C2V_257_1055),
	.C2V_17 (C2V_257_1104),
	.C2V_18 (C2V_257_1152),
	.C2V_19 (C2V_257_1408),
	.C2V_20 (C2V_257_1409),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU258 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_24_258),
	.V2C_2 (V2C_96_258),
	.V2C_3 (V2C_136_258),
	.V2C_4 (V2C_156_258),
	.V2C_5 (V2C_238_258),
	.V2C_6 (V2C_269_258),
	.V2C_7 (V2C_322_258),
	.V2C_8 (V2C_474_258),
	.V2C_9 (V2C_571_258),
	.V2C_10 (V2C_604_258),
	.V2C_11 (V2C_808_258),
	.V2C_12 (V2C_836_258),
	.V2C_13 (V2C_869_258),
	.V2C_14 (V2C_931_258),
	.V2C_15 (V2C_966_258),
	.V2C_16 (V2C_1033_258),
	.V2C_17 (V2C_1097_258),
	.V2C_18 (V2C_1147_258),
	.V2C_19 (V2C_1409_258),
	.V2C_20 (V2C_1410_258),
	.C2V_1 (C2V_258_24),
	.C2V_2 (C2V_258_96),
	.C2V_3 (C2V_258_136),
	.C2V_4 (C2V_258_156),
	.C2V_5 (C2V_258_238),
	.C2V_6 (C2V_258_269),
	.C2V_7 (C2V_258_322),
	.C2V_8 (C2V_258_474),
	.C2V_9 (C2V_258_571),
	.C2V_10 (C2V_258_604),
	.C2V_11 (C2V_258_808),
	.C2V_12 (C2V_258_836),
	.C2V_13 (C2V_258_869),
	.C2V_14 (C2V_258_931),
	.C2V_15 (C2V_258_966),
	.C2V_16 (C2V_258_1033),
	.C2V_17 (C2V_258_1097),
	.C2V_18 (C2V_258_1147),
	.C2V_19 (C2V_258_1409),
	.C2V_20 (C2V_258_1410),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU259 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_48_259),
	.V2C_2 (V2C_84_259),
	.V2C_3 (V2C_104_259),
	.V2C_4 (V2C_165_259),
	.V2C_5 (V2C_227_259),
	.V2C_6 (V2C_270_259),
	.V2C_7 (V2C_370_259),
	.V2C_8 (V2C_424_259),
	.V2C_9 (V2C_521_259),
	.V2C_10 (V2C_757_259),
	.V2C_11 (V2C_805_259),
	.V2C_12 (V2C_853_259),
	.V2C_13 (V2C_894_259),
	.V2C_14 (V2C_935_259),
	.V2C_15 (V2C_969_259),
	.V2C_16 (V2C_1056_259),
	.V2C_17 (V2C_1082_259),
	.V2C_18 (V2C_1141_259),
	.V2C_19 (V2C_1410_259),
	.V2C_20 (V2C_1411_259),
	.C2V_1 (C2V_259_48),
	.C2V_2 (C2V_259_84),
	.C2V_3 (C2V_259_104),
	.C2V_4 (C2V_259_165),
	.C2V_5 (C2V_259_227),
	.C2V_6 (C2V_259_270),
	.C2V_7 (C2V_259_370),
	.C2V_8 (C2V_259_424),
	.C2V_9 (C2V_259_521),
	.C2V_10 (C2V_259_757),
	.C2V_11 (C2V_259_805),
	.C2V_12 (C2V_259_853),
	.C2V_13 (C2V_259_894),
	.C2V_14 (C2V_259_935),
	.C2V_15 (C2V_259_969),
	.C2V_16 (C2V_259_1056),
	.C2V_17 (C2V_259_1082),
	.C2V_18 (C2V_259_1141),
	.C2V_19 (C2V_259_1410),
	.C2V_20 (C2V_259_1411),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU260 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_9_260),
	.V2C_2 (V2C_58_260),
	.V2C_3 (V2C_114_260),
	.V2C_4 (V2C_162_260),
	.V2C_5 (V2C_239_260),
	.V2C_6 (V2C_260_260),
	.V2C_7 (V2C_311_260),
	.V2C_8 (V2C_418_260),
	.V2C_9 (V2C_507_260),
	.V2C_10 (V2C_667_260),
	.V2C_11 (V2C_680_260),
	.V2C_12 (V2C_848_260),
	.V2C_13 (V2C_890_260),
	.V2C_14 (V2C_953_260),
	.V2C_15 (V2C_984_260),
	.V2C_16 (V2C_1016_260),
	.V2C_17 (V2C_1083_260),
	.V2C_18 (V2C_1114_260),
	.V2C_19 (V2C_1411_260),
	.V2C_20 (V2C_1412_260),
	.C2V_1 (C2V_260_9),
	.C2V_2 (C2V_260_58),
	.C2V_3 (C2V_260_114),
	.C2V_4 (C2V_260_162),
	.C2V_5 (C2V_260_239),
	.C2V_6 (C2V_260_260),
	.C2V_7 (C2V_260_311),
	.C2V_8 (C2V_260_418),
	.C2V_9 (C2V_260_507),
	.C2V_10 (C2V_260_667),
	.C2V_11 (C2V_260_680),
	.C2V_12 (C2V_260_848),
	.C2V_13 (C2V_260_890),
	.C2V_14 (C2V_260_953),
	.C2V_15 (C2V_260_984),
	.C2V_16 (C2V_260_1016),
	.C2V_17 (C2V_260_1083),
	.C2V_18 (C2V_260_1114),
	.C2V_19 (C2V_260_1411),
	.C2V_20 (C2V_260_1412),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU261 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_4_261),
	.V2C_2 (V2C_79_261),
	.V2C_3 (V2C_144_261),
	.V2C_4 (V2C_178_261),
	.V2C_5 (V2C_196_261),
	.V2C_6 (V2C_263_261),
	.V2C_7 (V2C_360_261),
	.V2C_8 (V2C_415_261),
	.V2C_9 (V2C_574_261),
	.V2C_10 (V2C_583_261),
	.V2C_11 (V2C_659_261),
	.V2C_12 (V2C_763_261),
	.V2C_13 (V2C_894_261),
	.V2C_14 (V2C_938_261),
	.V2C_15 (V2C_963_261),
	.V2C_16 (V2C_1023_261),
	.V2C_17 (V2C_1101_261),
	.V2C_18 (V2C_1146_261),
	.V2C_19 (V2C_1412_261),
	.V2C_20 (V2C_1413_261),
	.C2V_1 (C2V_261_4),
	.C2V_2 (C2V_261_79),
	.C2V_3 (C2V_261_144),
	.C2V_4 (C2V_261_178),
	.C2V_5 (C2V_261_196),
	.C2V_6 (C2V_261_263),
	.C2V_7 (C2V_261_360),
	.C2V_8 (C2V_261_415),
	.C2V_9 (C2V_261_574),
	.C2V_10 (C2V_261_583),
	.C2V_11 (C2V_261_659),
	.C2V_12 (C2V_261_763),
	.C2V_13 (C2V_261_894),
	.C2V_14 (C2V_261_938),
	.C2V_15 (C2V_261_963),
	.C2V_16 (C2V_261_1023),
	.C2V_17 (C2V_261_1101),
	.C2V_18 (C2V_261_1146),
	.C2V_19 (C2V_261_1412),
	.C2V_20 (C2V_261_1413),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU262 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_23_262),
	.V2C_2 (V2C_82_262),
	.V2C_3 (V2C_121_262),
	.V2C_4 (V2C_177_262),
	.V2C_5 (V2C_194_262),
	.V2C_6 (V2C_248_262),
	.V2C_7 (V2C_472_262),
	.V2C_8 (V2C_512_262),
	.V2C_9 (V2C_548_262),
	.V2C_10 (V2C_610_262),
	.V2C_11 (V2C_635_262),
	.V2C_12 (V2C_681_262),
	.V2C_13 (V2C_898_262),
	.V2C_14 (V2C_922_262),
	.V2C_15 (V2C_1006_262),
	.V2C_16 (V2C_1036_262),
	.V2C_17 (V2C_1063_262),
	.V2C_18 (V2C_1127_262),
	.V2C_19 (V2C_1413_262),
	.V2C_20 (V2C_1414_262),
	.C2V_1 (C2V_262_23),
	.C2V_2 (C2V_262_82),
	.C2V_3 (C2V_262_121),
	.C2V_4 (C2V_262_177),
	.C2V_5 (C2V_262_194),
	.C2V_6 (C2V_262_248),
	.C2V_7 (C2V_262_472),
	.C2V_8 (C2V_262_512),
	.C2V_9 (C2V_262_548),
	.C2V_10 (C2V_262_610),
	.C2V_11 (C2V_262_635),
	.C2V_12 (C2V_262_681),
	.C2V_13 (C2V_262_898),
	.C2V_14 (C2V_262_922),
	.C2V_15 (C2V_262_1006),
	.C2V_16 (C2V_262_1036),
	.C2V_17 (C2V_262_1063),
	.C2V_18 (C2V_262_1127),
	.C2V_19 (C2V_262_1413),
	.C2V_20 (C2V_262_1414),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU263 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_42_263),
	.V2C_2 (V2C_52_263),
	.V2C_3 (V2C_135_263),
	.V2C_4 (V2C_158_263),
	.V2C_5 (V2C_222_263),
	.V2C_6 (V2C_288_263),
	.V2C_7 (V2C_289_263),
	.V2C_8 (V2C_356_263),
	.V2C_9 (V2C_435_263),
	.V2C_10 (V2C_717_263),
	.V2C_11 (V2C_733_263),
	.V2C_12 (V2C_787_263),
	.V2C_13 (V2C_865_263),
	.V2C_14 (V2C_913_263),
	.V2C_15 (V2C_1004_263),
	.V2C_16 (V2C_1056_263),
	.V2C_17 (V2C_1057_263),
	.V2C_18 (V2C_1105_263),
	.V2C_19 (V2C_1414_263),
	.V2C_20 (V2C_1415_263),
	.C2V_1 (C2V_263_42),
	.C2V_2 (C2V_263_52),
	.C2V_3 (C2V_263_135),
	.C2V_4 (C2V_263_158),
	.C2V_5 (C2V_263_222),
	.C2V_6 (C2V_263_288),
	.C2V_7 (C2V_263_289),
	.C2V_8 (C2V_263_356),
	.C2V_9 (C2V_263_435),
	.C2V_10 (C2V_263_717),
	.C2V_11 (C2V_263_733),
	.C2V_12 (C2V_263_787),
	.C2V_13 (C2V_263_865),
	.C2V_14 (C2V_263_913),
	.C2V_15 (C2V_263_1004),
	.C2V_16 (C2V_263_1056),
	.C2V_17 (C2V_263_1057),
	.C2V_18 (C2V_263_1105),
	.C2V_19 (C2V_263_1414),
	.C2V_20 (C2V_263_1415),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU264 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_25_264),
	.V2C_2 (V2C_49_264),
	.V2C_3 (V2C_137_264),
	.V2C_4 (V2C_157_264),
	.V2C_5 (V2C_239_264),
	.V2C_6 (V2C_270_264),
	.V2C_7 (V2C_323_264),
	.V2C_8 (V2C_475_264),
	.V2C_9 (V2C_572_264),
	.V2C_10 (V2C_605_264),
	.V2C_11 (V2C_809_264),
	.V2C_12 (V2C_837_264),
	.V2C_13 (V2C_870_264),
	.V2C_14 (V2C_932_264),
	.V2C_15 (V2C_967_264),
	.V2C_16 (V2C_1034_264),
	.V2C_17 (V2C_1098_264),
	.V2C_18 (V2C_1148_264),
	.V2C_19 (V2C_1415_264),
	.V2C_20 (V2C_1416_264),
	.C2V_1 (C2V_264_25),
	.C2V_2 (C2V_264_49),
	.C2V_3 (C2V_264_137),
	.C2V_4 (C2V_264_157),
	.C2V_5 (C2V_264_239),
	.C2V_6 (C2V_264_270),
	.C2V_7 (C2V_264_323),
	.C2V_8 (C2V_264_475),
	.C2V_9 (C2V_264_572),
	.C2V_10 (C2V_264_605),
	.C2V_11 (C2V_264_809),
	.C2V_12 (C2V_264_837),
	.C2V_13 (C2V_264_870),
	.C2V_14 (C2V_264_932),
	.C2V_15 (C2V_264_967),
	.C2V_16 (C2V_264_1034),
	.C2V_17 (C2V_264_1098),
	.C2V_18 (C2V_264_1148),
	.C2V_19 (C2V_264_1415),
	.C2V_20 (C2V_264_1416),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU265 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_1_265),
	.V2C_2 (V2C_85_265),
	.V2C_3 (V2C_105_265),
	.V2C_4 (V2C_166_265),
	.V2C_5 (V2C_228_265),
	.V2C_6 (V2C_271_265),
	.V2C_7 (V2C_371_265),
	.V2C_8 (V2C_425_265),
	.V2C_9 (V2C_522_265),
	.V2C_10 (V2C_758_265),
	.V2C_11 (V2C_806_265),
	.V2C_12 (V2C_854_265),
	.V2C_13 (V2C_895_265),
	.V2C_14 (V2C_936_265),
	.V2C_15 (V2C_970_265),
	.V2C_16 (V2C_1009_265),
	.V2C_17 (V2C_1083_265),
	.V2C_18 (V2C_1142_265),
	.V2C_19 (V2C_1416_265),
	.V2C_20 (V2C_1417_265),
	.C2V_1 (C2V_265_1),
	.C2V_2 (C2V_265_85),
	.C2V_3 (C2V_265_105),
	.C2V_4 (C2V_265_166),
	.C2V_5 (C2V_265_228),
	.C2V_6 (C2V_265_271),
	.C2V_7 (C2V_265_371),
	.C2V_8 (C2V_265_425),
	.C2V_9 (C2V_265_522),
	.C2V_10 (C2V_265_758),
	.C2V_11 (C2V_265_806),
	.C2V_12 (C2V_265_854),
	.C2V_13 (C2V_265_895),
	.C2V_14 (C2V_265_936),
	.C2V_15 (C2V_265_970),
	.C2V_16 (C2V_265_1009),
	.C2V_17 (C2V_265_1083),
	.C2V_18 (C2V_265_1142),
	.C2V_19 (C2V_265_1416),
	.C2V_20 (C2V_265_1417),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU266 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_10_266),
	.V2C_2 (V2C_59_266),
	.V2C_3 (V2C_115_266),
	.V2C_4 (V2C_163_266),
	.V2C_5 (V2C_240_266),
	.V2C_6 (V2C_261_266),
	.V2C_7 (V2C_312_266),
	.V2C_8 (V2C_419_266),
	.V2C_9 (V2C_508_266),
	.V2C_10 (V2C_668_266),
	.V2C_11 (V2C_681_266),
	.V2C_12 (V2C_849_266),
	.V2C_13 (V2C_891_266),
	.V2C_14 (V2C_954_266),
	.V2C_15 (V2C_985_266),
	.V2C_16 (V2C_1017_266),
	.V2C_17 (V2C_1084_266),
	.V2C_18 (V2C_1115_266),
	.V2C_19 (V2C_1417_266),
	.V2C_20 (V2C_1418_266),
	.C2V_1 (C2V_266_10),
	.C2V_2 (C2V_266_59),
	.C2V_3 (C2V_266_115),
	.C2V_4 (C2V_266_163),
	.C2V_5 (C2V_266_240),
	.C2V_6 (C2V_266_261),
	.C2V_7 (C2V_266_312),
	.C2V_8 (C2V_266_419),
	.C2V_9 (C2V_266_508),
	.C2V_10 (C2V_266_668),
	.C2V_11 (C2V_266_681),
	.C2V_12 (C2V_266_849),
	.C2V_13 (C2V_266_891),
	.C2V_14 (C2V_266_954),
	.C2V_15 (C2V_266_985),
	.C2V_16 (C2V_266_1017),
	.C2V_17 (C2V_266_1084),
	.C2V_18 (C2V_266_1115),
	.C2V_19 (C2V_266_1417),
	.C2V_20 (C2V_266_1418),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU267 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_5_267),
	.V2C_2 (V2C_80_267),
	.V2C_3 (V2C_97_267),
	.V2C_4 (V2C_179_267),
	.V2C_5 (V2C_197_267),
	.V2C_6 (V2C_264_267),
	.V2C_7 (V2C_361_267),
	.V2C_8 (V2C_416_267),
	.V2C_9 (V2C_575_267),
	.V2C_10 (V2C_584_267),
	.V2C_11 (V2C_660_267),
	.V2C_12 (V2C_764_267),
	.V2C_13 (V2C_895_267),
	.V2C_14 (V2C_939_267),
	.V2C_15 (V2C_964_267),
	.V2C_16 (V2C_1024_267),
	.V2C_17 (V2C_1102_267),
	.V2C_18 (V2C_1147_267),
	.V2C_19 (V2C_1418_267),
	.V2C_20 (V2C_1419_267),
	.C2V_1 (C2V_267_5),
	.C2V_2 (C2V_267_80),
	.C2V_3 (C2V_267_97),
	.C2V_4 (C2V_267_179),
	.C2V_5 (C2V_267_197),
	.C2V_6 (C2V_267_264),
	.C2V_7 (C2V_267_361),
	.C2V_8 (C2V_267_416),
	.C2V_9 (C2V_267_575),
	.C2V_10 (C2V_267_584),
	.C2V_11 (C2V_267_660),
	.C2V_12 (C2V_267_764),
	.C2V_13 (C2V_267_895),
	.C2V_14 (C2V_267_939),
	.C2V_15 (C2V_267_964),
	.C2V_16 (C2V_267_1024),
	.C2V_17 (C2V_267_1102),
	.C2V_18 (C2V_267_1147),
	.C2V_19 (C2V_267_1418),
	.C2V_20 (C2V_267_1419),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU268 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_24_268),
	.V2C_2 (V2C_83_268),
	.V2C_3 (V2C_122_268),
	.V2C_4 (V2C_178_268),
	.V2C_5 (V2C_195_268),
	.V2C_6 (V2C_249_268),
	.V2C_7 (V2C_473_268),
	.V2C_8 (V2C_513_268),
	.V2C_9 (V2C_549_268),
	.V2C_10 (V2C_611_268),
	.V2C_11 (V2C_636_268),
	.V2C_12 (V2C_682_268),
	.V2C_13 (V2C_899_268),
	.V2C_14 (V2C_923_268),
	.V2C_15 (V2C_1007_268),
	.V2C_16 (V2C_1037_268),
	.V2C_17 (V2C_1064_268),
	.V2C_18 (V2C_1128_268),
	.V2C_19 (V2C_1419_268),
	.V2C_20 (V2C_1420_268),
	.C2V_1 (C2V_268_24),
	.C2V_2 (C2V_268_83),
	.C2V_3 (C2V_268_122),
	.C2V_4 (C2V_268_178),
	.C2V_5 (C2V_268_195),
	.C2V_6 (C2V_268_249),
	.C2V_7 (C2V_268_473),
	.C2V_8 (C2V_268_513),
	.C2V_9 (C2V_268_549),
	.C2V_10 (C2V_268_611),
	.C2V_11 (C2V_268_636),
	.C2V_12 (C2V_268_682),
	.C2V_13 (C2V_268_899),
	.C2V_14 (C2V_268_923),
	.C2V_15 (C2V_268_1007),
	.C2V_16 (C2V_268_1037),
	.C2V_17 (C2V_268_1064),
	.C2V_18 (C2V_268_1128),
	.C2V_19 (C2V_268_1419),
	.C2V_20 (C2V_268_1420),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU269 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_43_269),
	.V2C_2 (V2C_53_269),
	.V2C_3 (V2C_136_269),
	.V2C_4 (V2C_159_269),
	.V2C_5 (V2C_223_269),
	.V2C_6 (V2C_241_269),
	.V2C_7 (V2C_290_269),
	.V2C_8 (V2C_357_269),
	.V2C_9 (V2C_436_269),
	.V2C_10 (V2C_718_269),
	.V2C_11 (V2C_734_269),
	.V2C_12 (V2C_788_269),
	.V2C_13 (V2C_866_269),
	.V2C_14 (V2C_914_269),
	.V2C_15 (V2C_1005_269),
	.V2C_16 (V2C_1009_269),
	.V2C_17 (V2C_1058_269),
	.V2C_18 (V2C_1106_269),
	.V2C_19 (V2C_1420_269),
	.V2C_20 (V2C_1421_269),
	.C2V_1 (C2V_269_43),
	.C2V_2 (C2V_269_53),
	.C2V_3 (C2V_269_136),
	.C2V_4 (C2V_269_159),
	.C2V_5 (C2V_269_223),
	.C2V_6 (C2V_269_241),
	.C2V_7 (C2V_269_290),
	.C2V_8 (C2V_269_357),
	.C2V_9 (C2V_269_436),
	.C2V_10 (C2V_269_718),
	.C2V_11 (C2V_269_734),
	.C2V_12 (C2V_269_788),
	.C2V_13 (C2V_269_866),
	.C2V_14 (C2V_269_914),
	.C2V_15 (C2V_269_1005),
	.C2V_16 (C2V_269_1009),
	.C2V_17 (C2V_269_1058),
	.C2V_18 (C2V_269_1106),
	.C2V_19 (C2V_269_1420),
	.C2V_20 (C2V_269_1421),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU270 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_26_270),
	.V2C_2 (V2C_50_270),
	.V2C_3 (V2C_138_270),
	.V2C_4 (V2C_158_270),
	.V2C_5 (V2C_240_270),
	.V2C_6 (V2C_271_270),
	.V2C_7 (V2C_324_270),
	.V2C_8 (V2C_476_270),
	.V2C_9 (V2C_573_270),
	.V2C_10 (V2C_606_270),
	.V2C_11 (V2C_810_270),
	.V2C_12 (V2C_838_270),
	.V2C_13 (V2C_871_270),
	.V2C_14 (V2C_933_270),
	.V2C_15 (V2C_968_270),
	.V2C_16 (V2C_1035_270),
	.V2C_17 (V2C_1099_270),
	.V2C_18 (V2C_1149_270),
	.V2C_19 (V2C_1421_270),
	.V2C_20 (V2C_1422_270),
	.C2V_1 (C2V_270_26),
	.C2V_2 (C2V_270_50),
	.C2V_3 (C2V_270_138),
	.C2V_4 (C2V_270_158),
	.C2V_5 (C2V_270_240),
	.C2V_6 (C2V_270_271),
	.C2V_7 (C2V_270_324),
	.C2V_8 (C2V_270_476),
	.C2V_9 (C2V_270_573),
	.C2V_10 (C2V_270_606),
	.C2V_11 (C2V_270_810),
	.C2V_12 (C2V_270_838),
	.C2V_13 (C2V_270_871),
	.C2V_14 (C2V_270_933),
	.C2V_15 (C2V_270_968),
	.C2V_16 (C2V_270_1035),
	.C2V_17 (C2V_270_1099),
	.C2V_18 (C2V_270_1149),
	.C2V_19 (C2V_270_1421),
	.C2V_20 (C2V_270_1422),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU271 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_2_271),
	.V2C_2 (V2C_86_271),
	.V2C_3 (V2C_106_271),
	.V2C_4 (V2C_167_271),
	.V2C_5 (V2C_229_271),
	.V2C_6 (V2C_272_271),
	.V2C_7 (V2C_372_271),
	.V2C_8 (V2C_426_271),
	.V2C_9 (V2C_523_271),
	.V2C_10 (V2C_759_271),
	.V2C_11 (V2C_807_271),
	.V2C_12 (V2C_855_271),
	.V2C_13 (V2C_896_271),
	.V2C_14 (V2C_937_271),
	.V2C_15 (V2C_971_271),
	.V2C_16 (V2C_1010_271),
	.V2C_17 (V2C_1084_271),
	.V2C_18 (V2C_1143_271),
	.V2C_19 (V2C_1422_271),
	.V2C_20 (V2C_1423_271),
	.C2V_1 (C2V_271_2),
	.C2V_2 (C2V_271_86),
	.C2V_3 (C2V_271_106),
	.C2V_4 (C2V_271_167),
	.C2V_5 (C2V_271_229),
	.C2V_6 (C2V_271_272),
	.C2V_7 (C2V_271_372),
	.C2V_8 (C2V_271_426),
	.C2V_9 (C2V_271_523),
	.C2V_10 (C2V_271_759),
	.C2V_11 (C2V_271_807),
	.C2V_12 (C2V_271_855),
	.C2V_13 (C2V_271_896),
	.C2V_14 (C2V_271_937),
	.C2V_15 (C2V_271_971),
	.C2V_16 (C2V_271_1010),
	.C2V_17 (C2V_271_1084),
	.C2V_18 (C2V_271_1143),
	.C2V_19 (C2V_271_1422),
	.C2V_20 (C2V_271_1423),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU272 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_11_272),
	.V2C_2 (V2C_60_272),
	.V2C_3 (V2C_116_272),
	.V2C_4 (V2C_164_272),
	.V2C_5 (V2C_193_272),
	.V2C_6 (V2C_262_272),
	.V2C_7 (V2C_313_272),
	.V2C_8 (V2C_420_272),
	.V2C_9 (V2C_509_272),
	.V2C_10 (V2C_669_272),
	.V2C_11 (V2C_682_272),
	.V2C_12 (V2C_850_272),
	.V2C_13 (V2C_892_272),
	.V2C_14 (V2C_955_272),
	.V2C_15 (V2C_986_272),
	.V2C_16 (V2C_1018_272),
	.V2C_17 (V2C_1085_272),
	.V2C_18 (V2C_1116_272),
	.V2C_19 (V2C_1423_272),
	.V2C_20 (V2C_1424_272),
	.C2V_1 (C2V_272_11),
	.C2V_2 (C2V_272_60),
	.C2V_3 (C2V_272_116),
	.C2V_4 (C2V_272_164),
	.C2V_5 (C2V_272_193),
	.C2V_6 (C2V_272_262),
	.C2V_7 (C2V_272_313),
	.C2V_8 (C2V_272_420),
	.C2V_9 (C2V_272_509),
	.C2V_10 (C2V_272_669),
	.C2V_11 (C2V_272_682),
	.C2V_12 (C2V_272_850),
	.C2V_13 (C2V_272_892),
	.C2V_14 (C2V_272_955),
	.C2V_15 (C2V_272_986),
	.C2V_16 (C2V_272_1018),
	.C2V_17 (C2V_272_1085),
	.C2V_18 (C2V_272_1116),
	.C2V_19 (C2V_272_1423),
	.C2V_20 (C2V_272_1424),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU273 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_6_273),
	.V2C_2 (V2C_81_273),
	.V2C_3 (V2C_98_273),
	.V2C_4 (V2C_180_273),
	.V2C_5 (V2C_198_273),
	.V2C_6 (V2C_265_273),
	.V2C_7 (V2C_362_273),
	.V2C_8 (V2C_417_273),
	.V2C_9 (V2C_576_273),
	.V2C_10 (V2C_585_273),
	.V2C_11 (V2C_661_273),
	.V2C_12 (V2C_765_273),
	.V2C_13 (V2C_896_273),
	.V2C_14 (V2C_940_273),
	.V2C_15 (V2C_965_273),
	.V2C_16 (V2C_1025_273),
	.V2C_17 (V2C_1103_273),
	.V2C_18 (V2C_1148_273),
	.V2C_19 (V2C_1424_273),
	.V2C_20 (V2C_1425_273),
	.C2V_1 (C2V_273_6),
	.C2V_2 (C2V_273_81),
	.C2V_3 (C2V_273_98),
	.C2V_4 (C2V_273_180),
	.C2V_5 (C2V_273_198),
	.C2V_6 (C2V_273_265),
	.C2V_7 (C2V_273_362),
	.C2V_8 (C2V_273_417),
	.C2V_9 (C2V_273_576),
	.C2V_10 (C2V_273_585),
	.C2V_11 (C2V_273_661),
	.C2V_12 (C2V_273_765),
	.C2V_13 (C2V_273_896),
	.C2V_14 (C2V_273_940),
	.C2V_15 (C2V_273_965),
	.C2V_16 (C2V_273_1025),
	.C2V_17 (C2V_273_1103),
	.C2V_18 (C2V_273_1148),
	.C2V_19 (C2V_273_1424),
	.C2V_20 (C2V_273_1425),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU274 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_25_274),
	.V2C_2 (V2C_84_274),
	.V2C_3 (V2C_123_274),
	.V2C_4 (V2C_179_274),
	.V2C_5 (V2C_196_274),
	.V2C_6 (V2C_250_274),
	.V2C_7 (V2C_474_274),
	.V2C_8 (V2C_514_274),
	.V2C_9 (V2C_550_274),
	.V2C_10 (V2C_612_274),
	.V2C_11 (V2C_637_274),
	.V2C_12 (V2C_683_274),
	.V2C_13 (V2C_900_274),
	.V2C_14 (V2C_924_274),
	.V2C_15 (V2C_1008_274),
	.V2C_16 (V2C_1038_274),
	.V2C_17 (V2C_1065_274),
	.V2C_18 (V2C_1129_274),
	.V2C_19 (V2C_1425_274),
	.V2C_20 (V2C_1426_274),
	.C2V_1 (C2V_274_25),
	.C2V_2 (C2V_274_84),
	.C2V_3 (C2V_274_123),
	.C2V_4 (C2V_274_179),
	.C2V_5 (C2V_274_196),
	.C2V_6 (C2V_274_250),
	.C2V_7 (C2V_274_474),
	.C2V_8 (C2V_274_514),
	.C2V_9 (C2V_274_550),
	.C2V_10 (C2V_274_612),
	.C2V_11 (C2V_274_637),
	.C2V_12 (C2V_274_683),
	.C2V_13 (C2V_274_900),
	.C2V_14 (C2V_274_924),
	.C2V_15 (C2V_274_1008),
	.C2V_16 (C2V_274_1038),
	.C2V_17 (C2V_274_1065),
	.C2V_18 (C2V_274_1129),
	.C2V_19 (C2V_274_1425),
	.C2V_20 (C2V_274_1426),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU275 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_44_275),
	.V2C_2 (V2C_54_275),
	.V2C_3 (V2C_137_275),
	.V2C_4 (V2C_160_275),
	.V2C_5 (V2C_224_275),
	.V2C_6 (V2C_242_275),
	.V2C_7 (V2C_291_275),
	.V2C_8 (V2C_358_275),
	.V2C_9 (V2C_437_275),
	.V2C_10 (V2C_719_275),
	.V2C_11 (V2C_735_275),
	.V2C_12 (V2C_789_275),
	.V2C_13 (V2C_867_275),
	.V2C_14 (V2C_915_275),
	.V2C_15 (V2C_1006_275),
	.V2C_16 (V2C_1010_275),
	.V2C_17 (V2C_1059_275),
	.V2C_18 (V2C_1107_275),
	.V2C_19 (V2C_1426_275),
	.V2C_20 (V2C_1427_275),
	.C2V_1 (C2V_275_44),
	.C2V_2 (C2V_275_54),
	.C2V_3 (C2V_275_137),
	.C2V_4 (C2V_275_160),
	.C2V_5 (C2V_275_224),
	.C2V_6 (C2V_275_242),
	.C2V_7 (C2V_275_291),
	.C2V_8 (C2V_275_358),
	.C2V_9 (C2V_275_437),
	.C2V_10 (C2V_275_719),
	.C2V_11 (C2V_275_735),
	.C2V_12 (C2V_275_789),
	.C2V_13 (C2V_275_867),
	.C2V_14 (C2V_275_915),
	.C2V_15 (C2V_275_1006),
	.C2V_16 (C2V_275_1010),
	.C2V_17 (C2V_275_1059),
	.C2V_18 (C2V_275_1107),
	.C2V_19 (C2V_275_1426),
	.C2V_20 (C2V_275_1427),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU276 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_27_276),
	.V2C_2 (V2C_51_276),
	.V2C_3 (V2C_139_276),
	.V2C_4 (V2C_159_276),
	.V2C_5 (V2C_193_276),
	.V2C_6 (V2C_272_276),
	.V2C_7 (V2C_325_276),
	.V2C_8 (V2C_477_276),
	.V2C_9 (V2C_574_276),
	.V2C_10 (V2C_607_276),
	.V2C_11 (V2C_811_276),
	.V2C_12 (V2C_839_276),
	.V2C_13 (V2C_872_276),
	.V2C_14 (V2C_934_276),
	.V2C_15 (V2C_969_276),
	.V2C_16 (V2C_1036_276),
	.V2C_17 (V2C_1100_276),
	.V2C_18 (V2C_1150_276),
	.V2C_19 (V2C_1427_276),
	.V2C_20 (V2C_1428_276),
	.C2V_1 (C2V_276_27),
	.C2V_2 (C2V_276_51),
	.C2V_3 (C2V_276_139),
	.C2V_4 (C2V_276_159),
	.C2V_5 (C2V_276_193),
	.C2V_6 (C2V_276_272),
	.C2V_7 (C2V_276_325),
	.C2V_8 (C2V_276_477),
	.C2V_9 (C2V_276_574),
	.C2V_10 (C2V_276_607),
	.C2V_11 (C2V_276_811),
	.C2V_12 (C2V_276_839),
	.C2V_13 (C2V_276_872),
	.C2V_14 (C2V_276_934),
	.C2V_15 (C2V_276_969),
	.C2V_16 (C2V_276_1036),
	.C2V_17 (C2V_276_1100),
	.C2V_18 (C2V_276_1150),
	.C2V_19 (C2V_276_1427),
	.C2V_20 (C2V_276_1428),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU277 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_3_277),
	.V2C_2 (V2C_87_277),
	.V2C_3 (V2C_107_277),
	.V2C_4 (V2C_168_277),
	.V2C_5 (V2C_230_277),
	.V2C_6 (V2C_273_277),
	.V2C_7 (V2C_373_277),
	.V2C_8 (V2C_427_277),
	.V2C_9 (V2C_524_277),
	.V2C_10 (V2C_760_277),
	.V2C_11 (V2C_808_277),
	.V2C_12 (V2C_856_277),
	.V2C_13 (V2C_897_277),
	.V2C_14 (V2C_938_277),
	.V2C_15 (V2C_972_277),
	.V2C_16 (V2C_1011_277),
	.V2C_17 (V2C_1085_277),
	.V2C_18 (V2C_1144_277),
	.V2C_19 (V2C_1428_277),
	.V2C_20 (V2C_1429_277),
	.C2V_1 (C2V_277_3),
	.C2V_2 (C2V_277_87),
	.C2V_3 (C2V_277_107),
	.C2V_4 (C2V_277_168),
	.C2V_5 (C2V_277_230),
	.C2V_6 (C2V_277_273),
	.C2V_7 (C2V_277_373),
	.C2V_8 (C2V_277_427),
	.C2V_9 (C2V_277_524),
	.C2V_10 (C2V_277_760),
	.C2V_11 (C2V_277_808),
	.C2V_12 (C2V_277_856),
	.C2V_13 (C2V_277_897),
	.C2V_14 (C2V_277_938),
	.C2V_15 (C2V_277_972),
	.C2V_16 (C2V_277_1011),
	.C2V_17 (C2V_277_1085),
	.C2V_18 (C2V_277_1144),
	.C2V_19 (C2V_277_1428),
	.C2V_20 (C2V_277_1429),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU278 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_12_278),
	.V2C_2 (V2C_61_278),
	.V2C_3 (V2C_117_278),
	.V2C_4 (V2C_165_278),
	.V2C_5 (V2C_194_278),
	.V2C_6 (V2C_263_278),
	.V2C_7 (V2C_314_278),
	.V2C_8 (V2C_421_278),
	.V2C_9 (V2C_510_278),
	.V2C_10 (V2C_670_278),
	.V2C_11 (V2C_683_278),
	.V2C_12 (V2C_851_278),
	.V2C_13 (V2C_893_278),
	.V2C_14 (V2C_956_278),
	.V2C_15 (V2C_987_278),
	.V2C_16 (V2C_1019_278),
	.V2C_17 (V2C_1086_278),
	.V2C_18 (V2C_1117_278),
	.V2C_19 (V2C_1429_278),
	.V2C_20 (V2C_1430_278),
	.C2V_1 (C2V_278_12),
	.C2V_2 (C2V_278_61),
	.C2V_3 (C2V_278_117),
	.C2V_4 (C2V_278_165),
	.C2V_5 (C2V_278_194),
	.C2V_6 (C2V_278_263),
	.C2V_7 (C2V_278_314),
	.C2V_8 (C2V_278_421),
	.C2V_9 (C2V_278_510),
	.C2V_10 (C2V_278_670),
	.C2V_11 (C2V_278_683),
	.C2V_12 (C2V_278_851),
	.C2V_13 (C2V_278_893),
	.C2V_14 (C2V_278_956),
	.C2V_15 (C2V_278_987),
	.C2V_16 (C2V_278_1019),
	.C2V_17 (C2V_278_1086),
	.C2V_18 (C2V_278_1117),
	.C2V_19 (C2V_278_1429),
	.C2V_20 (C2V_278_1430),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU279 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_7_279),
	.V2C_2 (V2C_82_279),
	.V2C_3 (V2C_99_279),
	.V2C_4 (V2C_181_279),
	.V2C_5 (V2C_199_279),
	.V2C_6 (V2C_266_279),
	.V2C_7 (V2C_363_279),
	.V2C_8 (V2C_418_279),
	.V2C_9 (V2C_529_279),
	.V2C_10 (V2C_586_279),
	.V2C_11 (V2C_662_279),
	.V2C_12 (V2C_766_279),
	.V2C_13 (V2C_897_279),
	.V2C_14 (V2C_941_279),
	.V2C_15 (V2C_966_279),
	.V2C_16 (V2C_1026_279),
	.V2C_17 (V2C_1104_279),
	.V2C_18 (V2C_1149_279),
	.V2C_19 (V2C_1430_279),
	.V2C_20 (V2C_1431_279),
	.C2V_1 (C2V_279_7),
	.C2V_2 (C2V_279_82),
	.C2V_3 (C2V_279_99),
	.C2V_4 (C2V_279_181),
	.C2V_5 (C2V_279_199),
	.C2V_6 (C2V_279_266),
	.C2V_7 (C2V_279_363),
	.C2V_8 (C2V_279_418),
	.C2V_9 (C2V_279_529),
	.C2V_10 (C2V_279_586),
	.C2V_11 (C2V_279_662),
	.C2V_12 (C2V_279_766),
	.C2V_13 (C2V_279_897),
	.C2V_14 (C2V_279_941),
	.C2V_15 (C2V_279_966),
	.C2V_16 (C2V_279_1026),
	.C2V_17 (C2V_279_1104),
	.C2V_18 (C2V_279_1149),
	.C2V_19 (C2V_279_1430),
	.C2V_20 (C2V_279_1431),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU280 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_26_280),
	.V2C_2 (V2C_85_280),
	.V2C_3 (V2C_124_280),
	.V2C_4 (V2C_180_280),
	.V2C_5 (V2C_197_280),
	.V2C_6 (V2C_251_280),
	.V2C_7 (V2C_475_280),
	.V2C_8 (V2C_515_280),
	.V2C_9 (V2C_551_280),
	.V2C_10 (V2C_613_280),
	.V2C_11 (V2C_638_280),
	.V2C_12 (V2C_684_280),
	.V2C_13 (V2C_901_280),
	.V2C_14 (V2C_925_280),
	.V2C_15 (V2C_961_280),
	.V2C_16 (V2C_1039_280),
	.V2C_17 (V2C_1066_280),
	.V2C_18 (V2C_1130_280),
	.V2C_19 (V2C_1431_280),
	.V2C_20 (V2C_1432_280),
	.C2V_1 (C2V_280_26),
	.C2V_2 (C2V_280_85),
	.C2V_3 (C2V_280_124),
	.C2V_4 (C2V_280_180),
	.C2V_5 (C2V_280_197),
	.C2V_6 (C2V_280_251),
	.C2V_7 (C2V_280_475),
	.C2V_8 (C2V_280_515),
	.C2V_9 (C2V_280_551),
	.C2V_10 (C2V_280_613),
	.C2V_11 (C2V_280_638),
	.C2V_12 (C2V_280_684),
	.C2V_13 (C2V_280_901),
	.C2V_14 (C2V_280_925),
	.C2V_15 (C2V_280_961),
	.C2V_16 (C2V_280_1039),
	.C2V_17 (C2V_280_1066),
	.C2V_18 (C2V_280_1130),
	.C2V_19 (C2V_280_1431),
	.C2V_20 (C2V_280_1432),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU281 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_45_281),
	.V2C_2 (V2C_55_281),
	.V2C_3 (V2C_138_281),
	.V2C_4 (V2C_161_281),
	.V2C_5 (V2C_225_281),
	.V2C_6 (V2C_243_281),
	.V2C_7 (V2C_292_281),
	.V2C_8 (V2C_359_281),
	.V2C_9 (V2C_438_281),
	.V2C_10 (V2C_720_281),
	.V2C_11 (V2C_736_281),
	.V2C_12 (V2C_790_281),
	.V2C_13 (V2C_868_281),
	.V2C_14 (V2C_916_281),
	.V2C_15 (V2C_1007_281),
	.V2C_16 (V2C_1011_281),
	.V2C_17 (V2C_1060_281),
	.V2C_18 (V2C_1108_281),
	.V2C_19 (V2C_1432_281),
	.V2C_20 (V2C_1433_281),
	.C2V_1 (C2V_281_45),
	.C2V_2 (C2V_281_55),
	.C2V_3 (C2V_281_138),
	.C2V_4 (C2V_281_161),
	.C2V_5 (C2V_281_225),
	.C2V_6 (C2V_281_243),
	.C2V_7 (C2V_281_292),
	.C2V_8 (C2V_281_359),
	.C2V_9 (C2V_281_438),
	.C2V_10 (C2V_281_720),
	.C2V_11 (C2V_281_736),
	.C2V_12 (C2V_281_790),
	.C2V_13 (C2V_281_868),
	.C2V_14 (C2V_281_916),
	.C2V_15 (C2V_281_1007),
	.C2V_16 (C2V_281_1011),
	.C2V_17 (C2V_281_1060),
	.C2V_18 (C2V_281_1108),
	.C2V_19 (C2V_281_1432),
	.C2V_20 (C2V_281_1433),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU282 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_28_282),
	.V2C_2 (V2C_52_282),
	.V2C_3 (V2C_140_282),
	.V2C_4 (V2C_160_282),
	.V2C_5 (V2C_194_282),
	.V2C_6 (V2C_273_282),
	.V2C_7 (V2C_326_282),
	.V2C_8 (V2C_478_282),
	.V2C_9 (V2C_575_282),
	.V2C_10 (V2C_608_282),
	.V2C_11 (V2C_812_282),
	.V2C_12 (V2C_840_282),
	.V2C_13 (V2C_873_282),
	.V2C_14 (V2C_935_282),
	.V2C_15 (V2C_970_282),
	.V2C_16 (V2C_1037_282),
	.V2C_17 (V2C_1101_282),
	.V2C_18 (V2C_1151_282),
	.V2C_19 (V2C_1433_282),
	.V2C_20 (V2C_1434_282),
	.C2V_1 (C2V_282_28),
	.C2V_2 (C2V_282_52),
	.C2V_3 (C2V_282_140),
	.C2V_4 (C2V_282_160),
	.C2V_5 (C2V_282_194),
	.C2V_6 (C2V_282_273),
	.C2V_7 (C2V_282_326),
	.C2V_8 (C2V_282_478),
	.C2V_9 (C2V_282_575),
	.C2V_10 (C2V_282_608),
	.C2V_11 (C2V_282_812),
	.C2V_12 (C2V_282_840),
	.C2V_13 (C2V_282_873),
	.C2V_14 (C2V_282_935),
	.C2V_15 (C2V_282_970),
	.C2V_16 (C2V_282_1037),
	.C2V_17 (C2V_282_1101),
	.C2V_18 (C2V_282_1151),
	.C2V_19 (C2V_282_1433),
	.C2V_20 (C2V_282_1434),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU283 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_4_283),
	.V2C_2 (V2C_88_283),
	.V2C_3 (V2C_108_283),
	.V2C_4 (V2C_169_283),
	.V2C_5 (V2C_231_283),
	.V2C_6 (V2C_274_283),
	.V2C_7 (V2C_374_283),
	.V2C_8 (V2C_428_283),
	.V2C_9 (V2C_525_283),
	.V2C_10 (V2C_761_283),
	.V2C_11 (V2C_809_283),
	.V2C_12 (V2C_857_283),
	.V2C_13 (V2C_898_283),
	.V2C_14 (V2C_939_283),
	.V2C_15 (V2C_973_283),
	.V2C_16 (V2C_1012_283),
	.V2C_17 (V2C_1086_283),
	.V2C_18 (V2C_1145_283),
	.V2C_19 (V2C_1434_283),
	.V2C_20 (V2C_1435_283),
	.C2V_1 (C2V_283_4),
	.C2V_2 (C2V_283_88),
	.C2V_3 (C2V_283_108),
	.C2V_4 (C2V_283_169),
	.C2V_5 (C2V_283_231),
	.C2V_6 (C2V_283_274),
	.C2V_7 (C2V_283_374),
	.C2V_8 (C2V_283_428),
	.C2V_9 (C2V_283_525),
	.C2V_10 (C2V_283_761),
	.C2V_11 (C2V_283_809),
	.C2V_12 (C2V_283_857),
	.C2V_13 (C2V_283_898),
	.C2V_14 (C2V_283_939),
	.C2V_15 (C2V_283_973),
	.C2V_16 (C2V_283_1012),
	.C2V_17 (C2V_283_1086),
	.C2V_18 (C2V_283_1145),
	.C2V_19 (C2V_283_1434),
	.C2V_20 (C2V_283_1435),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU284 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_13_284),
	.V2C_2 (V2C_62_284),
	.V2C_3 (V2C_118_284),
	.V2C_4 (V2C_166_284),
	.V2C_5 (V2C_195_284),
	.V2C_6 (V2C_264_284),
	.V2C_7 (V2C_315_284),
	.V2C_8 (V2C_422_284),
	.V2C_9 (V2C_511_284),
	.V2C_10 (V2C_671_284),
	.V2C_11 (V2C_684_284),
	.V2C_12 (V2C_852_284),
	.V2C_13 (V2C_894_284),
	.V2C_14 (V2C_957_284),
	.V2C_15 (V2C_988_284),
	.V2C_16 (V2C_1020_284),
	.V2C_17 (V2C_1087_284),
	.V2C_18 (V2C_1118_284),
	.V2C_19 (V2C_1435_284),
	.V2C_20 (V2C_1436_284),
	.C2V_1 (C2V_284_13),
	.C2V_2 (C2V_284_62),
	.C2V_3 (C2V_284_118),
	.C2V_4 (C2V_284_166),
	.C2V_5 (C2V_284_195),
	.C2V_6 (C2V_284_264),
	.C2V_7 (C2V_284_315),
	.C2V_8 (C2V_284_422),
	.C2V_9 (C2V_284_511),
	.C2V_10 (C2V_284_671),
	.C2V_11 (C2V_284_684),
	.C2V_12 (C2V_284_852),
	.C2V_13 (C2V_284_894),
	.C2V_14 (C2V_284_957),
	.C2V_15 (C2V_284_988),
	.C2V_16 (C2V_284_1020),
	.C2V_17 (C2V_284_1087),
	.C2V_18 (C2V_284_1118),
	.C2V_19 (C2V_284_1435),
	.C2V_20 (C2V_284_1436),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU285 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_8_285),
	.V2C_2 (V2C_83_285),
	.V2C_3 (V2C_100_285),
	.V2C_4 (V2C_182_285),
	.V2C_5 (V2C_200_285),
	.V2C_6 (V2C_267_285),
	.V2C_7 (V2C_364_285),
	.V2C_8 (V2C_419_285),
	.V2C_9 (V2C_530_285),
	.V2C_10 (V2C_587_285),
	.V2C_11 (V2C_663_285),
	.V2C_12 (V2C_767_285),
	.V2C_13 (V2C_898_285),
	.V2C_14 (V2C_942_285),
	.V2C_15 (V2C_967_285),
	.V2C_16 (V2C_1027_285),
	.V2C_17 (V2C_1057_285),
	.V2C_18 (V2C_1150_285),
	.V2C_19 (V2C_1436_285),
	.V2C_20 (V2C_1437_285),
	.C2V_1 (C2V_285_8),
	.C2V_2 (C2V_285_83),
	.C2V_3 (C2V_285_100),
	.C2V_4 (C2V_285_182),
	.C2V_5 (C2V_285_200),
	.C2V_6 (C2V_285_267),
	.C2V_7 (C2V_285_364),
	.C2V_8 (C2V_285_419),
	.C2V_9 (C2V_285_530),
	.C2V_10 (C2V_285_587),
	.C2V_11 (C2V_285_663),
	.C2V_12 (C2V_285_767),
	.C2V_13 (C2V_285_898),
	.C2V_14 (C2V_285_942),
	.C2V_15 (C2V_285_967),
	.C2V_16 (C2V_285_1027),
	.C2V_17 (C2V_285_1057),
	.C2V_18 (C2V_285_1150),
	.C2V_19 (C2V_285_1436),
	.C2V_20 (C2V_285_1437),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU286 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_27_286),
	.V2C_2 (V2C_86_286),
	.V2C_3 (V2C_125_286),
	.V2C_4 (V2C_181_286),
	.V2C_5 (V2C_198_286),
	.V2C_6 (V2C_252_286),
	.V2C_7 (V2C_476_286),
	.V2C_8 (V2C_516_286),
	.V2C_9 (V2C_552_286),
	.V2C_10 (V2C_614_286),
	.V2C_11 (V2C_639_286),
	.V2C_12 (V2C_685_286),
	.V2C_13 (V2C_902_286),
	.V2C_14 (V2C_926_286),
	.V2C_15 (V2C_962_286),
	.V2C_16 (V2C_1040_286),
	.V2C_17 (V2C_1067_286),
	.V2C_18 (V2C_1131_286),
	.V2C_19 (V2C_1437_286),
	.V2C_20 (V2C_1438_286),
	.C2V_1 (C2V_286_27),
	.C2V_2 (C2V_286_86),
	.C2V_3 (C2V_286_125),
	.C2V_4 (C2V_286_181),
	.C2V_5 (C2V_286_198),
	.C2V_6 (C2V_286_252),
	.C2V_7 (C2V_286_476),
	.C2V_8 (C2V_286_516),
	.C2V_9 (C2V_286_552),
	.C2V_10 (C2V_286_614),
	.C2V_11 (C2V_286_639),
	.C2V_12 (C2V_286_685),
	.C2V_13 (C2V_286_902),
	.C2V_14 (C2V_286_926),
	.C2V_15 (C2V_286_962),
	.C2V_16 (C2V_286_1040),
	.C2V_17 (C2V_286_1067),
	.C2V_18 (C2V_286_1131),
	.C2V_19 (C2V_286_1437),
	.C2V_20 (C2V_286_1438),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU287 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_46_287),
	.V2C_2 (V2C_56_287),
	.V2C_3 (V2C_139_287),
	.V2C_4 (V2C_162_287),
	.V2C_5 (V2C_226_287),
	.V2C_6 (V2C_244_287),
	.V2C_7 (V2C_293_287),
	.V2C_8 (V2C_360_287),
	.V2C_9 (V2C_439_287),
	.V2C_10 (V2C_673_287),
	.V2C_11 (V2C_737_287),
	.V2C_12 (V2C_791_287),
	.V2C_13 (V2C_869_287),
	.V2C_14 (V2C_917_287),
	.V2C_15 (V2C_1008_287),
	.V2C_16 (V2C_1012_287),
	.V2C_17 (V2C_1061_287),
	.V2C_18 (V2C_1109_287),
	.V2C_19 (V2C_1438_287),
	.V2C_20 (V2C_1439_287),
	.C2V_1 (C2V_287_46),
	.C2V_2 (C2V_287_56),
	.C2V_3 (C2V_287_139),
	.C2V_4 (C2V_287_162),
	.C2V_5 (C2V_287_226),
	.C2V_6 (C2V_287_244),
	.C2V_7 (C2V_287_293),
	.C2V_8 (C2V_287_360),
	.C2V_9 (C2V_287_439),
	.C2V_10 (C2V_287_673),
	.C2V_11 (C2V_287_737),
	.C2V_12 (C2V_287_791),
	.C2V_13 (C2V_287_869),
	.C2V_14 (C2V_287_917),
	.C2V_15 (C2V_287_1008),
	.C2V_16 (C2V_287_1012),
	.C2V_17 (C2V_287_1061),
	.C2V_18 (C2V_287_1109),
	.C2V_19 (C2V_287_1438),
	.C2V_20 (C2V_287_1439),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU288 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_29_288),
	.V2C_2 (V2C_53_288),
	.V2C_3 (V2C_141_288),
	.V2C_4 (V2C_161_288),
	.V2C_5 (V2C_195_288),
	.V2C_6 (V2C_274_288),
	.V2C_7 (V2C_327_288),
	.V2C_8 (V2C_479_288),
	.V2C_9 (V2C_576_288),
	.V2C_10 (V2C_609_288),
	.V2C_11 (V2C_813_288),
	.V2C_12 (V2C_841_288),
	.V2C_13 (V2C_874_288),
	.V2C_14 (V2C_936_288),
	.V2C_15 (V2C_971_288),
	.V2C_16 (V2C_1038_288),
	.V2C_17 (V2C_1102_288),
	.V2C_18 (V2C_1152_288),
	.V2C_19 (V2C_1439_288),
	.V2C_20 (V2C_1440_288),
	.C2V_1 (C2V_288_29),
	.C2V_2 (C2V_288_53),
	.C2V_3 (C2V_288_141),
	.C2V_4 (C2V_288_161),
	.C2V_5 (C2V_288_195),
	.C2V_6 (C2V_288_274),
	.C2V_7 (C2V_288_327),
	.C2V_8 (C2V_288_479),
	.C2V_9 (C2V_288_576),
	.C2V_10 (C2V_288_609),
	.C2V_11 (C2V_288_813),
	.C2V_12 (C2V_288_841),
	.C2V_13 (C2V_288_874),
	.C2V_14 (C2V_288_936),
	.C2V_15 (C2V_288_971),
	.C2V_16 (C2V_288_1038),
	.C2V_17 (C2V_288_1102),
	.C2V_18 (C2V_288_1152),
	.C2V_19 (C2V_288_1439),
	.C2V_20 (C2V_288_1440),
	.init_cnt (8'd2)
);

VNU_6 #(quan_width) VNU1 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_1),
	.C2V_2 (C2V_120_1),
	.C2V_3 (C2V_130_1),
	.C2V_4 (C2V_212_1),
	.C2V_5 (C2V_243_1),
	.C2V_6 (C2V_265_1),
	.L (L[14:0]),
	.V2C_1 (V2C_1_17),
	.V2C_2 (V2C_1_120),
	.V2C_3 (V2C_1_130),
	.V2C_4 (V2C_1_212),
	.V2C_5 (V2C_1_243),
	.V2C_6 (V2C_1_265),
	.V (V_1)
);

VNU_6 #(quan_width) VNU2 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_2),
	.C2V_2 (C2V_126_2),
	.C2V_3 (C2V_136_2),
	.C2V_4 (C2V_218_2),
	.C2V_5 (C2V_249_2),
	.C2V_6 (C2V_271_2),
	.L (L[29:15]),
	.V2C_1 (V2C_2_23),
	.V2C_2 (V2C_2_126),
	.V2C_3 (V2C_2_136),
	.V2C_4 (V2C_2_218),
	.V2C_5 (V2C_2_249),
	.V2C_6 (V2C_2_271),
	.V (V_2)
);

VNU_6 #(quan_width) VNU3 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_3),
	.C2V_2 (C2V_132_3),
	.C2V_3 (C2V_142_3),
	.C2V_4 (C2V_224_3),
	.C2V_5 (C2V_255_3),
	.C2V_6 (C2V_277_3),
	.L (L[44:30]),
	.V2C_1 (V2C_3_29),
	.V2C_2 (V2C_3_132),
	.V2C_3 (V2C_3_142),
	.V2C_4 (V2C_3_224),
	.V2C_5 (V2C_3_255),
	.V2C_6 (V2C_3_277),
	.V (V_3)
);

VNU_6 #(quan_width) VNU4 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_4),
	.C2V_2 (C2V_138_4),
	.C2V_3 (C2V_148_4),
	.C2V_4 (C2V_230_4),
	.C2V_5 (C2V_261_4),
	.C2V_6 (C2V_283_4),
	.L (L[59:45]),
	.V2C_1 (V2C_4_35),
	.V2C_2 (V2C_4_138),
	.V2C_3 (V2C_4_148),
	.V2C_4 (V2C_4_230),
	.V2C_5 (V2C_4_261),
	.V2C_6 (V2C_4_283),
	.V (V_4)
);

VNU_6 #(quan_width) VNU5 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_5),
	.C2V_2 (C2V_41_5),
	.C2V_3 (C2V_144_5),
	.C2V_4 (C2V_154_5),
	.C2V_5 (C2V_236_5),
	.C2V_6 (C2V_267_5),
	.L (L[74:60]),
	.V2C_1 (V2C_5_1),
	.V2C_2 (V2C_5_41),
	.V2C_3 (V2C_5_144),
	.V2C_4 (V2C_5_154),
	.V2C_5 (V2C_5_236),
	.V2C_6 (V2C_5_267),
	.V (V_5)
);

VNU_6 #(quan_width) VNU6 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_6),
	.C2V_2 (C2V_47_6),
	.C2V_3 (C2V_150_6),
	.C2V_4 (C2V_160_6),
	.C2V_5 (C2V_242_6),
	.C2V_6 (C2V_273_6),
	.L (L[89:75]),
	.V2C_1 (V2C_6_7),
	.V2C_2 (V2C_6_47),
	.V2C_3 (V2C_6_150),
	.V2C_4 (V2C_6_160),
	.V2C_5 (V2C_6_242),
	.V2C_6 (V2C_6_273),
	.V (V_6)
);

VNU_6 #(quan_width) VNU7 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_7),
	.C2V_2 (C2V_53_7),
	.C2V_3 (C2V_156_7),
	.C2V_4 (C2V_166_7),
	.C2V_5 (C2V_248_7),
	.C2V_6 (C2V_279_7),
	.L (L[104:90]),
	.V2C_1 (V2C_7_13),
	.V2C_2 (V2C_7_53),
	.V2C_3 (V2C_7_156),
	.V2C_4 (V2C_7_166),
	.V2C_5 (V2C_7_248),
	.V2C_6 (V2C_7_279),
	.V (V_7)
);

VNU_6 #(quan_width) VNU8 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_8),
	.C2V_2 (C2V_59_8),
	.C2V_3 (C2V_162_8),
	.C2V_4 (C2V_172_8),
	.C2V_5 (C2V_254_8),
	.C2V_6 (C2V_285_8),
	.L (L[119:105]),
	.V2C_1 (V2C_8_19),
	.V2C_2 (V2C_8_59),
	.V2C_3 (V2C_8_162),
	.V2C_4 (V2C_8_172),
	.V2C_5 (V2C_8_254),
	.V2C_6 (V2C_8_285),
	.V (V_8)
);

VNU_6 #(quan_width) VNU9 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_9),
	.C2V_2 (C2V_25_9),
	.C2V_3 (C2V_65_9),
	.C2V_4 (C2V_168_9),
	.C2V_5 (C2V_178_9),
	.C2V_6 (C2V_260_9),
	.L (L[134:120]),
	.V2C_1 (V2C_9_3),
	.V2C_2 (V2C_9_25),
	.V2C_3 (V2C_9_65),
	.V2C_4 (V2C_9_168),
	.V2C_5 (V2C_9_178),
	.V2C_6 (V2C_9_260),
	.V (V_9)
);

VNU_6 #(quan_width) VNU10 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_10),
	.C2V_2 (C2V_31_10),
	.C2V_3 (C2V_71_10),
	.C2V_4 (C2V_174_10),
	.C2V_5 (C2V_184_10),
	.C2V_6 (C2V_266_10),
	.L (L[149:135]),
	.V2C_1 (V2C_10_9),
	.V2C_2 (V2C_10_31),
	.V2C_3 (V2C_10_71),
	.V2C_4 (V2C_10_174),
	.V2C_5 (V2C_10_184),
	.V2C_6 (V2C_10_266),
	.V (V_10)
);

VNU_6 #(quan_width) VNU11 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_11),
	.C2V_2 (C2V_37_11),
	.C2V_3 (C2V_77_11),
	.C2V_4 (C2V_180_11),
	.C2V_5 (C2V_190_11),
	.C2V_6 (C2V_272_11),
	.L (L[164:150]),
	.V2C_1 (V2C_11_15),
	.V2C_2 (V2C_11_37),
	.V2C_3 (V2C_11_77),
	.V2C_4 (V2C_11_180),
	.V2C_5 (V2C_11_190),
	.V2C_6 (V2C_11_272),
	.V (V_11)
);

VNU_6 #(quan_width) VNU12 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_12),
	.C2V_2 (C2V_43_12),
	.C2V_3 (C2V_83_12),
	.C2V_4 (C2V_186_12),
	.C2V_5 (C2V_196_12),
	.C2V_6 (C2V_278_12),
	.L (L[179:165]),
	.V2C_1 (V2C_12_21),
	.V2C_2 (V2C_12_43),
	.V2C_3 (V2C_12_83),
	.V2C_4 (V2C_12_186),
	.V2C_5 (V2C_12_196),
	.V2C_6 (V2C_12_278),
	.V (V_12)
);

VNU_6 #(quan_width) VNU13 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_13),
	.C2V_2 (C2V_49_13),
	.C2V_3 (C2V_89_13),
	.C2V_4 (C2V_192_13),
	.C2V_5 (C2V_202_13),
	.C2V_6 (C2V_284_13),
	.L (L[194:180]),
	.V2C_1 (V2C_13_27),
	.V2C_2 (V2C_13_49),
	.V2C_3 (V2C_13_89),
	.V2C_4 (V2C_13_192),
	.V2C_5 (V2C_13_202),
	.V2C_6 (V2C_13_284),
	.V (V_13)
);

VNU_6 #(quan_width) VNU14 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_14),
	.C2V_2 (C2V_33_14),
	.C2V_3 (C2V_55_14),
	.C2V_4 (C2V_95_14),
	.C2V_5 (C2V_198_14),
	.C2V_6 (C2V_208_14),
	.L (L[209:195]),
	.V2C_1 (V2C_14_2),
	.V2C_2 (V2C_14_33),
	.V2C_3 (V2C_14_55),
	.V2C_4 (V2C_14_95),
	.V2C_5 (V2C_14_198),
	.V2C_6 (V2C_14_208),
	.V (V_14)
);

VNU_6 #(quan_width) VNU15 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_15),
	.C2V_2 (C2V_39_15),
	.C2V_3 (C2V_61_15),
	.C2V_4 (C2V_101_15),
	.C2V_5 (C2V_204_15),
	.C2V_6 (C2V_214_15),
	.L (L[224:210]),
	.V2C_1 (V2C_15_8),
	.V2C_2 (V2C_15_39),
	.V2C_3 (V2C_15_61),
	.V2C_4 (V2C_15_101),
	.V2C_5 (V2C_15_204),
	.V2C_6 (V2C_15_214),
	.V (V_15)
);

VNU_6 #(quan_width) VNU16 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_16),
	.C2V_2 (C2V_45_16),
	.C2V_3 (C2V_67_16),
	.C2V_4 (C2V_107_16),
	.C2V_5 (C2V_210_16),
	.C2V_6 (C2V_220_16),
	.L (L[239:225]),
	.V2C_1 (V2C_16_14),
	.V2C_2 (V2C_16_45),
	.V2C_3 (V2C_16_67),
	.V2C_4 (V2C_16_107),
	.V2C_5 (V2C_16_210),
	.V2C_6 (V2C_16_220),
	.V (V_16)
);

VNU_6 #(quan_width) VNU17 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_17),
	.C2V_2 (C2V_51_17),
	.C2V_3 (C2V_73_17),
	.C2V_4 (C2V_113_17),
	.C2V_5 (C2V_216_17),
	.C2V_6 (C2V_226_17),
	.L (L[254:240]),
	.V2C_1 (V2C_17_20),
	.V2C_2 (V2C_17_51),
	.V2C_3 (V2C_17_73),
	.V2C_4 (V2C_17_113),
	.V2C_5 (V2C_17_216),
	.V2C_6 (V2C_17_226),
	.V (V_17)
);

VNU_6 #(quan_width) VNU18 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_18),
	.C2V_2 (C2V_57_18),
	.C2V_3 (C2V_79_18),
	.C2V_4 (C2V_119_18),
	.C2V_5 (C2V_222_18),
	.C2V_6 (C2V_232_18),
	.L (L[269:255]),
	.V2C_1 (V2C_18_26),
	.V2C_2 (V2C_18_57),
	.V2C_3 (V2C_18_79),
	.V2C_4 (V2C_18_119),
	.V2C_5 (V2C_18_222),
	.V2C_6 (V2C_18_232),
	.V (V_18)
);

VNU_6 #(quan_width) VNU19 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_19),
	.C2V_2 (C2V_63_19),
	.C2V_3 (C2V_85_19),
	.C2V_4 (C2V_125_19),
	.C2V_5 (C2V_228_19),
	.C2V_6 (C2V_238_19),
	.L (L[284:270]),
	.V2C_1 (V2C_19_32),
	.V2C_2 (V2C_19_63),
	.V2C_3 (V2C_19_85),
	.V2C_4 (V2C_19_125),
	.V2C_5 (V2C_19_228),
	.V2C_6 (V2C_19_238),
	.V (V_19)
);

VNU_6 #(quan_width) VNU20 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_20),
	.C2V_2 (C2V_69_20),
	.C2V_3 (C2V_91_20),
	.C2V_4 (C2V_131_20),
	.C2V_5 (C2V_234_20),
	.C2V_6 (C2V_244_20),
	.L (L[299:285]),
	.V2C_1 (V2C_20_38),
	.V2C_2 (V2C_20_69),
	.V2C_3 (V2C_20_91),
	.V2C_4 (V2C_20_131),
	.V2C_5 (V2C_20_234),
	.V2C_6 (V2C_20_244),
	.V (V_20)
);

VNU_6 #(quan_width) VNU21 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_21),
	.C2V_2 (C2V_75_21),
	.C2V_3 (C2V_97_21),
	.C2V_4 (C2V_137_21),
	.C2V_5 (C2V_240_21),
	.C2V_6 (C2V_250_21),
	.L (L[314:300]),
	.V2C_1 (V2C_21_44),
	.V2C_2 (V2C_21_75),
	.V2C_3 (V2C_21_97),
	.V2C_4 (V2C_21_137),
	.V2C_5 (V2C_21_240),
	.V2C_6 (V2C_21_250),
	.V (V_21)
);

VNU_6 #(quan_width) VNU22 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_22),
	.C2V_2 (C2V_81_22),
	.C2V_3 (C2V_103_22),
	.C2V_4 (C2V_143_22),
	.C2V_5 (C2V_246_22),
	.C2V_6 (C2V_256_22),
	.L (L[329:315]),
	.V2C_1 (V2C_22_50),
	.V2C_2 (V2C_22_81),
	.V2C_3 (V2C_22_103),
	.V2C_4 (V2C_22_143),
	.V2C_5 (V2C_22_246),
	.V2C_6 (V2C_22_256),
	.V (V_22)
);

VNU_6 #(quan_width) VNU23 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_23),
	.C2V_2 (C2V_87_23),
	.C2V_3 (C2V_109_23),
	.C2V_4 (C2V_149_23),
	.C2V_5 (C2V_252_23),
	.C2V_6 (C2V_262_23),
	.L (L[344:330]),
	.V2C_1 (V2C_23_56),
	.V2C_2 (V2C_23_87),
	.V2C_3 (V2C_23_109),
	.V2C_4 (V2C_23_149),
	.V2C_5 (V2C_23_252),
	.V2C_6 (V2C_23_262),
	.V (V_23)
);

VNU_6 #(quan_width) VNU24 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_24),
	.C2V_2 (C2V_93_24),
	.C2V_3 (C2V_115_24),
	.C2V_4 (C2V_155_24),
	.C2V_5 (C2V_258_24),
	.C2V_6 (C2V_268_24),
	.L (L[359:345]),
	.V2C_1 (V2C_24_62),
	.V2C_2 (V2C_24_93),
	.V2C_3 (V2C_24_115),
	.V2C_4 (V2C_24_155),
	.V2C_5 (V2C_24_258),
	.V2C_6 (V2C_24_268),
	.V (V_24)
);

VNU_6 #(quan_width) VNU25 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_25),
	.C2V_2 (C2V_99_25),
	.C2V_3 (C2V_121_25),
	.C2V_4 (C2V_161_25),
	.C2V_5 (C2V_264_25),
	.C2V_6 (C2V_274_25),
	.L (L[374:360]),
	.V2C_1 (V2C_25_68),
	.V2C_2 (V2C_25_99),
	.V2C_3 (V2C_25_121),
	.V2C_4 (V2C_25_161),
	.V2C_5 (V2C_25_264),
	.V2C_6 (V2C_25_274),
	.V (V_25)
);

VNU_6 #(quan_width) VNU26 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_26),
	.C2V_2 (C2V_105_26),
	.C2V_3 (C2V_127_26),
	.C2V_4 (C2V_167_26),
	.C2V_5 (C2V_270_26),
	.C2V_6 (C2V_280_26),
	.L (L[389:375]),
	.V2C_1 (V2C_26_74),
	.V2C_2 (V2C_26_105),
	.V2C_3 (V2C_26_127),
	.V2C_4 (V2C_26_167),
	.V2C_5 (V2C_26_270),
	.V2C_6 (V2C_26_280),
	.V (V_26)
);

VNU_6 #(quan_width) VNU27 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_80_27),
	.C2V_2 (C2V_111_27),
	.C2V_3 (C2V_133_27),
	.C2V_4 (C2V_173_27),
	.C2V_5 (C2V_276_27),
	.C2V_6 (C2V_286_27),
	.L (L[404:390]),
	.V2C_1 (V2C_27_80),
	.V2C_2 (V2C_27_111),
	.V2C_3 (V2C_27_133),
	.V2C_4 (V2C_27_173),
	.V2C_5 (V2C_27_276),
	.V2C_6 (V2C_27_286),
	.V (V_27)
);

VNU_6 #(quan_width) VNU28 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_28),
	.C2V_2 (C2V_86_28),
	.C2V_3 (C2V_117_28),
	.C2V_4 (C2V_139_28),
	.C2V_5 (C2V_179_28),
	.C2V_6 (C2V_282_28),
	.L (L[419:405]),
	.V2C_1 (V2C_28_4),
	.V2C_2 (V2C_28_86),
	.V2C_3 (V2C_28_117),
	.V2C_4 (V2C_28_139),
	.V2C_5 (V2C_28_179),
	.V2C_6 (V2C_28_282),
	.V (V_28)
);

VNU_6 #(quan_width) VNU29 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_29),
	.C2V_2 (C2V_92_29),
	.C2V_3 (C2V_123_29),
	.C2V_4 (C2V_145_29),
	.C2V_5 (C2V_185_29),
	.C2V_6 (C2V_288_29),
	.L (L[434:420]),
	.V2C_1 (V2C_29_10),
	.V2C_2 (V2C_29_92),
	.V2C_3 (V2C_29_123),
	.V2C_4 (V2C_29_145),
	.V2C_5 (V2C_29_185),
	.V2C_6 (V2C_29_288),
	.V (V_29)
);

VNU_6 #(quan_width) VNU30 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_30),
	.C2V_2 (C2V_16_30),
	.C2V_3 (C2V_98_30),
	.C2V_4 (C2V_129_30),
	.C2V_5 (C2V_151_30),
	.C2V_6 (C2V_191_30),
	.L (L[449:435]),
	.V2C_1 (V2C_30_6),
	.V2C_2 (V2C_30_16),
	.V2C_3 (V2C_30_98),
	.V2C_4 (V2C_30_129),
	.V2C_5 (V2C_30_151),
	.V2C_6 (V2C_30_191),
	.V (V_30)
);

VNU_6 #(quan_width) VNU31 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_31),
	.C2V_2 (C2V_22_31),
	.C2V_3 (C2V_104_31),
	.C2V_4 (C2V_135_31),
	.C2V_5 (C2V_157_31),
	.C2V_6 (C2V_197_31),
	.L (L[464:450]),
	.V2C_1 (V2C_31_12),
	.V2C_2 (V2C_31_22),
	.V2C_3 (V2C_31_104),
	.V2C_4 (V2C_31_135),
	.V2C_5 (V2C_31_157),
	.V2C_6 (V2C_31_197),
	.V (V_31)
);

VNU_6 #(quan_width) VNU32 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_32),
	.C2V_2 (C2V_28_32),
	.C2V_3 (C2V_110_32),
	.C2V_4 (C2V_141_32),
	.C2V_5 (C2V_163_32),
	.C2V_6 (C2V_203_32),
	.L (L[479:465]),
	.V2C_1 (V2C_32_18),
	.V2C_2 (V2C_32_28),
	.V2C_3 (V2C_32_110),
	.V2C_4 (V2C_32_141),
	.V2C_5 (V2C_32_163),
	.V2C_6 (V2C_32_203),
	.V (V_32)
);

VNU_6 #(quan_width) VNU33 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_33),
	.C2V_2 (C2V_34_33),
	.C2V_3 (C2V_116_33),
	.C2V_4 (C2V_147_33),
	.C2V_5 (C2V_169_33),
	.C2V_6 (C2V_209_33),
	.L (L[494:480]),
	.V2C_1 (V2C_33_24),
	.V2C_2 (V2C_33_34),
	.V2C_3 (V2C_33_116),
	.V2C_4 (V2C_33_147),
	.V2C_5 (V2C_33_169),
	.V2C_6 (V2C_33_209),
	.V (V_33)
);

VNU_6 #(quan_width) VNU34 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_34),
	.C2V_2 (C2V_40_34),
	.C2V_3 (C2V_122_34),
	.C2V_4 (C2V_153_34),
	.C2V_5 (C2V_175_34),
	.C2V_6 (C2V_215_34),
	.L (L[509:495]),
	.V2C_1 (V2C_34_30),
	.V2C_2 (V2C_34_40),
	.V2C_3 (V2C_34_122),
	.V2C_4 (V2C_34_153),
	.V2C_5 (V2C_34_175),
	.V2C_6 (V2C_34_215),
	.V (V_34)
);

VNU_6 #(quan_width) VNU35 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_35),
	.C2V_2 (C2V_46_35),
	.C2V_3 (C2V_128_35),
	.C2V_4 (C2V_159_35),
	.C2V_5 (C2V_181_35),
	.C2V_6 (C2V_221_35),
	.L (L[524:510]),
	.V2C_1 (V2C_35_36),
	.V2C_2 (V2C_35_46),
	.V2C_3 (V2C_35_128),
	.V2C_4 (V2C_35_159),
	.V2C_5 (V2C_35_181),
	.V2C_6 (V2C_35_221),
	.V (V_35)
);

VNU_6 #(quan_width) VNU36 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_36),
	.C2V_2 (C2V_52_36),
	.C2V_3 (C2V_134_36),
	.C2V_4 (C2V_165_36),
	.C2V_5 (C2V_187_36),
	.C2V_6 (C2V_227_36),
	.L (L[539:525]),
	.V2C_1 (V2C_36_42),
	.V2C_2 (V2C_36_52),
	.V2C_3 (V2C_36_134),
	.V2C_4 (V2C_36_165),
	.V2C_5 (V2C_36_187),
	.V2C_6 (V2C_36_227),
	.V (V_36)
);

VNU_6 #(quan_width) VNU37 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_37),
	.C2V_2 (C2V_58_37),
	.C2V_3 (C2V_140_37),
	.C2V_4 (C2V_171_37),
	.C2V_5 (C2V_193_37),
	.C2V_6 (C2V_233_37),
	.L (L[554:540]),
	.V2C_1 (V2C_37_48),
	.V2C_2 (V2C_37_58),
	.V2C_3 (V2C_37_140),
	.V2C_4 (V2C_37_171),
	.V2C_5 (V2C_37_193),
	.V2C_6 (V2C_37_233),
	.V (V_37)
);

VNU_6 #(quan_width) VNU38 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_54_38),
	.C2V_2 (C2V_64_38),
	.C2V_3 (C2V_146_38),
	.C2V_4 (C2V_177_38),
	.C2V_5 (C2V_199_38),
	.C2V_6 (C2V_239_38),
	.L (L[569:555]),
	.V2C_1 (V2C_38_54),
	.V2C_2 (V2C_38_64),
	.V2C_3 (V2C_38_146),
	.V2C_4 (V2C_38_177),
	.V2C_5 (V2C_38_199),
	.V2C_6 (V2C_38_239),
	.V (V_38)
);

VNU_6 #(quan_width) VNU39 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_60_39),
	.C2V_2 (C2V_70_39),
	.C2V_3 (C2V_152_39),
	.C2V_4 (C2V_183_39),
	.C2V_5 (C2V_205_39),
	.C2V_6 (C2V_245_39),
	.L (L[584:570]),
	.V2C_1 (V2C_39_60),
	.V2C_2 (V2C_39_70),
	.V2C_3 (V2C_39_152),
	.V2C_4 (V2C_39_183),
	.V2C_5 (V2C_39_205),
	.V2C_6 (V2C_39_245),
	.V (V_39)
);

VNU_6 #(quan_width) VNU40 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_66_40),
	.C2V_2 (C2V_76_40),
	.C2V_3 (C2V_158_40),
	.C2V_4 (C2V_189_40),
	.C2V_5 (C2V_211_40),
	.C2V_6 (C2V_251_40),
	.L (L[599:585]),
	.V2C_1 (V2C_40_66),
	.V2C_2 (V2C_40_76),
	.V2C_3 (V2C_40_158),
	.V2C_4 (V2C_40_189),
	.V2C_5 (V2C_40_211),
	.V2C_6 (V2C_40_251),
	.V (V_40)
);

VNU_6 #(quan_width) VNU41 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_72_41),
	.C2V_2 (C2V_82_41),
	.C2V_3 (C2V_164_41),
	.C2V_4 (C2V_195_41),
	.C2V_5 (C2V_217_41),
	.C2V_6 (C2V_257_41),
	.L (L[614:600]),
	.V2C_1 (V2C_41_72),
	.V2C_2 (V2C_41_82),
	.V2C_3 (V2C_41_164),
	.V2C_4 (V2C_41_195),
	.V2C_5 (V2C_41_217),
	.V2C_6 (V2C_41_257),
	.V (V_41)
);

VNU_6 #(quan_width) VNU42 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_78_42),
	.C2V_2 (C2V_88_42),
	.C2V_3 (C2V_170_42),
	.C2V_4 (C2V_201_42),
	.C2V_5 (C2V_223_42),
	.C2V_6 (C2V_263_42),
	.L (L[629:615]),
	.V2C_1 (V2C_42_78),
	.V2C_2 (V2C_42_88),
	.V2C_3 (V2C_42_170),
	.V2C_4 (V2C_42_201),
	.V2C_5 (V2C_42_223),
	.V2C_6 (V2C_42_263),
	.V (V_42)
);

VNU_6 #(quan_width) VNU43 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_84_43),
	.C2V_2 (C2V_94_43),
	.C2V_3 (C2V_176_43),
	.C2V_4 (C2V_207_43),
	.C2V_5 (C2V_229_43),
	.C2V_6 (C2V_269_43),
	.L (L[644:630]),
	.V2C_1 (V2C_43_84),
	.V2C_2 (V2C_43_94),
	.V2C_3 (V2C_43_176),
	.V2C_4 (V2C_43_207),
	.V2C_5 (V2C_43_229),
	.V2C_6 (V2C_43_269),
	.V (V_43)
);

VNU_6 #(quan_width) VNU44 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_90_44),
	.C2V_2 (C2V_100_44),
	.C2V_3 (C2V_182_44),
	.C2V_4 (C2V_213_44),
	.C2V_5 (C2V_235_44),
	.C2V_6 (C2V_275_44),
	.L (L[659:645]),
	.V2C_1 (V2C_44_90),
	.V2C_2 (V2C_44_100),
	.V2C_3 (V2C_44_182),
	.V2C_4 (V2C_44_213),
	.V2C_5 (V2C_44_235),
	.V2C_6 (V2C_44_275),
	.V (V_44)
);

VNU_6 #(quan_width) VNU45 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_96_45),
	.C2V_2 (C2V_106_45),
	.C2V_3 (C2V_188_45),
	.C2V_4 (C2V_219_45),
	.C2V_5 (C2V_241_45),
	.C2V_6 (C2V_281_45),
	.L (L[674:660]),
	.V2C_1 (V2C_45_96),
	.V2C_2 (V2C_45_106),
	.V2C_3 (V2C_45_188),
	.V2C_4 (V2C_45_219),
	.V2C_5 (V2C_45_241),
	.V2C_6 (V2C_45_281),
	.V (V_45)
);

VNU_6 #(quan_width) VNU46 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_102_46),
	.C2V_2 (C2V_112_46),
	.C2V_3 (C2V_194_46),
	.C2V_4 (C2V_225_46),
	.C2V_5 (C2V_247_46),
	.C2V_6 (C2V_287_46),
	.L (L[689:675]),
	.V2C_1 (V2C_46_102),
	.V2C_2 (V2C_46_112),
	.V2C_3 (V2C_46_194),
	.V2C_4 (V2C_46_225),
	.V2C_5 (V2C_46_247),
	.V2C_6 (V2C_46_287),
	.V (V_46)
);

VNU_6 #(quan_width) VNU47 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_47),
	.C2V_2 (C2V_108_47),
	.C2V_3 (C2V_118_47),
	.C2V_4 (C2V_200_47),
	.C2V_5 (C2V_231_47),
	.C2V_6 (C2V_253_47),
	.L (L[704:690]),
	.V2C_1 (V2C_47_5),
	.V2C_2 (V2C_47_108),
	.V2C_3 (V2C_47_118),
	.V2C_4 (V2C_47_200),
	.V2C_5 (V2C_47_231),
	.V2C_6 (V2C_47_253),
	.V (V_47)
);

VNU_6 #(quan_width) VNU48 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_48),
	.C2V_2 (C2V_114_48),
	.C2V_3 (C2V_124_48),
	.C2V_4 (C2V_206_48),
	.C2V_5 (C2V_237_48),
	.C2V_6 (C2V_259_48),
	.L (L[719:705]),
	.V2C_1 (V2C_48_11),
	.V2C_2 (V2C_48_114),
	.V2C_3 (V2C_48_124),
	.V2C_4 (V2C_48_206),
	.V2C_5 (V2C_48_237),
	.V2C_6 (V2C_48_259),
	.V (V_48)
);

VNU_6 #(quan_width) VNU49 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_49),
	.C2V_2 (C2V_64_49),
	.C2V_3 (C2V_81_49),
	.C2V_4 (C2V_206_49),
	.C2V_5 (C2V_245_49),
	.C2V_6 (C2V_264_49),
	.L (L[734:720]),
	.V2C_1 (V2C_49_49),
	.V2C_2 (V2C_49_64),
	.V2C_3 (V2C_49_81),
	.V2C_4 (V2C_49_206),
	.V2C_5 (V2C_49_245),
	.V2C_6 (V2C_49_264),
	.V (V_49)
);

VNU_6 #(quan_width) VNU50 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_50),
	.C2V_2 (C2V_70_50),
	.C2V_3 (C2V_87_50),
	.C2V_4 (C2V_212_50),
	.C2V_5 (C2V_251_50),
	.C2V_6 (C2V_270_50),
	.L (L[749:735]),
	.V2C_1 (V2C_50_55),
	.V2C_2 (V2C_50_70),
	.V2C_3 (V2C_50_87),
	.V2C_4 (V2C_50_212),
	.V2C_5 (V2C_50_251),
	.V2C_6 (V2C_50_270),
	.V (V_50)
);

VNU_6 #(quan_width) VNU51 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_51),
	.C2V_2 (C2V_76_51),
	.C2V_3 (C2V_93_51),
	.C2V_4 (C2V_218_51),
	.C2V_5 (C2V_257_51),
	.C2V_6 (C2V_276_51),
	.L (L[764:750]),
	.V2C_1 (V2C_51_61),
	.V2C_2 (V2C_51_76),
	.V2C_3 (V2C_51_93),
	.V2C_4 (V2C_51_218),
	.V2C_5 (V2C_51_257),
	.V2C_6 (V2C_51_276),
	.V (V_51)
);

VNU_6 #(quan_width) VNU52 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_52),
	.C2V_2 (C2V_82_52),
	.C2V_3 (C2V_99_52),
	.C2V_4 (C2V_224_52),
	.C2V_5 (C2V_263_52),
	.C2V_6 (C2V_282_52),
	.L (L[779:765]),
	.V2C_1 (V2C_52_67),
	.V2C_2 (V2C_52_82),
	.V2C_3 (V2C_52_99),
	.V2C_4 (V2C_52_224),
	.V2C_5 (V2C_52_263),
	.V2C_6 (V2C_52_282),
	.V (V_52)
);

VNU_6 #(quan_width) VNU53 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_53),
	.C2V_2 (C2V_88_53),
	.C2V_3 (C2V_105_53),
	.C2V_4 (C2V_230_53),
	.C2V_5 (C2V_269_53),
	.C2V_6 (C2V_288_53),
	.L (L[794:780]),
	.V2C_1 (V2C_53_73),
	.V2C_2 (V2C_53_88),
	.V2C_3 (V2C_53_105),
	.V2C_4 (V2C_53_230),
	.V2C_5 (V2C_53_269),
	.V2C_6 (V2C_53_288),
	.V (V_53)
);

VNU_6 #(quan_width) VNU54 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_54),
	.C2V_2 (C2V_79_54),
	.C2V_3 (C2V_94_54),
	.C2V_4 (C2V_111_54),
	.C2V_5 (C2V_236_54),
	.C2V_6 (C2V_275_54),
	.L (L[809:795]),
	.V2C_1 (V2C_54_6),
	.V2C_2 (V2C_54_79),
	.V2C_3 (V2C_54_94),
	.V2C_4 (V2C_54_111),
	.V2C_5 (V2C_54_236),
	.V2C_6 (V2C_54_275),
	.V (V_54)
);

VNU_6 #(quan_width) VNU55 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_55),
	.C2V_2 (C2V_85_55),
	.C2V_3 (C2V_100_55),
	.C2V_4 (C2V_117_55),
	.C2V_5 (C2V_242_55),
	.C2V_6 (C2V_281_55),
	.L (L[824:810]),
	.V2C_1 (V2C_55_12),
	.V2C_2 (V2C_55_85),
	.V2C_3 (V2C_55_100),
	.V2C_4 (V2C_55_117),
	.V2C_5 (V2C_55_242),
	.V2C_6 (V2C_55_281),
	.V (V_55)
);

VNU_6 #(quan_width) VNU56 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_56),
	.C2V_2 (C2V_91_56),
	.C2V_3 (C2V_106_56),
	.C2V_4 (C2V_123_56),
	.C2V_5 (C2V_248_56),
	.C2V_6 (C2V_287_56),
	.L (L[839:825]),
	.V2C_1 (V2C_56_18),
	.V2C_2 (V2C_56_91),
	.V2C_3 (V2C_56_106),
	.V2C_4 (V2C_56_123),
	.V2C_5 (V2C_56_248),
	.V2C_6 (V2C_56_287),
	.V (V_56)
);

VNU_6 #(quan_width) VNU57 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_57),
	.C2V_2 (C2V_24_57),
	.C2V_3 (C2V_97_57),
	.C2V_4 (C2V_112_57),
	.C2V_5 (C2V_129_57),
	.C2V_6 (C2V_254_57),
	.L (L[854:840]),
	.V2C_1 (V2C_57_5),
	.V2C_2 (V2C_57_24),
	.V2C_3 (V2C_57_97),
	.V2C_4 (V2C_57_112),
	.V2C_5 (V2C_57_129),
	.V2C_6 (V2C_57_254),
	.V (V_57)
);

VNU_6 #(quan_width) VNU58 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_58),
	.C2V_2 (C2V_30_58),
	.C2V_3 (C2V_103_58),
	.C2V_4 (C2V_118_58),
	.C2V_5 (C2V_135_58),
	.C2V_6 (C2V_260_58),
	.L (L[869:855]),
	.V2C_1 (V2C_58_11),
	.V2C_2 (V2C_58_30),
	.V2C_3 (V2C_58_103),
	.V2C_4 (V2C_58_118),
	.V2C_5 (V2C_58_135),
	.V2C_6 (V2C_58_260),
	.V (V_58)
);

VNU_6 #(quan_width) VNU59 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_59),
	.C2V_2 (C2V_36_59),
	.C2V_3 (C2V_109_59),
	.C2V_4 (C2V_124_59),
	.C2V_5 (C2V_141_59),
	.C2V_6 (C2V_266_59),
	.L (L[884:870]),
	.V2C_1 (V2C_59_17),
	.V2C_2 (V2C_59_36),
	.V2C_3 (V2C_59_109),
	.V2C_4 (V2C_59_124),
	.V2C_5 (V2C_59_141),
	.V2C_6 (V2C_59_266),
	.V (V_59)
);

VNU_6 #(quan_width) VNU60 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_60),
	.C2V_2 (C2V_42_60),
	.C2V_3 (C2V_115_60),
	.C2V_4 (C2V_130_60),
	.C2V_5 (C2V_147_60),
	.C2V_6 (C2V_272_60),
	.L (L[899:885]),
	.V2C_1 (V2C_60_23),
	.V2C_2 (V2C_60_42),
	.V2C_3 (V2C_60_115),
	.V2C_4 (V2C_60_130),
	.V2C_5 (V2C_60_147),
	.V2C_6 (V2C_60_272),
	.V (V_60)
);

VNU_6 #(quan_width) VNU61 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_61),
	.C2V_2 (C2V_48_61),
	.C2V_3 (C2V_121_61),
	.C2V_4 (C2V_136_61),
	.C2V_5 (C2V_153_61),
	.C2V_6 (C2V_278_61),
	.L (L[914:900]),
	.V2C_1 (V2C_61_29),
	.V2C_2 (V2C_61_48),
	.V2C_3 (V2C_61_121),
	.V2C_4 (V2C_61_136),
	.V2C_5 (V2C_61_153),
	.V2C_6 (V2C_61_278),
	.V (V_61)
);

VNU_6 #(quan_width) VNU62 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_62),
	.C2V_2 (C2V_54_62),
	.C2V_3 (C2V_127_62),
	.C2V_4 (C2V_142_62),
	.C2V_5 (C2V_159_62),
	.C2V_6 (C2V_284_62),
	.L (L[929:915]),
	.V2C_1 (V2C_62_35),
	.V2C_2 (V2C_62_54),
	.V2C_3 (V2C_62_127),
	.V2C_4 (V2C_62_142),
	.V2C_5 (V2C_62_159),
	.V2C_6 (V2C_62_284),
	.V (V_62)
);

VNU_6 #(quan_width) VNU63 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_63),
	.C2V_2 (C2V_41_63),
	.C2V_3 (C2V_60_63),
	.C2V_4 (C2V_133_63),
	.C2V_5 (C2V_148_63),
	.C2V_6 (C2V_165_63),
	.L (L[944:930]),
	.V2C_1 (V2C_63_2),
	.V2C_2 (V2C_63_41),
	.V2C_3 (V2C_63_60),
	.V2C_4 (V2C_63_133),
	.V2C_5 (V2C_63_148),
	.V2C_6 (V2C_63_165),
	.V (V_63)
);

VNU_6 #(quan_width) VNU64 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_64),
	.C2V_2 (C2V_47_64),
	.C2V_3 (C2V_66_64),
	.C2V_4 (C2V_139_64),
	.C2V_5 (C2V_154_64),
	.C2V_6 (C2V_171_64),
	.L (L[959:945]),
	.V2C_1 (V2C_64_8),
	.V2C_2 (V2C_64_47),
	.V2C_3 (V2C_64_66),
	.V2C_4 (V2C_64_139),
	.V2C_5 (V2C_64_154),
	.V2C_6 (V2C_64_171),
	.V (V_64)
);

VNU_6 #(quan_width) VNU65 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_65),
	.C2V_2 (C2V_53_65),
	.C2V_3 (C2V_72_65),
	.C2V_4 (C2V_145_65),
	.C2V_5 (C2V_160_65),
	.C2V_6 (C2V_177_65),
	.L (L[974:960]),
	.V2C_1 (V2C_65_14),
	.V2C_2 (V2C_65_53),
	.V2C_3 (V2C_65_72),
	.V2C_4 (V2C_65_145),
	.V2C_5 (V2C_65_160),
	.V2C_6 (V2C_65_177),
	.V (V_65)
);

VNU_6 #(quan_width) VNU66 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_66),
	.C2V_2 (C2V_59_66),
	.C2V_3 (C2V_78_66),
	.C2V_4 (C2V_151_66),
	.C2V_5 (C2V_166_66),
	.C2V_6 (C2V_183_66),
	.L (L[989:975]),
	.V2C_1 (V2C_66_20),
	.V2C_2 (V2C_66_59),
	.V2C_3 (V2C_66_78),
	.V2C_4 (V2C_66_151),
	.V2C_5 (V2C_66_166),
	.V2C_6 (V2C_66_183),
	.V (V_66)
);

VNU_6 #(quan_width) VNU67 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_67),
	.C2V_2 (C2V_65_67),
	.C2V_3 (C2V_84_67),
	.C2V_4 (C2V_157_67),
	.C2V_5 (C2V_172_67),
	.C2V_6 (C2V_189_67),
	.L (L[1004:990]),
	.V2C_1 (V2C_67_26),
	.V2C_2 (V2C_67_65),
	.V2C_3 (V2C_67_84),
	.V2C_4 (V2C_67_157),
	.V2C_5 (V2C_67_172),
	.V2C_6 (V2C_67_189),
	.V (V_67)
);

VNU_6 #(quan_width) VNU68 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_68),
	.C2V_2 (C2V_71_68),
	.C2V_3 (C2V_90_68),
	.C2V_4 (C2V_163_68),
	.C2V_5 (C2V_178_68),
	.C2V_6 (C2V_195_68),
	.L (L[1019:1005]),
	.V2C_1 (V2C_68_32),
	.V2C_2 (V2C_68_71),
	.V2C_3 (V2C_68_90),
	.V2C_4 (V2C_68_163),
	.V2C_5 (V2C_68_178),
	.V2C_6 (V2C_68_195),
	.V (V_68)
);

VNU_6 #(quan_width) VNU69 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_69),
	.C2V_2 (C2V_77_69),
	.C2V_3 (C2V_96_69),
	.C2V_4 (C2V_169_69),
	.C2V_5 (C2V_184_69),
	.C2V_6 (C2V_201_69),
	.L (L[1034:1020]),
	.V2C_1 (V2C_69_38),
	.V2C_2 (V2C_69_77),
	.V2C_3 (V2C_69_96),
	.V2C_4 (V2C_69_169),
	.V2C_5 (V2C_69_184),
	.V2C_6 (V2C_69_201),
	.V (V_69)
);

VNU_6 #(quan_width) VNU70 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_70),
	.C2V_2 (C2V_83_70),
	.C2V_3 (C2V_102_70),
	.C2V_4 (C2V_175_70),
	.C2V_5 (C2V_190_70),
	.C2V_6 (C2V_207_70),
	.L (L[1049:1035]),
	.V2C_1 (V2C_70_44),
	.V2C_2 (V2C_70_83),
	.V2C_3 (V2C_70_102),
	.V2C_4 (V2C_70_175),
	.V2C_5 (V2C_70_190),
	.V2C_6 (V2C_70_207),
	.V (V_70)
);

VNU_6 #(quan_width) VNU71 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_71),
	.C2V_2 (C2V_89_71),
	.C2V_3 (C2V_108_71),
	.C2V_4 (C2V_181_71),
	.C2V_5 (C2V_196_71),
	.C2V_6 (C2V_213_71),
	.L (L[1064:1050]),
	.V2C_1 (V2C_71_50),
	.V2C_2 (V2C_71_89),
	.V2C_3 (V2C_71_108),
	.V2C_4 (V2C_71_181),
	.V2C_5 (V2C_71_196),
	.V2C_6 (V2C_71_213),
	.V (V_71)
);

VNU_6 #(quan_width) VNU72 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_72),
	.C2V_2 (C2V_95_72),
	.C2V_3 (C2V_114_72),
	.C2V_4 (C2V_187_72),
	.C2V_5 (C2V_202_72),
	.C2V_6 (C2V_219_72),
	.L (L[1079:1065]),
	.V2C_1 (V2C_72_56),
	.V2C_2 (V2C_72_95),
	.V2C_3 (V2C_72_114),
	.V2C_4 (V2C_72_187),
	.V2C_5 (V2C_72_202),
	.V2C_6 (V2C_72_219),
	.V (V_72)
);

VNU_6 #(quan_width) VNU73 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_73),
	.C2V_2 (C2V_101_73),
	.C2V_3 (C2V_120_73),
	.C2V_4 (C2V_193_73),
	.C2V_5 (C2V_208_73),
	.C2V_6 (C2V_225_73),
	.L (L[1094:1080]),
	.V2C_1 (V2C_73_62),
	.V2C_2 (V2C_73_101),
	.V2C_3 (V2C_73_120),
	.V2C_4 (V2C_73_193),
	.V2C_5 (V2C_73_208),
	.V2C_6 (V2C_73_225),
	.V (V_73)
);

VNU_6 #(quan_width) VNU74 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_74),
	.C2V_2 (C2V_107_74),
	.C2V_3 (C2V_126_74),
	.C2V_4 (C2V_199_74),
	.C2V_5 (C2V_214_74),
	.C2V_6 (C2V_231_74),
	.L (L[1109:1095]),
	.V2C_1 (V2C_74_68),
	.V2C_2 (V2C_74_107),
	.V2C_3 (V2C_74_126),
	.V2C_4 (V2C_74_199),
	.V2C_5 (V2C_74_214),
	.V2C_6 (V2C_74_231),
	.V (V_74)
);

VNU_6 #(quan_width) VNU75 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_75),
	.C2V_2 (C2V_113_75),
	.C2V_3 (C2V_132_75),
	.C2V_4 (C2V_205_75),
	.C2V_5 (C2V_220_75),
	.C2V_6 (C2V_237_75),
	.L (L[1124:1110]),
	.V2C_1 (V2C_75_74),
	.V2C_2 (V2C_75_113),
	.V2C_3 (V2C_75_132),
	.V2C_4 (V2C_75_205),
	.V2C_5 (V2C_75_220),
	.V2C_6 (V2C_75_237),
	.V (V_75)
);

VNU_6 #(quan_width) VNU76 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_80_76),
	.C2V_2 (C2V_119_76),
	.C2V_3 (C2V_138_76),
	.C2V_4 (C2V_211_76),
	.C2V_5 (C2V_226_76),
	.C2V_6 (C2V_243_76),
	.L (L[1139:1125]),
	.V2C_1 (V2C_76_80),
	.V2C_2 (V2C_76_119),
	.V2C_3 (V2C_76_138),
	.V2C_4 (V2C_76_211),
	.V2C_5 (V2C_76_226),
	.V2C_6 (V2C_76_243),
	.V (V_76)
);

VNU_6 #(quan_width) VNU77 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_86_77),
	.C2V_2 (C2V_125_77),
	.C2V_3 (C2V_144_77),
	.C2V_4 (C2V_217_77),
	.C2V_5 (C2V_232_77),
	.C2V_6 (C2V_249_77),
	.L (L[1154:1140]),
	.V2C_1 (V2C_77_86),
	.V2C_2 (V2C_77_125),
	.V2C_3 (V2C_77_144),
	.V2C_4 (V2C_77_217),
	.V2C_5 (V2C_77_232),
	.V2C_6 (V2C_77_249),
	.V (V_77)
);

VNU_6 #(quan_width) VNU78 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_92_78),
	.C2V_2 (C2V_131_78),
	.C2V_3 (C2V_150_78),
	.C2V_4 (C2V_223_78),
	.C2V_5 (C2V_238_78),
	.C2V_6 (C2V_255_78),
	.L (L[1169:1155]),
	.V2C_1 (V2C_78_92),
	.V2C_2 (V2C_78_131),
	.V2C_3 (V2C_78_150),
	.V2C_4 (V2C_78_223),
	.V2C_5 (V2C_78_238),
	.V2C_6 (V2C_78_255),
	.V (V_78)
);

VNU_6 #(quan_width) VNU79 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_98_79),
	.C2V_2 (C2V_137_79),
	.C2V_3 (C2V_156_79),
	.C2V_4 (C2V_229_79),
	.C2V_5 (C2V_244_79),
	.C2V_6 (C2V_261_79),
	.L (L[1184:1170]),
	.V2C_1 (V2C_79_98),
	.V2C_2 (V2C_79_137),
	.V2C_3 (V2C_79_156),
	.V2C_4 (V2C_79_229),
	.V2C_5 (V2C_79_244),
	.V2C_6 (V2C_79_261),
	.V (V_79)
);

VNU_6 #(quan_width) VNU80 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_104_80),
	.C2V_2 (C2V_143_80),
	.C2V_3 (C2V_162_80),
	.C2V_4 (C2V_235_80),
	.C2V_5 (C2V_250_80),
	.C2V_6 (C2V_267_80),
	.L (L[1199:1185]),
	.V2C_1 (V2C_80_104),
	.V2C_2 (V2C_80_143),
	.V2C_3 (V2C_80_162),
	.V2C_4 (V2C_80_235),
	.V2C_5 (V2C_80_250),
	.V2C_6 (V2C_80_267),
	.V (V_80)
);

VNU_6 #(quan_width) VNU81 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_110_81),
	.C2V_2 (C2V_149_81),
	.C2V_3 (C2V_168_81),
	.C2V_4 (C2V_241_81),
	.C2V_5 (C2V_256_81),
	.C2V_6 (C2V_273_81),
	.L (L[1214:1200]),
	.V2C_1 (V2C_81_110),
	.V2C_2 (V2C_81_149),
	.V2C_3 (V2C_81_168),
	.V2C_4 (V2C_81_241),
	.V2C_5 (V2C_81_256),
	.V2C_6 (V2C_81_273),
	.V (V_81)
);

VNU_6 #(quan_width) VNU82 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_116_82),
	.C2V_2 (C2V_155_82),
	.C2V_3 (C2V_174_82),
	.C2V_4 (C2V_247_82),
	.C2V_5 (C2V_262_82),
	.C2V_6 (C2V_279_82),
	.L (L[1229:1215]),
	.V2C_1 (V2C_82_116),
	.V2C_2 (V2C_82_155),
	.V2C_3 (V2C_82_174),
	.V2C_4 (V2C_82_247),
	.V2C_5 (V2C_82_262),
	.V2C_6 (V2C_82_279),
	.V (V_82)
);

VNU_6 #(quan_width) VNU83 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_122_83),
	.C2V_2 (C2V_161_83),
	.C2V_3 (C2V_180_83),
	.C2V_4 (C2V_253_83),
	.C2V_5 (C2V_268_83),
	.C2V_6 (C2V_285_83),
	.L (L[1244:1230]),
	.V2C_1 (V2C_83_122),
	.V2C_2 (V2C_83_161),
	.V2C_3 (V2C_83_180),
	.V2C_4 (V2C_83_253),
	.V2C_5 (V2C_83_268),
	.V2C_6 (V2C_83_285),
	.V (V_83)
);

VNU_6 #(quan_width) VNU84 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_84),
	.C2V_2 (C2V_128_84),
	.C2V_3 (C2V_167_84),
	.C2V_4 (C2V_186_84),
	.C2V_5 (C2V_259_84),
	.C2V_6 (C2V_274_84),
	.L (L[1259:1245]),
	.V2C_1 (V2C_84_3),
	.V2C_2 (V2C_84_128),
	.V2C_3 (V2C_84_167),
	.V2C_4 (V2C_84_186),
	.V2C_5 (V2C_84_259),
	.V2C_6 (V2C_84_274),
	.V (V_84)
);

VNU_6 #(quan_width) VNU85 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_85),
	.C2V_2 (C2V_134_85),
	.C2V_3 (C2V_173_85),
	.C2V_4 (C2V_192_85),
	.C2V_5 (C2V_265_85),
	.C2V_6 (C2V_280_85),
	.L (L[1274:1260]),
	.V2C_1 (V2C_85_9),
	.V2C_2 (V2C_85_134),
	.V2C_3 (V2C_85_173),
	.V2C_4 (V2C_85_192),
	.V2C_5 (V2C_85_265),
	.V2C_6 (V2C_85_280),
	.V (V_85)
);

VNU_6 #(quan_width) VNU86 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_86),
	.C2V_2 (C2V_140_86),
	.C2V_3 (C2V_179_86),
	.C2V_4 (C2V_198_86),
	.C2V_5 (C2V_271_86),
	.C2V_6 (C2V_286_86),
	.L (L[1289:1275]),
	.V2C_1 (V2C_86_15),
	.V2C_2 (V2C_86_140),
	.V2C_3 (V2C_86_179),
	.V2C_4 (V2C_86_198),
	.V2C_5 (V2C_86_271),
	.V2C_6 (V2C_86_286),
	.V (V_86)
);

VNU_6 #(quan_width) VNU87 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_87),
	.C2V_2 (C2V_21_87),
	.C2V_3 (C2V_146_87),
	.C2V_4 (C2V_185_87),
	.C2V_5 (C2V_204_87),
	.C2V_6 (C2V_277_87),
	.L (L[1304:1290]),
	.V2C_1 (V2C_87_4),
	.V2C_2 (V2C_87_21),
	.V2C_3 (V2C_87_146),
	.V2C_4 (V2C_87_185),
	.V2C_5 (V2C_87_204),
	.V2C_6 (V2C_87_277),
	.V (V_87)
);

VNU_6 #(quan_width) VNU88 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_88),
	.C2V_2 (C2V_27_88),
	.C2V_3 (C2V_152_88),
	.C2V_4 (C2V_191_88),
	.C2V_5 (C2V_210_88),
	.C2V_6 (C2V_283_88),
	.L (L[1319:1305]),
	.V2C_1 (V2C_88_10),
	.V2C_2 (V2C_88_27),
	.V2C_3 (V2C_88_152),
	.V2C_4 (V2C_88_191),
	.V2C_5 (V2C_88_210),
	.V2C_6 (V2C_88_283),
	.V (V_88)
);

VNU_6 #(quan_width) VNU89 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_89),
	.C2V_2 (C2V_16_89),
	.C2V_3 (C2V_33_89),
	.C2V_4 (C2V_158_89),
	.C2V_5 (C2V_197_89),
	.C2V_6 (C2V_216_89),
	.L (L[1334:1320]),
	.V2C_1 (V2C_89_1),
	.V2C_2 (V2C_89_16),
	.V2C_3 (V2C_89_33),
	.V2C_4 (V2C_89_158),
	.V2C_5 (V2C_89_197),
	.V2C_6 (V2C_89_216),
	.V (V_89)
);

VNU_6 #(quan_width) VNU90 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_90),
	.C2V_2 (C2V_22_90),
	.C2V_3 (C2V_39_90),
	.C2V_4 (C2V_164_90),
	.C2V_5 (C2V_203_90),
	.C2V_6 (C2V_222_90),
	.L (L[1349:1335]),
	.V2C_1 (V2C_90_7),
	.V2C_2 (V2C_90_22),
	.V2C_3 (V2C_90_39),
	.V2C_4 (V2C_90_164),
	.V2C_5 (V2C_90_203),
	.V2C_6 (V2C_90_222),
	.V (V_90)
);

VNU_6 #(quan_width) VNU91 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_91),
	.C2V_2 (C2V_28_91),
	.C2V_3 (C2V_45_91),
	.C2V_4 (C2V_170_91),
	.C2V_5 (C2V_209_91),
	.C2V_6 (C2V_228_91),
	.L (L[1364:1350]),
	.V2C_1 (V2C_91_13),
	.V2C_2 (V2C_91_28),
	.V2C_3 (V2C_91_45),
	.V2C_4 (V2C_91_170),
	.V2C_5 (V2C_91_209),
	.V2C_6 (V2C_91_228),
	.V (V_91)
);

VNU_6 #(quan_width) VNU92 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_92),
	.C2V_2 (C2V_34_92),
	.C2V_3 (C2V_51_92),
	.C2V_4 (C2V_176_92),
	.C2V_5 (C2V_215_92),
	.C2V_6 (C2V_234_92),
	.L (L[1379:1365]),
	.V2C_1 (V2C_92_19),
	.V2C_2 (V2C_92_34),
	.V2C_3 (V2C_92_51),
	.V2C_4 (V2C_92_176),
	.V2C_5 (V2C_92_215),
	.V2C_6 (V2C_92_234),
	.V (V_92)
);

VNU_6 #(quan_width) VNU93 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_93),
	.C2V_2 (C2V_40_93),
	.C2V_3 (C2V_57_93),
	.C2V_4 (C2V_182_93),
	.C2V_5 (C2V_221_93),
	.C2V_6 (C2V_240_93),
	.L (L[1394:1380]),
	.V2C_1 (V2C_93_25),
	.V2C_2 (V2C_93_40),
	.V2C_3 (V2C_93_57),
	.V2C_4 (V2C_93_182),
	.V2C_5 (V2C_93_221),
	.V2C_6 (V2C_93_240),
	.V (V_93)
);

VNU_6 #(quan_width) VNU94 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_94),
	.C2V_2 (C2V_46_94),
	.C2V_3 (C2V_63_94),
	.C2V_4 (C2V_188_94),
	.C2V_5 (C2V_227_94),
	.C2V_6 (C2V_246_94),
	.L (L[1409:1395]),
	.V2C_1 (V2C_94_31),
	.V2C_2 (V2C_94_46),
	.V2C_3 (V2C_94_63),
	.V2C_4 (V2C_94_188),
	.V2C_5 (V2C_94_227),
	.V2C_6 (V2C_94_246),
	.V (V_94)
);

VNU_6 #(quan_width) VNU95 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_95),
	.C2V_2 (C2V_52_95),
	.C2V_3 (C2V_69_95),
	.C2V_4 (C2V_194_95),
	.C2V_5 (C2V_233_95),
	.C2V_6 (C2V_252_95),
	.L (L[1424:1410]),
	.V2C_1 (V2C_95_37),
	.V2C_2 (V2C_95_52),
	.V2C_3 (V2C_95_69),
	.V2C_4 (V2C_95_194),
	.V2C_5 (V2C_95_233),
	.V2C_6 (V2C_95_252),
	.V (V_95)
);

VNU_6 #(quan_width) VNU96 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_96),
	.C2V_2 (C2V_58_96),
	.C2V_3 (C2V_75_96),
	.C2V_4 (C2V_200_96),
	.C2V_5 (C2V_239_96),
	.C2V_6 (C2V_258_96),
	.L (L[1439:1425]),
	.V2C_1 (V2C_96_43),
	.V2C_2 (V2C_96_58),
	.V2C_3 (V2C_96_75),
	.V2C_4 (V2C_96_200),
	.V2C_5 (V2C_96_239),
	.V2C_6 (V2C_96_258),
	.V (V_96)
);

VNU_6 #(quan_width) VNU97 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_97),
	.C2V_2 (C2V_35_97),
	.C2V_3 (C2V_118_97),
	.C2V_4 (C2V_158_97),
	.C2V_5 (C2V_217_97),
	.C2V_6 (C2V_267_97),
	.L (L[1454:1440]),
	.V2C_1 (V2C_97_24),
	.V2C_2 (V2C_97_35),
	.V2C_3 (V2C_97_118),
	.V2C_4 (V2C_97_158),
	.V2C_5 (V2C_97_217),
	.V2C_6 (V2C_97_267),
	.V (V_97)
);

VNU_6 #(quan_width) VNU98 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_98),
	.C2V_2 (C2V_41_98),
	.C2V_3 (C2V_124_98),
	.C2V_4 (C2V_164_98),
	.C2V_5 (C2V_223_98),
	.C2V_6 (C2V_273_98),
	.L (L[1469:1455]),
	.V2C_1 (V2C_98_30),
	.V2C_2 (V2C_98_41),
	.V2C_3 (V2C_98_124),
	.V2C_4 (V2C_98_164),
	.V2C_5 (V2C_98_223),
	.V2C_6 (V2C_98_273),
	.V (V_98)
);

VNU_6 #(quan_width) VNU99 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_99),
	.C2V_2 (C2V_47_99),
	.C2V_3 (C2V_130_99),
	.C2V_4 (C2V_170_99),
	.C2V_5 (C2V_229_99),
	.C2V_6 (C2V_279_99),
	.L (L[1484:1470]),
	.V2C_1 (V2C_99_36),
	.V2C_2 (V2C_99_47),
	.V2C_3 (V2C_99_130),
	.V2C_4 (V2C_99_170),
	.V2C_5 (V2C_99_229),
	.V2C_6 (V2C_99_279),
	.V (V_99)
);

VNU_6 #(quan_width) VNU100 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_100),
	.C2V_2 (C2V_53_100),
	.C2V_3 (C2V_136_100),
	.C2V_4 (C2V_176_100),
	.C2V_5 (C2V_235_100),
	.C2V_6 (C2V_285_100),
	.L (L[1499:1485]),
	.V2C_1 (V2C_100_42),
	.V2C_2 (V2C_100_53),
	.V2C_3 (V2C_100_136),
	.V2C_4 (V2C_100_176),
	.V2C_5 (V2C_100_235),
	.V2C_6 (V2C_100_285),
	.V (V_100)
);

VNU_6 #(quan_width) VNU101 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_101),
	.C2V_2 (C2V_48_101),
	.C2V_3 (C2V_59_101),
	.C2V_4 (C2V_142_101),
	.C2V_5 (C2V_182_101),
	.C2V_6 (C2V_241_101),
	.L (L[1514:1500]),
	.V2C_1 (V2C_101_3),
	.V2C_2 (V2C_101_48),
	.V2C_3 (V2C_101_59),
	.V2C_4 (V2C_101_142),
	.V2C_5 (V2C_101_182),
	.V2C_6 (V2C_101_241),
	.V (V_101)
);

VNU_6 #(quan_width) VNU102 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_102),
	.C2V_2 (C2V_54_102),
	.C2V_3 (C2V_65_102),
	.C2V_4 (C2V_148_102),
	.C2V_5 (C2V_188_102),
	.C2V_6 (C2V_247_102),
	.L (L[1529:1515]),
	.V2C_1 (V2C_102_9),
	.V2C_2 (V2C_102_54),
	.V2C_3 (V2C_102_65),
	.V2C_4 (V2C_102_148),
	.V2C_5 (V2C_102_188),
	.V2C_6 (V2C_102_247),
	.V (V_102)
);

VNU_6 #(quan_width) VNU103 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_103),
	.C2V_2 (C2V_60_103),
	.C2V_3 (C2V_71_103),
	.C2V_4 (C2V_154_103),
	.C2V_5 (C2V_194_103),
	.C2V_6 (C2V_253_103),
	.L (L[1544:1530]),
	.V2C_1 (V2C_103_15),
	.V2C_2 (V2C_103_60),
	.V2C_3 (V2C_103_71),
	.V2C_4 (V2C_103_154),
	.V2C_5 (V2C_103_194),
	.V2C_6 (V2C_103_253),
	.V (V_103)
);

VNU_6 #(quan_width) VNU104 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_104),
	.C2V_2 (C2V_66_104),
	.C2V_3 (C2V_77_104),
	.C2V_4 (C2V_160_104),
	.C2V_5 (C2V_200_104),
	.C2V_6 (C2V_259_104),
	.L (L[1559:1545]),
	.V2C_1 (V2C_104_21),
	.V2C_2 (V2C_104_66),
	.V2C_3 (V2C_104_77),
	.V2C_4 (V2C_104_160),
	.V2C_5 (V2C_104_200),
	.V2C_6 (V2C_104_259),
	.V (V_104)
);

VNU_6 #(quan_width) VNU105 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_105),
	.C2V_2 (C2V_72_105),
	.C2V_3 (C2V_83_105),
	.C2V_4 (C2V_166_105),
	.C2V_5 (C2V_206_105),
	.C2V_6 (C2V_265_105),
	.L (L[1574:1560]),
	.V2C_1 (V2C_105_27),
	.V2C_2 (V2C_105_72),
	.V2C_3 (V2C_105_83),
	.V2C_4 (V2C_105_166),
	.V2C_5 (V2C_105_206),
	.V2C_6 (V2C_105_265),
	.V (V_105)
);

VNU_6 #(quan_width) VNU106 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_106),
	.C2V_2 (C2V_78_106),
	.C2V_3 (C2V_89_106),
	.C2V_4 (C2V_172_106),
	.C2V_5 (C2V_212_106),
	.C2V_6 (C2V_271_106),
	.L (L[1589:1575]),
	.V2C_1 (V2C_106_33),
	.V2C_2 (V2C_106_78),
	.V2C_3 (V2C_106_89),
	.V2C_4 (V2C_106_172),
	.V2C_5 (V2C_106_212),
	.V2C_6 (V2C_106_271),
	.V (V_106)
);

VNU_6 #(quan_width) VNU107 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_107),
	.C2V_2 (C2V_84_107),
	.C2V_3 (C2V_95_107),
	.C2V_4 (C2V_178_107),
	.C2V_5 (C2V_218_107),
	.C2V_6 (C2V_277_107),
	.L (L[1604:1590]),
	.V2C_1 (V2C_107_39),
	.V2C_2 (V2C_107_84),
	.V2C_3 (V2C_107_95),
	.V2C_4 (V2C_107_178),
	.V2C_5 (V2C_107_218),
	.V2C_6 (V2C_107_277),
	.V (V_107)
);

VNU_6 #(quan_width) VNU108 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_108),
	.C2V_2 (C2V_90_108),
	.C2V_3 (C2V_101_108),
	.C2V_4 (C2V_184_108),
	.C2V_5 (C2V_224_108),
	.C2V_6 (C2V_283_108),
	.L (L[1619:1605]),
	.V2C_1 (V2C_108_45),
	.V2C_2 (V2C_108_90),
	.V2C_3 (V2C_108_101),
	.V2C_4 (V2C_108_184),
	.V2C_5 (V2C_108_224),
	.V2C_6 (V2C_108_283),
	.V (V_108)
);

VNU_6 #(quan_width) VNU109 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_109),
	.C2V_2 (C2V_51_109),
	.C2V_3 (C2V_96_109),
	.C2V_4 (C2V_107_109),
	.C2V_5 (C2V_190_109),
	.C2V_6 (C2V_230_109),
	.L (L[1634:1620]),
	.V2C_1 (V2C_109_1),
	.V2C_2 (V2C_109_51),
	.V2C_3 (V2C_109_96),
	.V2C_4 (V2C_109_107),
	.V2C_5 (V2C_109_190),
	.V2C_6 (V2C_109_230),
	.V (V_109)
);

VNU_6 #(quan_width) VNU110 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_110),
	.C2V_2 (C2V_57_110),
	.C2V_3 (C2V_102_110),
	.C2V_4 (C2V_113_110),
	.C2V_5 (C2V_196_110),
	.C2V_6 (C2V_236_110),
	.L (L[1649:1635]),
	.V2C_1 (V2C_110_7),
	.V2C_2 (V2C_110_57),
	.V2C_3 (V2C_110_102),
	.V2C_4 (V2C_110_113),
	.V2C_5 (V2C_110_196),
	.V2C_6 (V2C_110_236),
	.V (V_110)
);

VNU_6 #(quan_width) VNU111 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_111),
	.C2V_2 (C2V_63_111),
	.C2V_3 (C2V_108_111),
	.C2V_4 (C2V_119_111),
	.C2V_5 (C2V_202_111),
	.C2V_6 (C2V_242_111),
	.L (L[1664:1650]),
	.V2C_1 (V2C_111_13),
	.V2C_2 (V2C_111_63),
	.V2C_3 (V2C_111_108),
	.V2C_4 (V2C_111_119),
	.V2C_5 (V2C_111_202),
	.V2C_6 (V2C_111_242),
	.V (V_111)
);

VNU_6 #(quan_width) VNU112 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_112),
	.C2V_2 (C2V_69_112),
	.C2V_3 (C2V_114_112),
	.C2V_4 (C2V_125_112),
	.C2V_5 (C2V_208_112),
	.C2V_6 (C2V_248_112),
	.L (L[1679:1665]),
	.V2C_1 (V2C_112_19),
	.V2C_2 (V2C_112_69),
	.V2C_3 (V2C_112_114),
	.V2C_4 (V2C_112_125),
	.V2C_5 (V2C_112_208),
	.V2C_6 (V2C_112_248),
	.V (V_112)
);

VNU_6 #(quan_width) VNU113 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_113),
	.C2V_2 (C2V_75_113),
	.C2V_3 (C2V_120_113),
	.C2V_4 (C2V_131_113),
	.C2V_5 (C2V_214_113),
	.C2V_6 (C2V_254_113),
	.L (L[1694:1680]),
	.V2C_1 (V2C_113_25),
	.V2C_2 (V2C_113_75),
	.V2C_3 (V2C_113_120),
	.V2C_4 (V2C_113_131),
	.V2C_5 (V2C_113_214),
	.V2C_6 (V2C_113_254),
	.V (V_113)
);

VNU_6 #(quan_width) VNU114 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_114),
	.C2V_2 (C2V_81_114),
	.C2V_3 (C2V_126_114),
	.C2V_4 (C2V_137_114),
	.C2V_5 (C2V_220_114),
	.C2V_6 (C2V_260_114),
	.L (L[1709:1695]),
	.V2C_1 (V2C_114_31),
	.V2C_2 (V2C_114_81),
	.V2C_3 (V2C_114_126),
	.V2C_4 (V2C_114_137),
	.V2C_5 (V2C_114_220),
	.V2C_6 (V2C_114_260),
	.V (V_114)
);

VNU_6 #(quan_width) VNU115 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_115),
	.C2V_2 (C2V_87_115),
	.C2V_3 (C2V_132_115),
	.C2V_4 (C2V_143_115),
	.C2V_5 (C2V_226_115),
	.C2V_6 (C2V_266_115),
	.L (L[1724:1710]),
	.V2C_1 (V2C_115_37),
	.V2C_2 (V2C_115_87),
	.V2C_3 (V2C_115_132),
	.V2C_4 (V2C_115_143),
	.V2C_5 (V2C_115_226),
	.V2C_6 (V2C_115_266),
	.V (V_115)
);

VNU_6 #(quan_width) VNU116 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_116),
	.C2V_2 (C2V_93_116),
	.C2V_3 (C2V_138_116),
	.C2V_4 (C2V_149_116),
	.C2V_5 (C2V_232_116),
	.C2V_6 (C2V_272_116),
	.L (L[1739:1725]),
	.V2C_1 (V2C_116_43),
	.V2C_2 (V2C_116_93),
	.V2C_3 (V2C_116_138),
	.V2C_4 (V2C_116_149),
	.V2C_5 (V2C_116_232),
	.V2C_6 (V2C_116_272),
	.V (V_116)
);

VNU_6 #(quan_width) VNU117 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_117),
	.C2V_2 (C2V_99_117),
	.C2V_3 (C2V_144_117),
	.C2V_4 (C2V_155_117),
	.C2V_5 (C2V_238_117),
	.C2V_6 (C2V_278_117),
	.L (L[1754:1740]),
	.V2C_1 (V2C_117_49),
	.V2C_2 (V2C_117_99),
	.V2C_3 (V2C_117_144),
	.V2C_4 (V2C_117_155),
	.V2C_5 (V2C_117_238),
	.V2C_6 (V2C_117_278),
	.V (V_117)
);

VNU_6 #(quan_width) VNU118 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_118),
	.C2V_2 (C2V_105_118),
	.C2V_3 (C2V_150_118),
	.C2V_4 (C2V_161_118),
	.C2V_5 (C2V_244_118),
	.C2V_6 (C2V_284_118),
	.L (L[1769:1755]),
	.V2C_1 (V2C_118_55),
	.V2C_2 (V2C_118_105),
	.V2C_3 (V2C_118_150),
	.V2C_4 (V2C_118_161),
	.V2C_5 (V2C_118_244),
	.V2C_6 (V2C_118_284),
	.V (V_118)
);

VNU_6 #(quan_width) VNU119 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_119),
	.C2V_2 (C2V_61_119),
	.C2V_3 (C2V_111_119),
	.C2V_4 (C2V_156_119),
	.C2V_5 (C2V_167_119),
	.C2V_6 (C2V_250_119),
	.L (L[1784:1770]),
	.V2C_1 (V2C_119_2),
	.V2C_2 (V2C_119_61),
	.V2C_3 (V2C_119_111),
	.V2C_4 (V2C_119_156),
	.V2C_5 (V2C_119_167),
	.V2C_6 (V2C_119_250),
	.V (V_119)
);

VNU_6 #(quan_width) VNU120 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_120),
	.C2V_2 (C2V_67_120),
	.C2V_3 (C2V_117_120),
	.C2V_4 (C2V_162_120),
	.C2V_5 (C2V_173_120),
	.C2V_6 (C2V_256_120),
	.L (L[1799:1785]),
	.V2C_1 (V2C_120_8),
	.V2C_2 (V2C_120_67),
	.V2C_3 (V2C_120_117),
	.V2C_4 (V2C_120_162),
	.V2C_5 (V2C_120_173),
	.V2C_6 (V2C_120_256),
	.V (V_120)
);

VNU_6 #(quan_width) VNU121 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_121),
	.C2V_2 (C2V_73_121),
	.C2V_3 (C2V_123_121),
	.C2V_4 (C2V_168_121),
	.C2V_5 (C2V_179_121),
	.C2V_6 (C2V_262_121),
	.L (L[1814:1800]),
	.V2C_1 (V2C_121_14),
	.V2C_2 (V2C_121_73),
	.V2C_3 (V2C_121_123),
	.V2C_4 (V2C_121_168),
	.V2C_5 (V2C_121_179),
	.V2C_6 (V2C_121_262),
	.V (V_121)
);

VNU_6 #(quan_width) VNU122 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_122),
	.C2V_2 (C2V_79_122),
	.C2V_3 (C2V_129_122),
	.C2V_4 (C2V_174_122),
	.C2V_5 (C2V_185_122),
	.C2V_6 (C2V_268_122),
	.L (L[1829:1815]),
	.V2C_1 (V2C_122_20),
	.V2C_2 (V2C_122_79),
	.V2C_3 (V2C_122_129),
	.V2C_4 (V2C_122_174),
	.V2C_5 (V2C_122_185),
	.V2C_6 (V2C_122_268),
	.V (V_122)
);

VNU_6 #(quan_width) VNU123 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_123),
	.C2V_2 (C2V_85_123),
	.C2V_3 (C2V_135_123),
	.C2V_4 (C2V_180_123),
	.C2V_5 (C2V_191_123),
	.C2V_6 (C2V_274_123),
	.L (L[1844:1830]),
	.V2C_1 (V2C_123_26),
	.V2C_2 (V2C_123_85),
	.V2C_3 (V2C_123_135),
	.V2C_4 (V2C_123_180),
	.V2C_5 (V2C_123_191),
	.V2C_6 (V2C_123_274),
	.V (V_123)
);

VNU_6 #(quan_width) VNU124 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_124),
	.C2V_2 (C2V_91_124),
	.C2V_3 (C2V_141_124),
	.C2V_4 (C2V_186_124),
	.C2V_5 (C2V_197_124),
	.C2V_6 (C2V_280_124),
	.L (L[1859:1845]),
	.V2C_1 (V2C_124_32),
	.V2C_2 (V2C_124_91),
	.V2C_3 (V2C_124_141),
	.V2C_4 (V2C_124_186),
	.V2C_5 (V2C_124_197),
	.V2C_6 (V2C_124_280),
	.V (V_124)
);

VNU_6 #(quan_width) VNU125 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_125),
	.C2V_2 (C2V_97_125),
	.C2V_3 (C2V_147_125),
	.C2V_4 (C2V_192_125),
	.C2V_5 (C2V_203_125),
	.C2V_6 (C2V_286_125),
	.L (L[1874:1860]),
	.V2C_1 (V2C_125_38),
	.V2C_2 (V2C_125_97),
	.V2C_3 (V2C_125_147),
	.V2C_4 (V2C_125_192),
	.V2C_5 (V2C_125_203),
	.V2C_6 (V2C_125_286),
	.V (V_125)
);

VNU_6 #(quan_width) VNU126 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_126),
	.C2V_2 (C2V_44_126),
	.C2V_3 (C2V_103_126),
	.C2V_4 (C2V_153_126),
	.C2V_5 (C2V_198_126),
	.C2V_6 (C2V_209_126),
	.L (L[1889:1875]),
	.V2C_1 (V2C_126_4),
	.V2C_2 (V2C_126_44),
	.V2C_3 (V2C_126_103),
	.V2C_4 (V2C_126_153),
	.V2C_5 (V2C_126_198),
	.V2C_6 (V2C_126_209),
	.V (V_126)
);

VNU_6 #(quan_width) VNU127 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_127),
	.C2V_2 (C2V_50_127),
	.C2V_3 (C2V_109_127),
	.C2V_4 (C2V_159_127),
	.C2V_5 (C2V_204_127),
	.C2V_6 (C2V_215_127),
	.L (L[1904:1890]),
	.V2C_1 (V2C_127_10),
	.V2C_2 (V2C_127_50),
	.V2C_3 (V2C_127_109),
	.V2C_4 (V2C_127_159),
	.V2C_5 (V2C_127_204),
	.V2C_6 (V2C_127_215),
	.V (V_127)
);

VNU_6 #(quan_width) VNU128 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_128),
	.C2V_2 (C2V_56_128),
	.C2V_3 (C2V_115_128),
	.C2V_4 (C2V_165_128),
	.C2V_5 (C2V_210_128),
	.C2V_6 (C2V_221_128),
	.L (L[1919:1905]),
	.V2C_1 (V2C_128_16),
	.V2C_2 (V2C_128_56),
	.V2C_3 (V2C_128_115),
	.V2C_4 (V2C_128_165),
	.V2C_5 (V2C_128_210),
	.V2C_6 (V2C_128_221),
	.V (V_128)
);

VNU_6 #(quan_width) VNU129 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_129),
	.C2V_2 (C2V_62_129),
	.C2V_3 (C2V_121_129),
	.C2V_4 (C2V_171_129),
	.C2V_5 (C2V_216_129),
	.C2V_6 (C2V_227_129),
	.L (L[1934:1920]),
	.V2C_1 (V2C_129_22),
	.V2C_2 (V2C_129_62),
	.V2C_3 (V2C_129_121),
	.V2C_4 (V2C_129_171),
	.V2C_5 (V2C_129_216),
	.V2C_6 (V2C_129_227),
	.V (V_129)
);

VNU_6 #(quan_width) VNU130 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_130),
	.C2V_2 (C2V_68_130),
	.C2V_3 (C2V_127_130),
	.C2V_4 (C2V_177_130),
	.C2V_5 (C2V_222_130),
	.C2V_6 (C2V_233_130),
	.L (L[1949:1935]),
	.V2C_1 (V2C_130_28),
	.V2C_2 (V2C_130_68),
	.V2C_3 (V2C_130_127),
	.V2C_4 (V2C_130_177),
	.V2C_5 (V2C_130_222),
	.V2C_6 (V2C_130_233),
	.V (V_130)
);

VNU_6 #(quan_width) VNU131 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_131),
	.C2V_2 (C2V_74_131),
	.C2V_3 (C2V_133_131),
	.C2V_4 (C2V_183_131),
	.C2V_5 (C2V_228_131),
	.C2V_6 (C2V_239_131),
	.L (L[1964:1950]),
	.V2C_1 (V2C_131_34),
	.V2C_2 (V2C_131_74),
	.V2C_3 (V2C_131_133),
	.V2C_4 (V2C_131_183),
	.V2C_5 (V2C_131_228),
	.V2C_6 (V2C_131_239),
	.V (V_131)
);

VNU_6 #(quan_width) VNU132 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_132),
	.C2V_2 (C2V_80_132),
	.C2V_3 (C2V_139_132),
	.C2V_4 (C2V_189_132),
	.C2V_5 (C2V_234_132),
	.C2V_6 (C2V_245_132),
	.L (L[1979:1965]),
	.V2C_1 (V2C_132_40),
	.V2C_2 (V2C_132_80),
	.V2C_3 (V2C_132_139),
	.V2C_4 (V2C_132_189),
	.V2C_5 (V2C_132_234),
	.V2C_6 (V2C_132_245),
	.V (V_132)
);

VNU_6 #(quan_width) VNU133 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_133),
	.C2V_2 (C2V_86_133),
	.C2V_3 (C2V_145_133),
	.C2V_4 (C2V_195_133),
	.C2V_5 (C2V_240_133),
	.C2V_6 (C2V_251_133),
	.L (L[1994:1980]),
	.V2C_1 (V2C_133_46),
	.V2C_2 (V2C_133_86),
	.V2C_3 (V2C_133_145),
	.V2C_4 (V2C_133_195),
	.V2C_5 (V2C_133_240),
	.V2C_6 (V2C_133_251),
	.V (V_133)
);

VNU_6 #(quan_width) VNU134 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_134),
	.C2V_2 (C2V_92_134),
	.C2V_3 (C2V_151_134),
	.C2V_4 (C2V_201_134),
	.C2V_5 (C2V_246_134),
	.C2V_6 (C2V_257_134),
	.L (L[2009:1995]),
	.V2C_1 (V2C_134_52),
	.V2C_2 (V2C_134_92),
	.V2C_3 (V2C_134_151),
	.V2C_4 (V2C_134_201),
	.V2C_5 (V2C_134_246),
	.V2C_6 (V2C_134_257),
	.V (V_134)
);

VNU_6 #(quan_width) VNU135 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_135),
	.C2V_2 (C2V_98_135),
	.C2V_3 (C2V_157_135),
	.C2V_4 (C2V_207_135),
	.C2V_5 (C2V_252_135),
	.C2V_6 (C2V_263_135),
	.L (L[2024:2010]),
	.V2C_1 (V2C_135_58),
	.V2C_2 (V2C_135_98),
	.V2C_3 (V2C_135_157),
	.V2C_4 (V2C_135_207),
	.V2C_5 (V2C_135_252),
	.V2C_6 (V2C_135_263),
	.V (V_135)
);

VNU_6 #(quan_width) VNU136 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_136),
	.C2V_2 (C2V_104_136),
	.C2V_3 (C2V_163_136),
	.C2V_4 (C2V_213_136),
	.C2V_5 (C2V_258_136),
	.C2V_6 (C2V_269_136),
	.L (L[2039:2025]),
	.V2C_1 (V2C_136_64),
	.V2C_2 (V2C_136_104),
	.V2C_3 (V2C_136_163),
	.V2C_4 (V2C_136_213),
	.V2C_5 (V2C_136_258),
	.V2C_6 (V2C_136_269),
	.V (V_136)
);

VNU_6 #(quan_width) VNU137 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_137),
	.C2V_2 (C2V_110_137),
	.C2V_3 (C2V_169_137),
	.C2V_4 (C2V_219_137),
	.C2V_5 (C2V_264_137),
	.C2V_6 (C2V_275_137),
	.L (L[2054:2040]),
	.V2C_1 (V2C_137_70),
	.V2C_2 (V2C_137_110),
	.V2C_3 (V2C_137_169),
	.V2C_4 (V2C_137_219),
	.V2C_5 (V2C_137_264),
	.V2C_6 (V2C_137_275),
	.V (V_137)
);

VNU_6 #(quan_width) VNU138 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_138),
	.C2V_2 (C2V_116_138),
	.C2V_3 (C2V_175_138),
	.C2V_4 (C2V_225_138),
	.C2V_5 (C2V_270_138),
	.C2V_6 (C2V_281_138),
	.L (L[2069:2055]),
	.V2C_1 (V2C_138_76),
	.V2C_2 (V2C_138_116),
	.V2C_3 (V2C_138_175),
	.V2C_4 (V2C_138_225),
	.V2C_5 (V2C_138_270),
	.V2C_6 (V2C_138_281),
	.V (V_138)
);

VNU_6 #(quan_width) VNU139 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_139),
	.C2V_2 (C2V_122_139),
	.C2V_3 (C2V_181_139),
	.C2V_4 (C2V_231_139),
	.C2V_5 (C2V_276_139),
	.C2V_6 (C2V_287_139),
	.L (L[2084:2070]),
	.V2C_1 (V2C_139_82),
	.V2C_2 (V2C_139_122),
	.V2C_3 (V2C_139_181),
	.V2C_4 (V2C_139_231),
	.V2C_5 (V2C_139_276),
	.V2C_6 (V2C_139_287),
	.V (V_139)
);

VNU_6 #(quan_width) VNU140 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_140),
	.C2V_2 (C2V_88_140),
	.C2V_3 (C2V_128_140),
	.C2V_4 (C2V_187_140),
	.C2V_5 (C2V_237_140),
	.C2V_6 (C2V_282_140),
	.L (L[2099:2085]),
	.V2C_1 (V2C_140_5),
	.V2C_2 (V2C_140_88),
	.V2C_3 (V2C_140_128),
	.V2C_4 (V2C_140_187),
	.V2C_5 (V2C_140_237),
	.V2C_6 (V2C_140_282),
	.V (V_140)
);

VNU_6 #(quan_width) VNU141 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_141),
	.C2V_2 (C2V_94_141),
	.C2V_3 (C2V_134_141),
	.C2V_4 (C2V_193_141),
	.C2V_5 (C2V_243_141),
	.C2V_6 (C2V_288_141),
	.L (L[2114:2100]),
	.V2C_1 (V2C_141_11),
	.V2C_2 (V2C_141_94),
	.V2C_3 (V2C_141_134),
	.V2C_4 (V2C_141_193),
	.V2C_5 (V2C_141_243),
	.V2C_6 (V2C_141_288),
	.V (V_141)
);

VNU_6 #(quan_width) VNU142 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_142),
	.C2V_2 (C2V_17_142),
	.C2V_3 (C2V_100_142),
	.C2V_4 (C2V_140_142),
	.C2V_5 (C2V_199_142),
	.C2V_6 (C2V_249_142),
	.L (L[2129:2115]),
	.V2C_1 (V2C_142_6),
	.V2C_2 (V2C_142_17),
	.V2C_3 (V2C_142_100),
	.V2C_4 (V2C_142_140),
	.V2C_5 (V2C_142_199),
	.V2C_6 (V2C_142_249),
	.V (V_142)
);

VNU_6 #(quan_width) VNU143 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_143),
	.C2V_2 (C2V_23_143),
	.C2V_3 (C2V_106_143),
	.C2V_4 (C2V_146_143),
	.C2V_5 (C2V_205_143),
	.C2V_6 (C2V_255_143),
	.L (L[2144:2130]),
	.V2C_1 (V2C_143_12),
	.V2C_2 (V2C_143_23),
	.V2C_3 (V2C_143_106),
	.V2C_4 (V2C_143_146),
	.V2C_5 (V2C_143_205),
	.V2C_6 (V2C_143_255),
	.V (V_143)
);

VNU_6 #(quan_width) VNU144 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_144),
	.C2V_2 (C2V_29_144),
	.C2V_3 (C2V_112_144),
	.C2V_4 (C2V_152_144),
	.C2V_5 (C2V_211_144),
	.C2V_6 (C2V_261_144),
	.L (L[2159:2145]),
	.V2C_1 (V2C_144_18),
	.V2C_2 (V2C_144_29),
	.V2C_3 (V2C_144_112),
	.V2C_4 (V2C_144_152),
	.V2C_5 (V2C_144_211),
	.V2C_6 (V2C_144_261),
	.V (V_144)
);

VNU_6 #(quan_width) VNU145 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_145),
	.C2V_2 (C2V_70_145),
	.C2V_3 (C2V_139_145),
	.C2V_4 (C2V_158_145),
	.C2V_5 (C2V_185_145),
	.C2V_6 (C2V_192_145),
	.L (L[2174:2160]),
	.V2C_1 (V2C_145_63),
	.V2C_2 (V2C_145_70),
	.V2C_3 (V2C_145_139),
	.V2C_4 (V2C_145_158),
	.V2C_5 (V2C_145_185),
	.V2C_6 (V2C_145_192),
	.V (V_145)
);

VNU_6 #(quan_width) VNU146 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_146),
	.C2V_2 (C2V_76_146),
	.C2V_3 (C2V_145_146),
	.C2V_4 (C2V_164_146),
	.C2V_5 (C2V_191_146),
	.C2V_6 (C2V_198_146),
	.L (L[2189:2175]),
	.V2C_1 (V2C_146_69),
	.V2C_2 (V2C_146_76),
	.V2C_3 (V2C_146_145),
	.V2C_4 (V2C_146_164),
	.V2C_5 (V2C_146_191),
	.V2C_6 (V2C_146_198),
	.V (V_146)
);

VNU_6 #(quan_width) VNU147 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_147),
	.C2V_2 (C2V_82_147),
	.C2V_3 (C2V_151_147),
	.C2V_4 (C2V_170_147),
	.C2V_5 (C2V_197_147),
	.C2V_6 (C2V_204_147),
	.L (L[2204:2190]),
	.V2C_1 (V2C_147_75),
	.V2C_2 (V2C_147_82),
	.V2C_3 (V2C_147_151),
	.V2C_4 (V2C_147_170),
	.V2C_5 (V2C_147_197),
	.V2C_6 (V2C_147_204),
	.V (V_147)
);

VNU_6 #(quan_width) VNU148 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_148),
	.C2V_2 (C2V_88_148),
	.C2V_3 (C2V_157_148),
	.C2V_4 (C2V_176_148),
	.C2V_5 (C2V_203_148),
	.C2V_6 (C2V_210_148),
	.L (L[2219:2205]),
	.V2C_1 (V2C_148_81),
	.V2C_2 (V2C_148_88),
	.V2C_3 (V2C_148_157),
	.V2C_4 (V2C_148_176),
	.V2C_5 (V2C_148_203),
	.V2C_6 (V2C_148_210),
	.V (V_148)
);

VNU_6 #(quan_width) VNU149 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_149),
	.C2V_2 (C2V_94_149),
	.C2V_3 (C2V_163_149),
	.C2V_4 (C2V_182_149),
	.C2V_5 (C2V_209_149),
	.C2V_6 (C2V_216_149),
	.L (L[2234:2220]),
	.V2C_1 (V2C_149_87),
	.V2C_2 (V2C_149_94),
	.V2C_3 (V2C_149_163),
	.V2C_4 (V2C_149_182),
	.V2C_5 (V2C_149_209),
	.V2C_6 (V2C_149_216),
	.V (V_149)
);

VNU_6 #(quan_width) VNU150 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_93_150),
	.C2V_2 (C2V_100_150),
	.C2V_3 (C2V_169_150),
	.C2V_4 (C2V_188_150),
	.C2V_5 (C2V_215_150),
	.C2V_6 (C2V_222_150),
	.L (L[2249:2235]),
	.V2C_1 (V2C_150_93),
	.V2C_2 (V2C_150_100),
	.V2C_3 (V2C_150_169),
	.V2C_4 (V2C_150_188),
	.V2C_5 (V2C_150_215),
	.V2C_6 (V2C_150_222),
	.V (V_150)
);

VNU_6 #(quan_width) VNU151 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_99_151),
	.C2V_2 (C2V_106_151),
	.C2V_3 (C2V_175_151),
	.C2V_4 (C2V_194_151),
	.C2V_5 (C2V_221_151),
	.C2V_6 (C2V_228_151),
	.L (L[2264:2250]),
	.V2C_1 (V2C_151_99),
	.V2C_2 (V2C_151_106),
	.V2C_3 (V2C_151_175),
	.V2C_4 (V2C_151_194),
	.V2C_5 (V2C_151_221),
	.V2C_6 (V2C_151_228),
	.V (V_151)
);

VNU_6 #(quan_width) VNU152 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_105_152),
	.C2V_2 (C2V_112_152),
	.C2V_3 (C2V_181_152),
	.C2V_4 (C2V_200_152),
	.C2V_5 (C2V_227_152),
	.C2V_6 (C2V_234_152),
	.L (L[2279:2265]),
	.V2C_1 (V2C_152_105),
	.V2C_2 (V2C_152_112),
	.V2C_3 (V2C_152_181),
	.V2C_4 (V2C_152_200),
	.V2C_5 (V2C_152_227),
	.V2C_6 (V2C_152_234),
	.V (V_152)
);

VNU_6 #(quan_width) VNU153 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_111_153),
	.C2V_2 (C2V_118_153),
	.C2V_3 (C2V_187_153),
	.C2V_4 (C2V_206_153),
	.C2V_5 (C2V_233_153),
	.C2V_6 (C2V_240_153),
	.L (L[2294:2280]),
	.V2C_1 (V2C_153_111),
	.V2C_2 (V2C_153_118),
	.V2C_3 (V2C_153_187),
	.V2C_4 (V2C_153_206),
	.V2C_5 (V2C_153_233),
	.V2C_6 (V2C_153_240),
	.V (V_153)
);

VNU_6 #(quan_width) VNU154 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_117_154),
	.C2V_2 (C2V_124_154),
	.C2V_3 (C2V_193_154),
	.C2V_4 (C2V_212_154),
	.C2V_5 (C2V_239_154),
	.C2V_6 (C2V_246_154),
	.L (L[2309:2295]),
	.V2C_1 (V2C_154_117),
	.V2C_2 (V2C_154_124),
	.V2C_3 (V2C_154_193),
	.V2C_4 (V2C_154_212),
	.V2C_5 (V2C_154_239),
	.V2C_6 (V2C_154_246),
	.V (V_154)
);

VNU_6 #(quan_width) VNU155 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_123_155),
	.C2V_2 (C2V_130_155),
	.C2V_3 (C2V_199_155),
	.C2V_4 (C2V_218_155),
	.C2V_5 (C2V_245_155),
	.C2V_6 (C2V_252_155),
	.L (L[2324:2310]),
	.V2C_1 (V2C_155_123),
	.V2C_2 (V2C_155_130),
	.V2C_3 (V2C_155_199),
	.V2C_4 (V2C_155_218),
	.V2C_5 (V2C_155_245),
	.V2C_6 (V2C_155_252),
	.V (V_155)
);

VNU_6 #(quan_width) VNU156 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_129_156),
	.C2V_2 (C2V_136_156),
	.C2V_3 (C2V_205_156),
	.C2V_4 (C2V_224_156),
	.C2V_5 (C2V_251_156),
	.C2V_6 (C2V_258_156),
	.L (L[2339:2325]),
	.V2C_1 (V2C_156_129),
	.V2C_2 (V2C_156_136),
	.V2C_3 (V2C_156_205),
	.V2C_4 (V2C_156_224),
	.V2C_5 (V2C_156_251),
	.V2C_6 (V2C_156_258),
	.V (V_156)
);

VNU_6 #(quan_width) VNU157 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_135_157),
	.C2V_2 (C2V_142_157),
	.C2V_3 (C2V_211_157),
	.C2V_4 (C2V_230_157),
	.C2V_5 (C2V_257_157),
	.C2V_6 (C2V_264_157),
	.L (L[2354:2340]),
	.V2C_1 (V2C_157_135),
	.V2C_2 (V2C_157_142),
	.V2C_3 (V2C_157_211),
	.V2C_4 (V2C_157_230),
	.V2C_5 (V2C_157_257),
	.V2C_6 (V2C_157_264),
	.V (V_157)
);

VNU_6 #(quan_width) VNU158 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_141_158),
	.C2V_2 (C2V_148_158),
	.C2V_3 (C2V_217_158),
	.C2V_4 (C2V_236_158),
	.C2V_5 (C2V_263_158),
	.C2V_6 (C2V_270_158),
	.L (L[2369:2355]),
	.V2C_1 (V2C_158_141),
	.V2C_2 (V2C_158_148),
	.V2C_3 (V2C_158_217),
	.V2C_4 (V2C_158_236),
	.V2C_5 (V2C_158_263),
	.V2C_6 (V2C_158_270),
	.V (V_158)
);

VNU_6 #(quan_width) VNU159 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_147_159),
	.C2V_2 (C2V_154_159),
	.C2V_3 (C2V_223_159),
	.C2V_4 (C2V_242_159),
	.C2V_5 (C2V_269_159),
	.C2V_6 (C2V_276_159),
	.L (L[2384:2370]),
	.V2C_1 (V2C_159_147),
	.V2C_2 (V2C_159_154),
	.V2C_3 (V2C_159_223),
	.V2C_4 (V2C_159_242),
	.V2C_5 (V2C_159_269),
	.V2C_6 (V2C_159_276),
	.V (V_159)
);

VNU_6 #(quan_width) VNU160 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_153_160),
	.C2V_2 (C2V_160_160),
	.C2V_3 (C2V_229_160),
	.C2V_4 (C2V_248_160),
	.C2V_5 (C2V_275_160),
	.C2V_6 (C2V_282_160),
	.L (L[2399:2385]),
	.V2C_1 (V2C_160_153),
	.V2C_2 (V2C_160_160),
	.V2C_3 (V2C_160_229),
	.V2C_4 (V2C_160_248),
	.V2C_5 (V2C_160_275),
	.V2C_6 (V2C_160_282),
	.V (V_160)
);

VNU_6 #(quan_width) VNU161 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_159_161),
	.C2V_2 (C2V_166_161),
	.C2V_3 (C2V_235_161),
	.C2V_4 (C2V_254_161),
	.C2V_5 (C2V_281_161),
	.C2V_6 (C2V_288_161),
	.L (L[2414:2400]),
	.V2C_1 (V2C_161_159),
	.V2C_2 (V2C_161_166),
	.V2C_3 (V2C_161_235),
	.V2C_4 (V2C_161_254),
	.V2C_5 (V2C_161_281),
	.V2C_6 (V2C_161_288),
	.V (V_161)
);

VNU_6 #(quan_width) VNU162 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_162),
	.C2V_2 (C2V_165_162),
	.C2V_3 (C2V_172_162),
	.C2V_4 (C2V_241_162),
	.C2V_5 (C2V_260_162),
	.C2V_6 (C2V_287_162),
	.L (L[2429:2415]),
	.V2C_1 (V2C_162_6),
	.V2C_2 (V2C_162_165),
	.V2C_3 (V2C_162_172),
	.V2C_4 (V2C_162_241),
	.V2C_5 (V2C_162_260),
	.V2C_6 (V2C_162_287),
	.V (V_162)
);

VNU_6 #(quan_width) VNU163 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_163),
	.C2V_2 (C2V_12_163),
	.C2V_3 (C2V_171_163),
	.C2V_4 (C2V_178_163),
	.C2V_5 (C2V_247_163),
	.C2V_6 (C2V_266_163),
	.L (L[2444:2430]),
	.V2C_1 (V2C_163_5),
	.V2C_2 (V2C_163_12),
	.V2C_3 (V2C_163_171),
	.V2C_4 (V2C_163_178),
	.V2C_5 (V2C_163_247),
	.V2C_6 (V2C_163_266),
	.V (V_163)
);

VNU_6 #(quan_width) VNU164 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_164),
	.C2V_2 (C2V_18_164),
	.C2V_3 (C2V_177_164),
	.C2V_4 (C2V_184_164),
	.C2V_5 (C2V_253_164),
	.C2V_6 (C2V_272_164),
	.L (L[2459:2445]),
	.V2C_1 (V2C_164_11),
	.V2C_2 (V2C_164_18),
	.V2C_3 (V2C_164_177),
	.V2C_4 (V2C_164_184),
	.V2C_5 (V2C_164_253),
	.V2C_6 (V2C_164_272),
	.V (V_164)
);

VNU_6 #(quan_width) VNU165 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_165),
	.C2V_2 (C2V_24_165),
	.C2V_3 (C2V_183_165),
	.C2V_4 (C2V_190_165),
	.C2V_5 (C2V_259_165),
	.C2V_6 (C2V_278_165),
	.L (L[2474:2460]),
	.V2C_1 (V2C_165_17),
	.V2C_2 (V2C_165_24),
	.V2C_3 (V2C_165_183),
	.V2C_4 (V2C_165_190),
	.V2C_5 (V2C_165_259),
	.V2C_6 (V2C_165_278),
	.V (V_165)
);

VNU_6 #(quan_width) VNU166 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_166),
	.C2V_2 (C2V_30_166),
	.C2V_3 (C2V_189_166),
	.C2V_4 (C2V_196_166),
	.C2V_5 (C2V_265_166),
	.C2V_6 (C2V_284_166),
	.L (L[2489:2475]),
	.V2C_1 (V2C_166_23),
	.V2C_2 (V2C_166_30),
	.V2C_3 (V2C_166_189),
	.V2C_4 (V2C_166_196),
	.V2C_5 (V2C_166_265),
	.V2C_6 (V2C_166_284),
	.V (V_166)
);

VNU_6 #(quan_width) VNU167 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_167),
	.C2V_2 (C2V_29_167),
	.C2V_3 (C2V_36_167),
	.C2V_4 (C2V_195_167),
	.C2V_5 (C2V_202_167),
	.C2V_6 (C2V_271_167),
	.L (L[2504:2490]),
	.V2C_1 (V2C_167_2),
	.V2C_2 (V2C_167_29),
	.V2C_3 (V2C_167_36),
	.V2C_4 (V2C_167_195),
	.V2C_5 (V2C_167_202),
	.V2C_6 (V2C_167_271),
	.V (V_167)
);

VNU_6 #(quan_width) VNU168 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_168),
	.C2V_2 (C2V_35_168),
	.C2V_3 (C2V_42_168),
	.C2V_4 (C2V_201_168),
	.C2V_5 (C2V_208_168),
	.C2V_6 (C2V_277_168),
	.L (L[2519:2505]),
	.V2C_1 (V2C_168_8),
	.V2C_2 (V2C_168_35),
	.V2C_3 (V2C_168_42),
	.V2C_4 (V2C_168_201),
	.V2C_5 (V2C_168_208),
	.V2C_6 (V2C_168_277),
	.V (V_168)
);

VNU_6 #(quan_width) VNU169 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_169),
	.C2V_2 (C2V_41_169),
	.C2V_3 (C2V_48_169),
	.C2V_4 (C2V_207_169),
	.C2V_5 (C2V_214_169),
	.C2V_6 (C2V_283_169),
	.L (L[2534:2520]),
	.V2C_1 (V2C_169_14),
	.V2C_2 (V2C_169_41),
	.V2C_3 (V2C_169_48),
	.V2C_4 (V2C_169_207),
	.V2C_5 (V2C_169_214),
	.V2C_6 (V2C_169_283),
	.V (V_169)
);

VNU_6 #(quan_width) VNU170 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_170),
	.C2V_2 (C2V_20_170),
	.C2V_3 (C2V_47_170),
	.C2V_4 (C2V_54_170),
	.C2V_5 (C2V_213_170),
	.C2V_6 (C2V_220_170),
	.L (L[2549:2535]),
	.V2C_1 (V2C_170_1),
	.V2C_2 (V2C_170_20),
	.V2C_3 (V2C_170_47),
	.V2C_4 (V2C_170_54),
	.V2C_5 (V2C_170_213),
	.V2C_6 (V2C_170_220),
	.V (V_170)
);

VNU_6 #(quan_width) VNU171 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_171),
	.C2V_2 (C2V_26_171),
	.C2V_3 (C2V_53_171),
	.C2V_4 (C2V_60_171),
	.C2V_5 (C2V_219_171),
	.C2V_6 (C2V_226_171),
	.L (L[2564:2550]),
	.V2C_1 (V2C_171_7),
	.V2C_2 (V2C_171_26),
	.V2C_3 (V2C_171_53),
	.V2C_4 (V2C_171_60),
	.V2C_5 (V2C_171_219),
	.V2C_6 (V2C_171_226),
	.V (V_171)
);

VNU_6 #(quan_width) VNU172 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_172),
	.C2V_2 (C2V_32_172),
	.C2V_3 (C2V_59_172),
	.C2V_4 (C2V_66_172),
	.C2V_5 (C2V_225_172),
	.C2V_6 (C2V_232_172),
	.L (L[2579:2565]),
	.V2C_1 (V2C_172_13),
	.V2C_2 (V2C_172_32),
	.V2C_3 (V2C_172_59),
	.V2C_4 (V2C_172_66),
	.V2C_5 (V2C_172_225),
	.V2C_6 (V2C_172_232),
	.V (V_172)
);

VNU_6 #(quan_width) VNU173 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_173),
	.C2V_2 (C2V_38_173),
	.C2V_3 (C2V_65_173),
	.C2V_4 (C2V_72_173),
	.C2V_5 (C2V_231_173),
	.C2V_6 (C2V_238_173),
	.L (L[2594:2580]),
	.V2C_1 (V2C_173_19),
	.V2C_2 (V2C_173_38),
	.V2C_3 (V2C_173_65),
	.V2C_4 (V2C_173_72),
	.V2C_5 (V2C_173_231),
	.V2C_6 (V2C_173_238),
	.V (V_173)
);

VNU_6 #(quan_width) VNU174 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_174),
	.C2V_2 (C2V_44_174),
	.C2V_3 (C2V_71_174),
	.C2V_4 (C2V_78_174),
	.C2V_5 (C2V_237_174),
	.C2V_6 (C2V_244_174),
	.L (L[2609:2595]),
	.V2C_1 (V2C_174_25),
	.V2C_2 (V2C_174_44),
	.V2C_3 (V2C_174_71),
	.V2C_4 (V2C_174_78),
	.V2C_5 (V2C_174_237),
	.V2C_6 (V2C_174_244),
	.V (V_174)
);

VNU_6 #(quan_width) VNU175 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_175),
	.C2V_2 (C2V_50_175),
	.C2V_3 (C2V_77_175),
	.C2V_4 (C2V_84_175),
	.C2V_5 (C2V_243_175),
	.C2V_6 (C2V_250_175),
	.L (L[2624:2610]),
	.V2C_1 (V2C_175_31),
	.V2C_2 (V2C_175_50),
	.V2C_3 (V2C_175_77),
	.V2C_4 (V2C_175_84),
	.V2C_5 (V2C_175_243),
	.V2C_6 (V2C_175_250),
	.V (V_175)
);

VNU_6 #(quan_width) VNU176 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_176),
	.C2V_2 (C2V_56_176),
	.C2V_3 (C2V_83_176),
	.C2V_4 (C2V_90_176),
	.C2V_5 (C2V_249_176),
	.C2V_6 (C2V_256_176),
	.L (L[2639:2625]),
	.V2C_1 (V2C_176_37),
	.V2C_2 (V2C_176_56),
	.V2C_3 (V2C_176_83),
	.V2C_4 (V2C_176_90),
	.V2C_5 (V2C_176_249),
	.V2C_6 (V2C_176_256),
	.V (V_176)
);

VNU_6 #(quan_width) VNU177 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_177),
	.C2V_2 (C2V_62_177),
	.C2V_3 (C2V_89_177),
	.C2V_4 (C2V_96_177),
	.C2V_5 (C2V_255_177),
	.C2V_6 (C2V_262_177),
	.L (L[2654:2640]),
	.V2C_1 (V2C_177_43),
	.V2C_2 (V2C_177_62),
	.V2C_3 (V2C_177_89),
	.V2C_4 (V2C_177_96),
	.V2C_5 (V2C_177_255),
	.V2C_6 (V2C_177_262),
	.V (V_177)
);

VNU_6 #(quan_width) VNU178 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_178),
	.C2V_2 (C2V_68_178),
	.C2V_3 (C2V_95_178),
	.C2V_4 (C2V_102_178),
	.C2V_5 (C2V_261_178),
	.C2V_6 (C2V_268_178),
	.L (L[2669:2655]),
	.V2C_1 (V2C_178_49),
	.V2C_2 (V2C_178_68),
	.V2C_3 (V2C_178_95),
	.V2C_4 (V2C_178_102),
	.V2C_5 (V2C_178_261),
	.V2C_6 (V2C_178_268),
	.V (V_178)
);

VNU_6 #(quan_width) VNU179 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_179),
	.C2V_2 (C2V_74_179),
	.C2V_3 (C2V_101_179),
	.C2V_4 (C2V_108_179),
	.C2V_5 (C2V_267_179),
	.C2V_6 (C2V_274_179),
	.L (L[2684:2670]),
	.V2C_1 (V2C_179_55),
	.V2C_2 (V2C_179_74),
	.V2C_3 (V2C_179_101),
	.V2C_4 (V2C_179_108),
	.V2C_5 (V2C_179_267),
	.V2C_6 (V2C_179_274),
	.V (V_179)
);

VNU_6 #(quan_width) VNU180 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_180),
	.C2V_2 (C2V_80_180),
	.C2V_3 (C2V_107_180),
	.C2V_4 (C2V_114_180),
	.C2V_5 (C2V_273_180),
	.C2V_6 (C2V_280_180),
	.L (L[2699:2685]),
	.V2C_1 (V2C_180_61),
	.V2C_2 (V2C_180_80),
	.V2C_3 (V2C_180_107),
	.V2C_4 (V2C_180_114),
	.V2C_5 (V2C_180_273),
	.V2C_6 (V2C_180_280),
	.V (V_180)
);

VNU_6 #(quan_width) VNU181 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_181),
	.C2V_2 (C2V_86_181),
	.C2V_3 (C2V_113_181),
	.C2V_4 (C2V_120_181),
	.C2V_5 (C2V_279_181),
	.C2V_6 (C2V_286_181),
	.L (L[2714:2700]),
	.V2C_1 (V2C_181_67),
	.V2C_2 (V2C_181_86),
	.V2C_3 (V2C_181_113),
	.V2C_4 (V2C_181_120),
	.V2C_5 (V2C_181_279),
	.V2C_6 (V2C_181_286),
	.V (V_181)
);

VNU_6 #(quan_width) VNU182 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_182),
	.C2V_2 (C2V_73_182),
	.C2V_3 (C2V_92_182),
	.C2V_4 (C2V_119_182),
	.C2V_5 (C2V_126_182),
	.C2V_6 (C2V_285_182),
	.L (L[2729:2715]),
	.V2C_1 (V2C_182_4),
	.V2C_2 (V2C_182_73),
	.V2C_3 (V2C_182_92),
	.V2C_4 (V2C_182_119),
	.V2C_5 (V2C_182_126),
	.V2C_6 (V2C_182_285),
	.V (V_182)
);

VNU_6 #(quan_width) VNU183 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_183),
	.C2V_2 (C2V_10_183),
	.C2V_3 (C2V_79_183),
	.C2V_4 (C2V_98_183),
	.C2V_5 (C2V_125_183),
	.C2V_6 (C2V_132_183),
	.L (L[2744:2730]),
	.V2C_1 (V2C_183_3),
	.V2C_2 (V2C_183_10),
	.V2C_3 (V2C_183_79),
	.V2C_4 (V2C_183_98),
	.V2C_5 (V2C_183_125),
	.V2C_6 (V2C_183_132),
	.V (V_183)
);

VNU_6 #(quan_width) VNU184 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_184),
	.C2V_2 (C2V_16_184),
	.C2V_3 (C2V_85_184),
	.C2V_4 (C2V_104_184),
	.C2V_5 (C2V_131_184),
	.C2V_6 (C2V_138_184),
	.L (L[2759:2745]),
	.V2C_1 (V2C_184_9),
	.V2C_2 (V2C_184_16),
	.V2C_3 (V2C_184_85),
	.V2C_4 (V2C_184_104),
	.V2C_5 (V2C_184_131),
	.V2C_6 (V2C_184_138),
	.V (V_184)
);

VNU_6 #(quan_width) VNU185 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_185),
	.C2V_2 (C2V_22_185),
	.C2V_3 (C2V_91_185),
	.C2V_4 (C2V_110_185),
	.C2V_5 (C2V_137_185),
	.C2V_6 (C2V_144_185),
	.L (L[2774:2760]),
	.V2C_1 (V2C_185_15),
	.V2C_2 (V2C_185_22),
	.V2C_3 (V2C_185_91),
	.V2C_4 (V2C_185_110),
	.V2C_5 (V2C_185_137),
	.V2C_6 (V2C_185_144),
	.V (V_185)
);

VNU_6 #(quan_width) VNU186 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_186),
	.C2V_2 (C2V_28_186),
	.C2V_3 (C2V_97_186),
	.C2V_4 (C2V_116_186),
	.C2V_5 (C2V_143_186),
	.C2V_6 (C2V_150_186),
	.L (L[2789:2775]),
	.V2C_1 (V2C_186_21),
	.V2C_2 (V2C_186_28),
	.V2C_3 (V2C_186_97),
	.V2C_4 (V2C_186_116),
	.V2C_5 (V2C_186_143),
	.V2C_6 (V2C_186_150),
	.V (V_186)
);

VNU_6 #(quan_width) VNU187 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_187),
	.C2V_2 (C2V_34_187),
	.C2V_3 (C2V_103_187),
	.C2V_4 (C2V_122_187),
	.C2V_5 (C2V_149_187),
	.C2V_6 (C2V_156_187),
	.L (L[2804:2790]),
	.V2C_1 (V2C_187_27),
	.V2C_2 (V2C_187_34),
	.V2C_3 (V2C_187_103),
	.V2C_4 (V2C_187_122),
	.V2C_5 (V2C_187_149),
	.V2C_6 (V2C_187_156),
	.V (V_187)
);

VNU_6 #(quan_width) VNU188 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_188),
	.C2V_2 (C2V_40_188),
	.C2V_3 (C2V_109_188),
	.C2V_4 (C2V_128_188),
	.C2V_5 (C2V_155_188),
	.C2V_6 (C2V_162_188),
	.L (L[2819:2805]),
	.V2C_1 (V2C_188_33),
	.V2C_2 (V2C_188_40),
	.V2C_3 (V2C_188_109),
	.V2C_4 (V2C_188_128),
	.V2C_5 (V2C_188_155),
	.V2C_6 (V2C_188_162),
	.V (V_188)
);

VNU_6 #(quan_width) VNU189 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_189),
	.C2V_2 (C2V_46_189),
	.C2V_3 (C2V_115_189),
	.C2V_4 (C2V_134_189),
	.C2V_5 (C2V_161_189),
	.C2V_6 (C2V_168_189),
	.L (L[2834:2820]),
	.V2C_1 (V2C_189_39),
	.V2C_2 (V2C_189_46),
	.V2C_3 (V2C_189_115),
	.V2C_4 (V2C_189_134),
	.V2C_5 (V2C_189_161),
	.V2C_6 (V2C_189_168),
	.V (V_189)
);

VNU_6 #(quan_width) VNU190 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_190),
	.C2V_2 (C2V_52_190),
	.C2V_3 (C2V_121_190),
	.C2V_4 (C2V_140_190),
	.C2V_5 (C2V_167_190),
	.C2V_6 (C2V_174_190),
	.L (L[2849:2835]),
	.V2C_1 (V2C_190_45),
	.V2C_2 (V2C_190_52),
	.V2C_3 (V2C_190_121),
	.V2C_4 (V2C_190_140),
	.V2C_5 (V2C_190_167),
	.V2C_6 (V2C_190_174),
	.V (V_190)
);

VNU_6 #(quan_width) VNU191 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_191),
	.C2V_2 (C2V_58_191),
	.C2V_3 (C2V_127_191),
	.C2V_4 (C2V_146_191),
	.C2V_5 (C2V_173_191),
	.C2V_6 (C2V_180_191),
	.L (L[2864:2850]),
	.V2C_1 (V2C_191_51),
	.V2C_2 (V2C_191_58),
	.V2C_3 (V2C_191_127),
	.V2C_4 (V2C_191_146),
	.V2C_5 (V2C_191_173),
	.V2C_6 (V2C_191_180),
	.V (V_191)
);

VNU_6 #(quan_width) VNU192 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_192),
	.C2V_2 (C2V_64_192),
	.C2V_3 (C2V_133_192),
	.C2V_4 (C2V_152_192),
	.C2V_5 (C2V_179_192),
	.C2V_6 (C2V_186_192),
	.L (L[2879:2865]),
	.V2C_1 (V2C_192_57),
	.V2C_2 (V2C_192_64),
	.V2C_3 (V2C_192_133),
	.V2C_4 (V2C_192_152),
	.V2C_5 (V2C_192_179),
	.V2C_6 (V2C_192_186),
	.V (V_192)
);

VNU_6 #(quan_width) VNU193 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_193),
	.C2V_2 (C2V_89_193),
	.C2V_3 (C2V_243_193),
	.C2V_4 (C2V_256_193),
	.C2V_5 (C2V_272_193),
	.C2V_6 (C2V_276_193),
	.L (L[2894:2880]),
	.V2C_1 (V2C_193_55),
	.V2C_2 (V2C_193_89),
	.V2C_3 (V2C_193_243),
	.V2C_4 (V2C_193_256),
	.V2C_5 (V2C_193_272),
	.V2C_6 (V2C_193_276),
	.V (V_193)
);

VNU_6 #(quan_width) VNU194 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_194),
	.C2V_2 (C2V_95_194),
	.C2V_3 (C2V_249_194),
	.C2V_4 (C2V_262_194),
	.C2V_5 (C2V_278_194),
	.C2V_6 (C2V_282_194),
	.L (L[2909:2895]),
	.V2C_1 (V2C_194_61),
	.V2C_2 (V2C_194_95),
	.V2C_3 (V2C_194_249),
	.V2C_4 (V2C_194_262),
	.V2C_5 (V2C_194_278),
	.V2C_6 (V2C_194_282),
	.V (V_194)
);

VNU_6 #(quan_width) VNU195 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_195),
	.C2V_2 (C2V_101_195),
	.C2V_3 (C2V_255_195),
	.C2V_4 (C2V_268_195),
	.C2V_5 (C2V_284_195),
	.C2V_6 (C2V_288_195),
	.L (L[2924:2910]),
	.V2C_1 (V2C_195_67),
	.V2C_2 (V2C_195_101),
	.V2C_3 (V2C_195_255),
	.V2C_4 (V2C_195_268),
	.V2C_5 (V2C_195_284),
	.V2C_6 (V2C_195_288),
	.V (V_195)
);

VNU_6 #(quan_width) VNU196 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_196),
	.C2V_2 (C2V_6_196),
	.C2V_3 (C2V_73_196),
	.C2V_4 (C2V_107_196),
	.C2V_5 (C2V_261_196),
	.C2V_6 (C2V_274_196),
	.L (L[2939:2925]),
	.V2C_1 (V2C_196_2),
	.V2C_2 (V2C_196_6),
	.V2C_3 (V2C_196_73),
	.V2C_4 (V2C_196_107),
	.V2C_5 (V2C_196_261),
	.V2C_6 (V2C_196_274),
	.V (V_196)
);

VNU_6 #(quan_width) VNU197 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_197),
	.C2V_2 (C2V_12_197),
	.C2V_3 (C2V_79_197),
	.C2V_4 (C2V_113_197),
	.C2V_5 (C2V_267_197),
	.C2V_6 (C2V_280_197),
	.L (L[2954:2940]),
	.V2C_1 (V2C_197_8),
	.V2C_2 (V2C_197_12),
	.V2C_3 (V2C_197_79),
	.V2C_4 (V2C_197_113),
	.V2C_5 (V2C_197_267),
	.V2C_6 (V2C_197_280),
	.V (V_197)
);

VNU_6 #(quan_width) VNU198 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_198),
	.C2V_2 (C2V_18_198),
	.C2V_3 (C2V_85_198),
	.C2V_4 (C2V_119_198),
	.C2V_5 (C2V_273_198),
	.C2V_6 (C2V_286_198),
	.L (L[2969:2955]),
	.V2C_1 (V2C_198_14),
	.V2C_2 (V2C_198_18),
	.V2C_3 (V2C_198_85),
	.V2C_4 (V2C_198_119),
	.V2C_5 (V2C_198_273),
	.V2C_6 (V2C_198_286),
	.V (V_198)
);

VNU_6 #(quan_width) VNU199 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_199),
	.C2V_2 (C2V_20_199),
	.C2V_3 (C2V_24_199),
	.C2V_4 (C2V_91_199),
	.C2V_5 (C2V_125_199),
	.C2V_6 (C2V_279_199),
	.L (L[2984:2970]),
	.V2C_1 (V2C_199_4),
	.V2C_2 (V2C_199_20),
	.V2C_3 (V2C_199_24),
	.V2C_4 (V2C_199_91),
	.V2C_5 (V2C_199_125),
	.V2C_6 (V2C_199_279),
	.V (V_199)
);

VNU_6 #(quan_width) VNU200 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_200),
	.C2V_2 (C2V_26_200),
	.C2V_3 (C2V_30_200),
	.C2V_4 (C2V_97_200),
	.C2V_5 (C2V_131_200),
	.C2V_6 (C2V_285_200),
	.L (L[2999:2985]),
	.V2C_1 (V2C_200_10),
	.V2C_2 (V2C_200_26),
	.V2C_3 (V2C_200_30),
	.V2C_4 (V2C_200_97),
	.V2C_5 (V2C_200_131),
	.V2C_6 (V2C_200_285),
	.V (V_200)
);

VNU_6 #(quan_width) VNU201 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_201),
	.C2V_2 (C2V_16_201),
	.C2V_3 (C2V_32_201),
	.C2V_4 (C2V_36_201),
	.C2V_5 (C2V_103_201),
	.C2V_6 (C2V_137_201),
	.L (L[3014:3000]),
	.V2C_1 (V2C_201_3),
	.V2C_2 (V2C_201_16),
	.V2C_3 (V2C_201_32),
	.V2C_4 (V2C_201_36),
	.V2C_5 (V2C_201_103),
	.V2C_6 (V2C_201_137),
	.V (V_201)
);

VNU_6 #(quan_width) VNU202 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_202),
	.C2V_2 (C2V_22_202),
	.C2V_3 (C2V_38_202),
	.C2V_4 (C2V_42_202),
	.C2V_5 (C2V_109_202),
	.C2V_6 (C2V_143_202),
	.L (L[3029:3015]),
	.V2C_1 (V2C_202_9),
	.V2C_2 (V2C_202_22),
	.V2C_3 (V2C_202_38),
	.V2C_4 (V2C_202_42),
	.V2C_5 (V2C_202_109),
	.V2C_6 (V2C_202_143),
	.V (V_202)
);

VNU_6 #(quan_width) VNU203 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_203),
	.C2V_2 (C2V_28_203),
	.C2V_3 (C2V_44_203),
	.C2V_4 (C2V_48_203),
	.C2V_5 (C2V_115_203),
	.C2V_6 (C2V_149_203),
	.L (L[3044:3030]),
	.V2C_1 (V2C_203_15),
	.V2C_2 (V2C_203_28),
	.V2C_3 (V2C_203_44),
	.V2C_4 (V2C_203_48),
	.V2C_5 (V2C_203_115),
	.V2C_6 (V2C_203_149),
	.V (V_203)
);

VNU_6 #(quan_width) VNU204 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_204),
	.C2V_2 (C2V_34_204),
	.C2V_3 (C2V_50_204),
	.C2V_4 (C2V_54_204),
	.C2V_5 (C2V_121_204),
	.C2V_6 (C2V_155_204),
	.L (L[3059:3045]),
	.V2C_1 (V2C_204_21),
	.V2C_2 (V2C_204_34),
	.V2C_3 (V2C_204_50),
	.V2C_4 (V2C_204_54),
	.V2C_5 (V2C_204_121),
	.V2C_6 (V2C_204_155),
	.V (V_204)
);

VNU_6 #(quan_width) VNU205 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_205),
	.C2V_2 (C2V_40_205),
	.C2V_3 (C2V_56_205),
	.C2V_4 (C2V_60_205),
	.C2V_5 (C2V_127_205),
	.C2V_6 (C2V_161_205),
	.L (L[3074:3060]),
	.V2C_1 (V2C_205_27),
	.V2C_2 (V2C_205_40),
	.V2C_3 (V2C_205_56),
	.V2C_4 (V2C_205_60),
	.V2C_5 (V2C_205_127),
	.V2C_6 (V2C_205_161),
	.V (V_205)
);

VNU_6 #(quan_width) VNU206 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_206),
	.C2V_2 (C2V_46_206),
	.C2V_3 (C2V_62_206),
	.C2V_4 (C2V_66_206),
	.C2V_5 (C2V_133_206),
	.C2V_6 (C2V_167_206),
	.L (L[3089:3075]),
	.V2C_1 (V2C_206_33),
	.V2C_2 (V2C_206_46),
	.V2C_3 (V2C_206_62),
	.V2C_4 (V2C_206_66),
	.V2C_5 (V2C_206_133),
	.V2C_6 (V2C_206_167),
	.V (V_206)
);

VNU_6 #(quan_width) VNU207 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_207),
	.C2V_2 (C2V_52_207),
	.C2V_3 (C2V_68_207),
	.C2V_4 (C2V_72_207),
	.C2V_5 (C2V_139_207),
	.C2V_6 (C2V_173_207),
	.L (L[3104:3090]),
	.V2C_1 (V2C_207_39),
	.V2C_2 (V2C_207_52),
	.V2C_3 (V2C_207_68),
	.V2C_4 (V2C_207_72),
	.V2C_5 (V2C_207_139),
	.V2C_6 (V2C_207_173),
	.V (V_207)
);

VNU_6 #(quan_width) VNU208 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_208),
	.C2V_2 (C2V_58_208),
	.C2V_3 (C2V_74_208),
	.C2V_4 (C2V_78_208),
	.C2V_5 (C2V_145_208),
	.C2V_6 (C2V_179_208),
	.L (L[3119:3105]),
	.V2C_1 (V2C_208_45),
	.V2C_2 (V2C_208_58),
	.V2C_3 (V2C_208_74),
	.V2C_4 (V2C_208_78),
	.V2C_5 (V2C_208_145),
	.V2C_6 (V2C_208_179),
	.V (V_208)
);

VNU_6 #(quan_width) VNU209 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_209),
	.C2V_2 (C2V_64_209),
	.C2V_3 (C2V_80_209),
	.C2V_4 (C2V_84_209),
	.C2V_5 (C2V_151_209),
	.C2V_6 (C2V_185_209),
	.L (L[3134:3120]),
	.V2C_1 (V2C_209_51),
	.V2C_2 (V2C_209_64),
	.V2C_3 (V2C_209_80),
	.V2C_4 (V2C_209_84),
	.V2C_5 (V2C_209_151),
	.V2C_6 (V2C_209_185),
	.V (V_209)
);

VNU_6 #(quan_width) VNU210 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_210),
	.C2V_2 (C2V_70_210),
	.C2V_3 (C2V_86_210),
	.C2V_4 (C2V_90_210),
	.C2V_5 (C2V_157_210),
	.C2V_6 (C2V_191_210),
	.L (L[3149:3135]),
	.V2C_1 (V2C_210_57),
	.V2C_2 (V2C_210_70),
	.V2C_3 (V2C_210_86),
	.V2C_4 (V2C_210_90),
	.V2C_5 (V2C_210_157),
	.V2C_6 (V2C_210_191),
	.V (V_210)
);

VNU_6 #(quan_width) VNU211 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_211),
	.C2V_2 (C2V_76_211),
	.C2V_3 (C2V_92_211),
	.C2V_4 (C2V_96_211),
	.C2V_5 (C2V_163_211),
	.C2V_6 (C2V_197_211),
	.L (L[3164:3150]),
	.V2C_1 (V2C_211_63),
	.V2C_2 (V2C_211_76),
	.V2C_3 (V2C_211_92),
	.V2C_4 (V2C_211_96),
	.V2C_5 (V2C_211_163),
	.V2C_6 (V2C_211_197),
	.V (V_211)
);

VNU_6 #(quan_width) VNU212 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_212),
	.C2V_2 (C2V_82_212),
	.C2V_3 (C2V_98_212),
	.C2V_4 (C2V_102_212),
	.C2V_5 (C2V_169_212),
	.C2V_6 (C2V_203_212),
	.L (L[3179:3165]),
	.V2C_1 (V2C_212_69),
	.V2C_2 (V2C_212_82),
	.V2C_3 (V2C_212_98),
	.V2C_4 (V2C_212_102),
	.V2C_5 (V2C_212_169),
	.V2C_6 (V2C_212_203),
	.V (V_212)
);

VNU_6 #(quan_width) VNU213 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_213),
	.C2V_2 (C2V_88_213),
	.C2V_3 (C2V_104_213),
	.C2V_4 (C2V_108_213),
	.C2V_5 (C2V_175_213),
	.C2V_6 (C2V_209_213),
	.L (L[3194:3180]),
	.V2C_1 (V2C_213_75),
	.V2C_2 (V2C_213_88),
	.V2C_3 (V2C_213_104),
	.V2C_4 (V2C_213_108),
	.V2C_5 (V2C_213_175),
	.V2C_6 (V2C_213_209),
	.V (V_213)
);

VNU_6 #(quan_width) VNU214 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_214),
	.C2V_2 (C2V_94_214),
	.C2V_3 (C2V_110_214),
	.C2V_4 (C2V_114_214),
	.C2V_5 (C2V_181_214),
	.C2V_6 (C2V_215_214),
	.L (L[3209:3195]),
	.V2C_1 (V2C_214_81),
	.V2C_2 (V2C_214_94),
	.V2C_3 (V2C_214_110),
	.V2C_4 (V2C_214_114),
	.V2C_5 (V2C_214_181),
	.V2C_6 (V2C_214_215),
	.V (V_214)
);

VNU_6 #(quan_width) VNU215 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_215),
	.C2V_2 (C2V_100_215),
	.C2V_3 (C2V_116_215),
	.C2V_4 (C2V_120_215),
	.C2V_5 (C2V_187_215),
	.C2V_6 (C2V_221_215),
	.L (L[3224:3210]),
	.V2C_1 (V2C_215_87),
	.V2C_2 (V2C_215_100),
	.V2C_3 (V2C_215_116),
	.V2C_4 (V2C_215_120),
	.V2C_5 (V2C_215_187),
	.V2C_6 (V2C_215_221),
	.V (V_215)
);

VNU_6 #(quan_width) VNU216 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_93_216),
	.C2V_2 (C2V_106_216),
	.C2V_3 (C2V_122_216),
	.C2V_4 (C2V_126_216),
	.C2V_5 (C2V_193_216),
	.C2V_6 (C2V_227_216),
	.L (L[3239:3225]),
	.V2C_1 (V2C_216_93),
	.V2C_2 (V2C_216_106),
	.V2C_3 (V2C_216_122),
	.V2C_4 (V2C_216_126),
	.V2C_5 (V2C_216_193),
	.V2C_6 (V2C_216_227),
	.V (V_216)
);

VNU_6 #(quan_width) VNU217 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_99_217),
	.C2V_2 (C2V_112_217),
	.C2V_3 (C2V_128_217),
	.C2V_4 (C2V_132_217),
	.C2V_5 (C2V_199_217),
	.C2V_6 (C2V_233_217),
	.L (L[3254:3240]),
	.V2C_1 (V2C_217_99),
	.V2C_2 (V2C_217_112),
	.V2C_3 (V2C_217_128),
	.V2C_4 (V2C_217_132),
	.V2C_5 (V2C_217_199),
	.V2C_6 (V2C_217_233),
	.V (V_217)
);

VNU_6 #(quan_width) VNU218 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_105_218),
	.C2V_2 (C2V_118_218),
	.C2V_3 (C2V_134_218),
	.C2V_4 (C2V_138_218),
	.C2V_5 (C2V_205_218),
	.C2V_6 (C2V_239_218),
	.L (L[3269:3255]),
	.V2C_1 (V2C_218_105),
	.V2C_2 (V2C_218_118),
	.V2C_3 (V2C_218_134),
	.V2C_4 (V2C_218_138),
	.V2C_5 (V2C_218_205),
	.V2C_6 (V2C_218_239),
	.V (V_218)
);

VNU_6 #(quan_width) VNU219 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_111_219),
	.C2V_2 (C2V_124_219),
	.C2V_3 (C2V_140_219),
	.C2V_4 (C2V_144_219),
	.C2V_5 (C2V_211_219),
	.C2V_6 (C2V_245_219),
	.L (L[3284:3270]),
	.V2C_1 (V2C_219_111),
	.V2C_2 (V2C_219_124),
	.V2C_3 (V2C_219_140),
	.V2C_4 (V2C_219_144),
	.V2C_5 (V2C_219_211),
	.V2C_6 (V2C_219_245),
	.V (V_219)
);

VNU_6 #(quan_width) VNU220 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_117_220),
	.C2V_2 (C2V_130_220),
	.C2V_3 (C2V_146_220),
	.C2V_4 (C2V_150_220),
	.C2V_5 (C2V_217_220),
	.C2V_6 (C2V_251_220),
	.L (L[3299:3285]),
	.V2C_1 (V2C_220_117),
	.V2C_2 (V2C_220_130),
	.V2C_3 (V2C_220_146),
	.V2C_4 (V2C_220_150),
	.V2C_5 (V2C_220_217),
	.V2C_6 (V2C_220_251),
	.V (V_220)
);

VNU_6 #(quan_width) VNU221 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_123_221),
	.C2V_2 (C2V_136_221),
	.C2V_3 (C2V_152_221),
	.C2V_4 (C2V_156_221),
	.C2V_5 (C2V_223_221),
	.C2V_6 (C2V_257_221),
	.L (L[3314:3300]),
	.V2C_1 (V2C_221_123),
	.V2C_2 (V2C_221_136),
	.V2C_3 (V2C_221_152),
	.V2C_4 (V2C_221_156),
	.V2C_5 (V2C_221_223),
	.V2C_6 (V2C_221_257),
	.V (V_221)
);

VNU_6 #(quan_width) VNU222 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_129_222),
	.C2V_2 (C2V_142_222),
	.C2V_3 (C2V_158_222),
	.C2V_4 (C2V_162_222),
	.C2V_5 (C2V_229_222),
	.C2V_6 (C2V_263_222),
	.L (L[3329:3315]),
	.V2C_1 (V2C_222_129),
	.V2C_2 (V2C_222_142),
	.V2C_3 (V2C_222_158),
	.V2C_4 (V2C_222_162),
	.V2C_5 (V2C_222_229),
	.V2C_6 (V2C_222_263),
	.V (V_222)
);

VNU_6 #(quan_width) VNU223 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_135_223),
	.C2V_2 (C2V_148_223),
	.C2V_3 (C2V_164_223),
	.C2V_4 (C2V_168_223),
	.C2V_5 (C2V_235_223),
	.C2V_6 (C2V_269_223),
	.L (L[3344:3330]),
	.V2C_1 (V2C_223_135),
	.V2C_2 (V2C_223_148),
	.V2C_3 (V2C_223_164),
	.V2C_4 (V2C_223_168),
	.V2C_5 (V2C_223_235),
	.V2C_6 (V2C_223_269),
	.V (V_223)
);

VNU_6 #(quan_width) VNU224 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_141_224),
	.C2V_2 (C2V_154_224),
	.C2V_3 (C2V_170_224),
	.C2V_4 (C2V_174_224),
	.C2V_5 (C2V_241_224),
	.C2V_6 (C2V_275_224),
	.L (L[3359:3345]),
	.V2C_1 (V2C_224_141),
	.V2C_2 (V2C_224_154),
	.V2C_3 (V2C_224_170),
	.V2C_4 (V2C_224_174),
	.V2C_5 (V2C_224_241),
	.V2C_6 (V2C_224_275),
	.V (V_224)
);

VNU_6 #(quan_width) VNU225 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_147_225),
	.C2V_2 (C2V_160_225),
	.C2V_3 (C2V_176_225),
	.C2V_4 (C2V_180_225),
	.C2V_5 (C2V_247_225),
	.C2V_6 (C2V_281_225),
	.L (L[3374:3360]),
	.V2C_1 (V2C_225_147),
	.V2C_2 (V2C_225_160),
	.V2C_3 (V2C_225_176),
	.V2C_4 (V2C_225_180),
	.V2C_5 (V2C_225_247),
	.V2C_6 (V2C_225_281),
	.V (V_225)
);

VNU_6 #(quan_width) VNU226 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_153_226),
	.C2V_2 (C2V_166_226),
	.C2V_3 (C2V_182_226),
	.C2V_4 (C2V_186_226),
	.C2V_5 (C2V_253_226),
	.C2V_6 (C2V_287_226),
	.L (L[3389:3375]),
	.V2C_1 (V2C_226_153),
	.V2C_2 (V2C_226_166),
	.V2C_3 (V2C_226_182),
	.V2C_4 (V2C_226_186),
	.V2C_5 (V2C_226_253),
	.V2C_6 (V2C_226_287),
	.V (V_226)
);

VNU_6 #(quan_width) VNU227 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_227),
	.C2V_2 (C2V_159_227),
	.C2V_3 (C2V_172_227),
	.C2V_4 (C2V_188_227),
	.C2V_5 (C2V_192_227),
	.C2V_6 (C2V_259_227),
	.L (L[3404:3390]),
	.V2C_1 (V2C_227_5),
	.V2C_2 (V2C_227_159),
	.V2C_3 (V2C_227_172),
	.V2C_4 (V2C_227_188),
	.V2C_5 (V2C_227_192),
	.V2C_6 (V2C_227_259),
	.V (V_227)
);

VNU_6 #(quan_width) VNU228 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_228),
	.C2V_2 (C2V_165_228),
	.C2V_3 (C2V_178_228),
	.C2V_4 (C2V_194_228),
	.C2V_5 (C2V_198_228),
	.C2V_6 (C2V_265_228),
	.L (L[3419:3405]),
	.V2C_1 (V2C_228_11),
	.V2C_2 (V2C_228_165),
	.V2C_3 (V2C_228_178),
	.V2C_4 (V2C_228_194),
	.V2C_5 (V2C_228_198),
	.V2C_6 (V2C_228_265),
	.V (V_228)
);

VNU_6 #(quan_width) VNU229 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_229),
	.C2V_2 (C2V_171_229),
	.C2V_3 (C2V_184_229),
	.C2V_4 (C2V_200_229),
	.C2V_5 (C2V_204_229),
	.C2V_6 (C2V_271_229),
	.L (L[3434:3420]),
	.V2C_1 (V2C_229_17),
	.V2C_2 (V2C_229_171),
	.V2C_3 (V2C_229_184),
	.V2C_4 (V2C_229_200),
	.V2C_5 (V2C_229_204),
	.V2C_6 (V2C_229_271),
	.V (V_229)
);

VNU_6 #(quan_width) VNU230 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_230),
	.C2V_2 (C2V_177_230),
	.C2V_3 (C2V_190_230),
	.C2V_4 (C2V_206_230),
	.C2V_5 (C2V_210_230),
	.C2V_6 (C2V_277_230),
	.L (L[3449:3435]),
	.V2C_1 (V2C_230_23),
	.V2C_2 (V2C_230_177),
	.V2C_3 (V2C_230_190),
	.V2C_4 (V2C_230_206),
	.V2C_5 (V2C_230_210),
	.V2C_6 (V2C_230_277),
	.V (V_230)
);

VNU_6 #(quan_width) VNU231 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_231),
	.C2V_2 (C2V_183_231),
	.C2V_3 (C2V_196_231),
	.C2V_4 (C2V_212_231),
	.C2V_5 (C2V_216_231),
	.C2V_6 (C2V_283_231),
	.L (L[3464:3450]),
	.V2C_1 (V2C_231_29),
	.V2C_2 (V2C_231_183),
	.V2C_3 (V2C_231_196),
	.V2C_4 (V2C_231_212),
	.V2C_5 (V2C_231_216),
	.V2C_6 (V2C_231_283),
	.V (V_231)
);

VNU_6 #(quan_width) VNU232 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_232),
	.C2V_2 (C2V_35_232),
	.C2V_3 (C2V_189_232),
	.C2V_4 (C2V_202_232),
	.C2V_5 (C2V_218_232),
	.C2V_6 (C2V_222_232),
	.L (L[3479:3465]),
	.V2C_1 (V2C_232_1),
	.V2C_2 (V2C_232_35),
	.V2C_3 (V2C_232_189),
	.V2C_4 (V2C_232_202),
	.V2C_5 (V2C_232_218),
	.V2C_6 (V2C_232_222),
	.V (V_232)
);

VNU_6 #(quan_width) VNU233 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_233),
	.C2V_2 (C2V_41_233),
	.C2V_3 (C2V_195_233),
	.C2V_4 (C2V_208_233),
	.C2V_5 (C2V_224_233),
	.C2V_6 (C2V_228_233),
	.L (L[3494:3480]),
	.V2C_1 (V2C_233_7),
	.V2C_2 (V2C_233_41),
	.V2C_3 (V2C_233_195),
	.V2C_4 (V2C_233_208),
	.V2C_5 (V2C_233_224),
	.V2C_6 (V2C_233_228),
	.V (V_233)
);

VNU_6 #(quan_width) VNU234 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_234),
	.C2V_2 (C2V_47_234),
	.C2V_3 (C2V_201_234),
	.C2V_4 (C2V_214_234),
	.C2V_5 (C2V_230_234),
	.C2V_6 (C2V_234_234),
	.L (L[3509:3495]),
	.V2C_1 (V2C_234_13),
	.V2C_2 (V2C_234_47),
	.V2C_3 (V2C_234_201),
	.V2C_4 (V2C_234_214),
	.V2C_5 (V2C_234_230),
	.V2C_6 (V2C_234_234),
	.V (V_234)
);

VNU_6 #(quan_width) VNU235 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_235),
	.C2V_2 (C2V_53_235),
	.C2V_3 (C2V_207_235),
	.C2V_4 (C2V_220_235),
	.C2V_5 (C2V_236_235),
	.C2V_6 (C2V_240_235),
	.L (L[3524:3510]),
	.V2C_1 (V2C_235_19),
	.V2C_2 (V2C_235_53),
	.V2C_3 (V2C_235_207),
	.V2C_4 (V2C_235_220),
	.V2C_5 (V2C_235_236),
	.V2C_6 (V2C_235_240),
	.V (V_235)
);

VNU_6 #(quan_width) VNU236 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_236),
	.C2V_2 (C2V_59_236),
	.C2V_3 (C2V_213_236),
	.C2V_4 (C2V_226_236),
	.C2V_5 (C2V_242_236),
	.C2V_6 (C2V_246_236),
	.L (L[3539:3525]),
	.V2C_1 (V2C_236_25),
	.V2C_2 (V2C_236_59),
	.V2C_3 (V2C_236_213),
	.V2C_4 (V2C_236_226),
	.V2C_5 (V2C_236_242),
	.V2C_6 (V2C_236_246),
	.V (V_236)
);

VNU_6 #(quan_width) VNU237 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_237),
	.C2V_2 (C2V_65_237),
	.C2V_3 (C2V_219_237),
	.C2V_4 (C2V_232_237),
	.C2V_5 (C2V_248_237),
	.C2V_6 (C2V_252_237),
	.L (L[3554:3540]),
	.V2C_1 (V2C_237_31),
	.V2C_2 (V2C_237_65),
	.V2C_3 (V2C_237_219),
	.V2C_4 (V2C_237_232),
	.V2C_5 (V2C_237_248),
	.V2C_6 (V2C_237_252),
	.V (V_237)
);

VNU_6 #(quan_width) VNU238 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_238),
	.C2V_2 (C2V_71_238),
	.C2V_3 (C2V_225_238),
	.C2V_4 (C2V_238_238),
	.C2V_5 (C2V_254_238),
	.C2V_6 (C2V_258_238),
	.L (L[3569:3555]),
	.V2C_1 (V2C_238_37),
	.V2C_2 (V2C_238_71),
	.V2C_3 (V2C_238_225),
	.V2C_4 (V2C_238_238),
	.V2C_5 (V2C_238_254),
	.V2C_6 (V2C_238_258),
	.V (V_238)
);

VNU_6 #(quan_width) VNU239 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_239),
	.C2V_2 (C2V_77_239),
	.C2V_3 (C2V_231_239),
	.C2V_4 (C2V_244_239),
	.C2V_5 (C2V_260_239),
	.C2V_6 (C2V_264_239),
	.L (L[3584:3570]),
	.V2C_1 (V2C_239_43),
	.V2C_2 (V2C_239_77),
	.V2C_3 (V2C_239_231),
	.V2C_4 (V2C_239_244),
	.V2C_5 (V2C_239_260),
	.V2C_6 (V2C_239_264),
	.V (V_239)
);

VNU_6 #(quan_width) VNU240 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_240),
	.C2V_2 (C2V_83_240),
	.C2V_3 (C2V_237_240),
	.C2V_4 (C2V_250_240),
	.C2V_5 (C2V_266_240),
	.C2V_6 (C2V_270_240),
	.L (L[3599:3585]),
	.V2C_1 (V2C_240_49),
	.V2C_2 (V2C_240_83),
	.V2C_3 (V2C_240_237),
	.V2C_4 (V2C_240_250),
	.V2C_5 (V2C_240_266),
	.V2C_6 (V2C_240_270),
	.V (V_240)
);

VNU_6 #(quan_width) VNU241 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_241),
	.C2V_2 (C2V_90_241),
	.C2V_3 (C2V_129_241),
	.C2V_4 (C2V_146_241),
	.C2V_5 (C2V_220_241),
	.C2V_6 (C2V_269_241),
	.L (L[3614:3600]),
	.V2C_1 (V2C_241_85),
	.V2C_2 (V2C_241_90),
	.V2C_3 (V2C_241_129),
	.V2C_4 (V2C_241_146),
	.V2C_5 (V2C_241_220),
	.V2C_6 (V2C_241_269),
	.V (V_241)
);

VNU_6 #(quan_width) VNU242 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_91_242),
	.C2V_2 (C2V_96_242),
	.C2V_3 (C2V_135_242),
	.C2V_4 (C2V_152_242),
	.C2V_5 (C2V_226_242),
	.C2V_6 (C2V_275_242),
	.L (L[3629:3615]),
	.V2C_1 (V2C_242_91),
	.V2C_2 (V2C_242_96),
	.V2C_3 (V2C_242_135),
	.V2C_4 (V2C_242_152),
	.V2C_5 (V2C_242_226),
	.V2C_6 (V2C_242_275),
	.V (V_242)
);

VNU_6 #(quan_width) VNU243 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_97_243),
	.C2V_2 (C2V_102_243),
	.C2V_3 (C2V_141_243),
	.C2V_4 (C2V_158_243),
	.C2V_5 (C2V_232_243),
	.C2V_6 (C2V_281_243),
	.L (L[3644:3630]),
	.V2C_1 (V2C_243_97),
	.V2C_2 (V2C_243_102),
	.V2C_3 (V2C_243_141),
	.V2C_4 (V2C_243_158),
	.V2C_5 (V2C_243_232),
	.V2C_6 (V2C_243_281),
	.V (V_243)
);

VNU_6 #(quan_width) VNU244 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_103_244),
	.C2V_2 (C2V_108_244),
	.C2V_3 (C2V_147_244),
	.C2V_4 (C2V_164_244),
	.C2V_5 (C2V_238_244),
	.C2V_6 (C2V_287_244),
	.L (L[3659:3645]),
	.V2C_1 (V2C_244_103),
	.V2C_2 (V2C_244_108),
	.V2C_3 (V2C_244_147),
	.V2C_4 (V2C_244_164),
	.V2C_5 (V2C_244_238),
	.V2C_6 (V2C_244_287),
	.V (V_244)
);

VNU_6 #(quan_width) VNU245 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_245),
	.C2V_2 (C2V_109_245),
	.C2V_3 (C2V_114_245),
	.C2V_4 (C2V_153_245),
	.C2V_5 (C2V_170_245),
	.C2V_6 (C2V_244_245),
	.L (L[3674:3660]),
	.V2C_1 (V2C_245_5),
	.V2C_2 (V2C_245_109),
	.V2C_3 (V2C_245_114),
	.V2C_4 (V2C_245_153),
	.V2C_5 (V2C_245_170),
	.V2C_6 (V2C_245_244),
	.V (V_245)
);

VNU_6 #(quan_width) VNU246 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_246),
	.C2V_2 (C2V_115_246),
	.C2V_3 (C2V_120_246),
	.C2V_4 (C2V_159_246),
	.C2V_5 (C2V_176_246),
	.C2V_6 (C2V_250_246),
	.L (L[3689:3675]),
	.V2C_1 (V2C_246_11),
	.V2C_2 (V2C_246_115),
	.V2C_3 (V2C_246_120),
	.V2C_4 (V2C_246_159),
	.V2C_5 (V2C_246_176),
	.V2C_6 (V2C_246_250),
	.V (V_246)
);

VNU_6 #(quan_width) VNU247 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_247),
	.C2V_2 (C2V_121_247),
	.C2V_3 (C2V_126_247),
	.C2V_4 (C2V_165_247),
	.C2V_5 (C2V_182_247),
	.C2V_6 (C2V_256_247),
	.L (L[3704:3690]),
	.V2C_1 (V2C_247_17),
	.V2C_2 (V2C_247_121),
	.V2C_3 (V2C_247_126),
	.V2C_4 (V2C_247_165),
	.V2C_5 (V2C_247_182),
	.V2C_6 (V2C_247_256),
	.V (V_247)
);

VNU_6 #(quan_width) VNU248 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_248),
	.C2V_2 (C2V_127_248),
	.C2V_3 (C2V_132_248),
	.C2V_4 (C2V_171_248),
	.C2V_5 (C2V_188_248),
	.C2V_6 (C2V_262_248),
	.L (L[3719:3705]),
	.V2C_1 (V2C_248_23),
	.V2C_2 (V2C_248_127),
	.V2C_3 (V2C_248_132),
	.V2C_4 (V2C_248_171),
	.V2C_5 (V2C_248_188),
	.V2C_6 (V2C_248_262),
	.V (V_248)
);

VNU_6 #(quan_width) VNU249 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_249),
	.C2V_2 (C2V_133_249),
	.C2V_3 (C2V_138_249),
	.C2V_4 (C2V_177_249),
	.C2V_5 (C2V_194_249),
	.C2V_6 (C2V_268_249),
	.L (L[3734:3720]),
	.V2C_1 (V2C_249_29),
	.V2C_2 (V2C_249_133),
	.V2C_3 (V2C_249_138),
	.V2C_4 (V2C_249_177),
	.V2C_5 (V2C_249_194),
	.V2C_6 (V2C_249_268),
	.V (V_249)
);

VNU_6 #(quan_width) VNU250 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_250),
	.C2V_2 (C2V_139_250),
	.C2V_3 (C2V_144_250),
	.C2V_4 (C2V_183_250),
	.C2V_5 (C2V_200_250),
	.C2V_6 (C2V_274_250),
	.L (L[3749:3735]),
	.V2C_1 (V2C_250_35),
	.V2C_2 (V2C_250_139),
	.V2C_3 (V2C_250_144),
	.V2C_4 (V2C_250_183),
	.V2C_5 (V2C_250_200),
	.V2C_6 (V2C_250_274),
	.V (V_250)
);

VNU_6 #(quan_width) VNU251 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_251),
	.C2V_2 (C2V_145_251),
	.C2V_3 (C2V_150_251),
	.C2V_4 (C2V_189_251),
	.C2V_5 (C2V_206_251),
	.C2V_6 (C2V_280_251),
	.L (L[3764:3750]),
	.V2C_1 (V2C_251_41),
	.V2C_2 (V2C_251_145),
	.V2C_3 (V2C_251_150),
	.V2C_4 (V2C_251_189),
	.V2C_5 (V2C_251_206),
	.V2C_6 (V2C_251_280),
	.V (V_251)
);

VNU_6 #(quan_width) VNU252 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_252),
	.C2V_2 (C2V_151_252),
	.C2V_3 (C2V_156_252),
	.C2V_4 (C2V_195_252),
	.C2V_5 (C2V_212_252),
	.C2V_6 (C2V_286_252),
	.L (L[3779:3765]),
	.V2C_1 (V2C_252_47),
	.V2C_2 (V2C_252_151),
	.V2C_3 (V2C_252_156),
	.V2C_4 (V2C_252_195),
	.V2C_5 (V2C_252_212),
	.V2C_6 (V2C_252_286),
	.V (V_252)
);

VNU_6 #(quan_width) VNU253 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_253),
	.C2V_2 (C2V_53_253),
	.C2V_3 (C2V_157_253),
	.C2V_4 (C2V_162_253),
	.C2V_5 (C2V_201_253),
	.C2V_6 (C2V_218_253),
	.L (L[3794:3780]),
	.V2C_1 (V2C_253_4),
	.V2C_2 (V2C_253_53),
	.V2C_3 (V2C_253_157),
	.V2C_4 (V2C_253_162),
	.V2C_5 (V2C_253_201),
	.V2C_6 (V2C_253_218),
	.V (V_253)
);

VNU_6 #(quan_width) VNU254 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_254),
	.C2V_2 (C2V_59_254),
	.C2V_3 (C2V_163_254),
	.C2V_4 (C2V_168_254),
	.C2V_5 (C2V_207_254),
	.C2V_6 (C2V_224_254),
	.L (L[3809:3795]),
	.V2C_1 (V2C_254_10),
	.V2C_2 (V2C_254_59),
	.V2C_3 (V2C_254_163),
	.V2C_4 (V2C_254_168),
	.V2C_5 (V2C_254_207),
	.V2C_6 (V2C_254_224),
	.V (V_254)
);

VNU_6 #(quan_width) VNU255 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_255),
	.C2V_2 (C2V_65_255),
	.C2V_3 (C2V_169_255),
	.C2V_4 (C2V_174_255),
	.C2V_5 (C2V_213_255),
	.C2V_6 (C2V_230_255),
	.L (L[3824:3810]),
	.V2C_1 (V2C_255_16),
	.V2C_2 (V2C_255_65),
	.V2C_3 (V2C_255_169),
	.V2C_4 (V2C_255_174),
	.V2C_5 (V2C_255_213),
	.V2C_6 (V2C_255_230),
	.V (V_255)
);

VNU_6 #(quan_width) VNU256 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_256),
	.C2V_2 (C2V_71_256),
	.C2V_3 (C2V_175_256),
	.C2V_4 (C2V_180_256),
	.C2V_5 (C2V_219_256),
	.C2V_6 (C2V_236_256),
	.L (L[3839:3825]),
	.V2C_1 (V2C_256_22),
	.V2C_2 (V2C_256_71),
	.V2C_3 (V2C_256_175),
	.V2C_4 (V2C_256_180),
	.V2C_5 (V2C_256_219),
	.V2C_6 (V2C_256_236),
	.V (V_256)
);

VNU_6 #(quan_width) VNU257 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_257),
	.C2V_2 (C2V_77_257),
	.C2V_3 (C2V_181_257),
	.C2V_4 (C2V_186_257),
	.C2V_5 (C2V_225_257),
	.C2V_6 (C2V_242_257),
	.L (L[3854:3840]),
	.V2C_1 (V2C_257_28),
	.V2C_2 (V2C_257_77),
	.V2C_3 (V2C_257_181),
	.V2C_4 (V2C_257_186),
	.V2C_5 (V2C_257_225),
	.V2C_6 (V2C_257_242),
	.V (V_257)
);

VNU_6 #(quan_width) VNU258 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_258),
	.C2V_2 (C2V_83_258),
	.C2V_3 (C2V_187_258),
	.C2V_4 (C2V_192_258),
	.C2V_5 (C2V_231_258),
	.C2V_6 (C2V_248_258),
	.L (L[3869:3855]),
	.V2C_1 (V2C_258_34),
	.V2C_2 (V2C_258_83),
	.V2C_3 (V2C_258_187),
	.V2C_4 (V2C_258_192),
	.V2C_5 (V2C_258_231),
	.V2C_6 (V2C_258_248),
	.V (V_258)
);

VNU_6 #(quan_width) VNU259 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_259),
	.C2V_2 (C2V_89_259),
	.C2V_3 (C2V_193_259),
	.C2V_4 (C2V_198_259),
	.C2V_5 (C2V_237_259),
	.C2V_6 (C2V_254_259),
	.L (L[3884:3870]),
	.V2C_1 (V2C_259_40),
	.V2C_2 (V2C_259_89),
	.V2C_3 (V2C_259_193),
	.V2C_4 (V2C_259_198),
	.V2C_5 (V2C_259_237),
	.V2C_6 (V2C_259_254),
	.V (V_259)
);

VNU_6 #(quan_width) VNU260 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_260),
	.C2V_2 (C2V_95_260),
	.C2V_3 (C2V_199_260),
	.C2V_4 (C2V_204_260),
	.C2V_5 (C2V_243_260),
	.C2V_6 (C2V_260_260),
	.L (L[3899:3885]),
	.V2C_1 (V2C_260_46),
	.V2C_2 (V2C_260_95),
	.V2C_3 (V2C_260_199),
	.V2C_4 (V2C_260_204),
	.V2C_5 (V2C_260_243),
	.V2C_6 (V2C_260_260),
	.V (V_260)
);

VNU_6 #(quan_width) VNU261 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_261),
	.C2V_2 (C2V_101_261),
	.C2V_3 (C2V_205_261),
	.C2V_4 (C2V_210_261),
	.C2V_5 (C2V_249_261),
	.C2V_6 (C2V_266_261),
	.L (L[3914:3900]),
	.V2C_1 (V2C_261_52),
	.V2C_2 (V2C_261_101),
	.V2C_3 (V2C_261_205),
	.V2C_4 (V2C_261_210),
	.V2C_5 (V2C_261_249),
	.V2C_6 (V2C_261_266),
	.V (V_261)
);

VNU_6 #(quan_width) VNU262 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_262),
	.C2V_2 (C2V_107_262),
	.C2V_3 (C2V_211_262),
	.C2V_4 (C2V_216_262),
	.C2V_5 (C2V_255_262),
	.C2V_6 (C2V_272_262),
	.L (L[3929:3915]),
	.V2C_1 (V2C_262_58),
	.V2C_2 (V2C_262_107),
	.V2C_3 (V2C_262_211),
	.V2C_4 (V2C_262_216),
	.V2C_5 (V2C_262_255),
	.V2C_6 (V2C_262_272),
	.V (V_262)
);

VNU_6 #(quan_width) VNU263 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_263),
	.C2V_2 (C2V_113_263),
	.C2V_3 (C2V_217_263),
	.C2V_4 (C2V_222_263),
	.C2V_5 (C2V_261_263),
	.C2V_6 (C2V_278_263),
	.L (L[3944:3930]),
	.V2C_1 (V2C_263_64),
	.V2C_2 (V2C_263_113),
	.V2C_3 (V2C_263_217),
	.V2C_4 (V2C_263_222),
	.V2C_5 (V2C_263_261),
	.V2C_6 (V2C_263_278),
	.V (V_263)
);

VNU_6 #(quan_width) VNU264 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_264),
	.C2V_2 (C2V_119_264),
	.C2V_3 (C2V_223_264),
	.C2V_4 (C2V_228_264),
	.C2V_5 (C2V_267_264),
	.C2V_6 (C2V_284_264),
	.L (L[3959:3945]),
	.V2C_1 (V2C_264_70),
	.V2C_2 (V2C_264_119),
	.V2C_3 (V2C_264_223),
	.V2C_4 (V2C_264_228),
	.V2C_5 (V2C_264_267),
	.V2C_6 (V2C_264_284),
	.V (V_264)
);

VNU_6 #(quan_width) VNU265 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_265),
	.C2V_2 (C2V_76_265),
	.C2V_3 (C2V_125_265),
	.C2V_4 (C2V_229_265),
	.C2V_5 (C2V_234_265),
	.C2V_6 (C2V_273_265),
	.L (L[3974:3960]),
	.V2C_1 (V2C_265_2),
	.V2C_2 (V2C_265_76),
	.V2C_3 (V2C_265_125),
	.V2C_4 (V2C_265_229),
	.V2C_5 (V2C_265_234),
	.V2C_6 (V2C_265_273),
	.V (V_265)
);

VNU_6 #(quan_width) VNU266 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_266),
	.C2V_2 (C2V_82_266),
	.C2V_3 (C2V_131_266),
	.C2V_4 (C2V_235_266),
	.C2V_5 (C2V_240_266),
	.C2V_6 (C2V_279_266),
	.L (L[3989:3975]),
	.V2C_1 (V2C_266_8),
	.V2C_2 (V2C_266_82),
	.V2C_3 (V2C_266_131),
	.V2C_4 (V2C_266_235),
	.V2C_5 (V2C_266_240),
	.V2C_6 (V2C_266_279),
	.V (V_266)
);

VNU_6 #(quan_width) VNU267 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_267),
	.C2V_2 (C2V_88_267),
	.C2V_3 (C2V_137_267),
	.C2V_4 (C2V_241_267),
	.C2V_5 (C2V_246_267),
	.C2V_6 (C2V_285_267),
	.L (L[4004:3990]),
	.V2C_1 (V2C_267_14),
	.V2C_2 (V2C_267_88),
	.V2C_3 (V2C_267_137),
	.V2C_4 (V2C_267_241),
	.V2C_5 (V2C_267_246),
	.V2C_6 (V2C_267_285),
	.V (V_267)
);

VNU_6 #(quan_width) VNU268 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_268),
	.C2V_2 (C2V_20_268),
	.C2V_3 (C2V_94_268),
	.C2V_4 (C2V_143_268),
	.C2V_5 (C2V_247_268),
	.C2V_6 (C2V_252_268),
	.L (L[4019:4005]),
	.V2C_1 (V2C_268_3),
	.V2C_2 (V2C_268_20),
	.V2C_3 (V2C_268_94),
	.V2C_4 (V2C_268_143),
	.V2C_5 (V2C_268_247),
	.V2C_6 (V2C_268_252),
	.V (V_268)
);

VNU_6 #(quan_width) VNU269 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_269),
	.C2V_2 (C2V_26_269),
	.C2V_3 (C2V_100_269),
	.C2V_4 (C2V_149_269),
	.C2V_5 (C2V_253_269),
	.C2V_6 (C2V_258_269),
	.L (L[4034:4020]),
	.V2C_1 (V2C_269_9),
	.V2C_2 (V2C_269_26),
	.V2C_3 (V2C_269_100),
	.V2C_4 (V2C_269_149),
	.V2C_5 (V2C_269_253),
	.V2C_6 (V2C_269_258),
	.V (V_269)
);

VNU_6 #(quan_width) VNU270 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_270),
	.C2V_2 (C2V_32_270),
	.C2V_3 (C2V_106_270),
	.C2V_4 (C2V_155_270),
	.C2V_5 (C2V_259_270),
	.C2V_6 (C2V_264_270),
	.L (L[4049:4035]),
	.V2C_1 (V2C_270_15),
	.V2C_2 (V2C_270_32),
	.V2C_3 (V2C_270_106),
	.V2C_4 (V2C_270_155),
	.V2C_5 (V2C_270_259),
	.V2C_6 (V2C_270_264),
	.V (V_270)
);

VNU_6 #(quan_width) VNU271 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_271),
	.C2V_2 (C2V_38_271),
	.C2V_3 (C2V_112_271),
	.C2V_4 (C2V_161_271),
	.C2V_5 (C2V_265_271),
	.C2V_6 (C2V_270_271),
	.L (L[4064:4050]),
	.V2C_1 (V2C_271_21),
	.V2C_2 (V2C_271_38),
	.V2C_3 (V2C_271_112),
	.V2C_4 (V2C_271_161),
	.V2C_5 (V2C_271_265),
	.V2C_6 (V2C_271_270),
	.V (V_271)
);

VNU_6 #(quan_width) VNU272 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_272),
	.C2V_2 (C2V_44_272),
	.C2V_3 (C2V_118_272),
	.C2V_4 (C2V_167_272),
	.C2V_5 (C2V_271_272),
	.C2V_6 (C2V_276_272),
	.L (L[4079:4065]),
	.V2C_1 (V2C_272_27),
	.V2C_2 (V2C_272_44),
	.V2C_3 (V2C_272_118),
	.V2C_4 (V2C_272_167),
	.V2C_5 (V2C_272_271),
	.V2C_6 (V2C_272_276),
	.V (V_272)
);

VNU_6 #(quan_width) VNU273 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_273),
	.C2V_2 (C2V_50_273),
	.C2V_3 (C2V_124_273),
	.C2V_4 (C2V_173_273),
	.C2V_5 (C2V_277_273),
	.C2V_6 (C2V_282_273),
	.L (L[4094:4080]),
	.V2C_1 (V2C_273_33),
	.V2C_2 (V2C_273_50),
	.V2C_3 (V2C_273_124),
	.V2C_4 (V2C_273_173),
	.V2C_5 (V2C_273_277),
	.V2C_6 (V2C_273_282),
	.V (V_273)
);

VNU_6 #(quan_width) VNU274 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_274),
	.C2V_2 (C2V_56_274),
	.C2V_3 (C2V_130_274),
	.C2V_4 (C2V_179_274),
	.C2V_5 (C2V_283_274),
	.C2V_6 (C2V_288_274),
	.L (L[4109:4095]),
	.V2C_1 (V2C_274_39),
	.V2C_2 (V2C_274_56),
	.V2C_3 (V2C_274_130),
	.V2C_4 (V2C_274_179),
	.V2C_5 (V2C_274_283),
	.V2C_6 (V2C_274_288),
	.V (V_274)
);

VNU_6 #(quan_width) VNU275 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_275),
	.C2V_2 (C2V_6_275),
	.C2V_3 (C2V_45_275),
	.C2V_4 (C2V_62_275),
	.C2V_5 (C2V_136_275),
	.C2V_6 (C2V_185_275),
	.L (L[4124:4110]),
	.V2C_1 (V2C_275_1),
	.V2C_2 (V2C_275_6),
	.V2C_3 (V2C_275_45),
	.V2C_4 (V2C_275_62),
	.V2C_5 (V2C_275_136),
	.V2C_6 (V2C_275_185),
	.V (V_275)
);

VNU_6 #(quan_width) VNU276 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_276),
	.C2V_2 (C2V_12_276),
	.C2V_3 (C2V_51_276),
	.C2V_4 (C2V_68_276),
	.C2V_5 (C2V_142_276),
	.C2V_6 (C2V_191_276),
	.L (L[4139:4125]),
	.V2C_1 (V2C_276_7),
	.V2C_2 (V2C_276_12),
	.V2C_3 (V2C_276_51),
	.V2C_4 (V2C_276_68),
	.V2C_5 (V2C_276_142),
	.V2C_6 (V2C_276_191),
	.V (V_276)
);

VNU_6 #(quan_width) VNU277 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_277),
	.C2V_2 (C2V_18_277),
	.C2V_3 (C2V_57_277),
	.C2V_4 (C2V_74_277),
	.C2V_5 (C2V_148_277),
	.C2V_6 (C2V_197_277),
	.L (L[4154:4140]),
	.V2C_1 (V2C_277_13),
	.V2C_2 (V2C_277_18),
	.V2C_3 (V2C_277_57),
	.V2C_4 (V2C_277_74),
	.V2C_5 (V2C_277_148),
	.V2C_6 (V2C_277_197),
	.V (V_277)
);

VNU_6 #(quan_width) VNU278 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_278),
	.C2V_2 (C2V_24_278),
	.C2V_3 (C2V_63_278),
	.C2V_4 (C2V_80_278),
	.C2V_5 (C2V_154_278),
	.C2V_6 (C2V_203_278),
	.L (L[4169:4155]),
	.V2C_1 (V2C_278_19),
	.V2C_2 (V2C_278_24),
	.V2C_3 (V2C_278_63),
	.V2C_4 (V2C_278_80),
	.V2C_5 (V2C_278_154),
	.V2C_6 (V2C_278_203),
	.V (V_278)
);

VNU_6 #(quan_width) VNU279 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_279),
	.C2V_2 (C2V_30_279),
	.C2V_3 (C2V_69_279),
	.C2V_4 (C2V_86_279),
	.C2V_5 (C2V_160_279),
	.C2V_6 (C2V_209_279),
	.L (L[4184:4170]),
	.V2C_1 (V2C_279_25),
	.V2C_2 (V2C_279_30),
	.V2C_3 (V2C_279_69),
	.V2C_4 (V2C_279_86),
	.V2C_5 (V2C_279_160),
	.V2C_6 (V2C_279_209),
	.V (V_279)
);

VNU_6 #(quan_width) VNU280 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_280),
	.C2V_2 (C2V_36_280),
	.C2V_3 (C2V_75_280),
	.C2V_4 (C2V_92_280),
	.C2V_5 (C2V_166_280),
	.C2V_6 (C2V_215_280),
	.L (L[4199:4185]),
	.V2C_1 (V2C_280_31),
	.V2C_2 (V2C_280_36),
	.V2C_3 (V2C_280_75),
	.V2C_4 (V2C_280_92),
	.V2C_5 (V2C_280_166),
	.V2C_6 (V2C_280_215),
	.V (V_280)
);

VNU_6 #(quan_width) VNU281 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_281),
	.C2V_2 (C2V_42_281),
	.C2V_3 (C2V_81_281),
	.C2V_4 (C2V_98_281),
	.C2V_5 (C2V_172_281),
	.C2V_6 (C2V_221_281),
	.L (L[4214:4200]),
	.V2C_1 (V2C_281_37),
	.V2C_2 (V2C_281_42),
	.V2C_3 (V2C_281_81),
	.V2C_4 (V2C_281_98),
	.V2C_5 (V2C_281_172),
	.V2C_6 (V2C_281_221),
	.V (V_281)
);

VNU_6 #(quan_width) VNU282 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_282),
	.C2V_2 (C2V_48_282),
	.C2V_3 (C2V_87_282),
	.C2V_4 (C2V_104_282),
	.C2V_5 (C2V_178_282),
	.C2V_6 (C2V_227_282),
	.L (L[4229:4215]),
	.V2C_1 (V2C_282_43),
	.V2C_2 (V2C_282_48),
	.V2C_3 (V2C_282_87),
	.V2C_4 (V2C_282_104),
	.V2C_5 (V2C_282_178),
	.V2C_6 (V2C_282_227),
	.V (V_282)
);

VNU_6 #(quan_width) VNU283 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_283),
	.C2V_2 (C2V_54_283),
	.C2V_3 (C2V_93_283),
	.C2V_4 (C2V_110_283),
	.C2V_5 (C2V_184_283),
	.C2V_6 (C2V_233_283),
	.L (L[4244:4230]),
	.V2C_1 (V2C_283_49),
	.V2C_2 (V2C_283_54),
	.V2C_3 (V2C_283_93),
	.V2C_4 (V2C_283_110),
	.V2C_5 (V2C_283_184),
	.V2C_6 (V2C_283_233),
	.V (V_283)
);

VNU_6 #(quan_width) VNU284 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_284),
	.C2V_2 (C2V_60_284),
	.C2V_3 (C2V_99_284),
	.C2V_4 (C2V_116_284),
	.C2V_5 (C2V_190_284),
	.C2V_6 (C2V_239_284),
	.L (L[4259:4245]),
	.V2C_1 (V2C_284_55),
	.V2C_2 (V2C_284_60),
	.V2C_3 (V2C_284_99),
	.V2C_4 (V2C_284_116),
	.V2C_5 (V2C_284_190),
	.V2C_6 (V2C_284_239),
	.V (V_284)
);

VNU_6 #(quan_width) VNU285 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_285),
	.C2V_2 (C2V_66_285),
	.C2V_3 (C2V_105_285),
	.C2V_4 (C2V_122_285),
	.C2V_5 (C2V_196_285),
	.C2V_6 (C2V_245_285),
	.L (L[4274:4260]),
	.V2C_1 (V2C_285_61),
	.V2C_2 (V2C_285_66),
	.V2C_3 (V2C_285_105),
	.V2C_4 (V2C_285_122),
	.V2C_5 (V2C_285_196),
	.V2C_6 (V2C_285_245),
	.V (V_285)
);

VNU_6 #(quan_width) VNU286 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_286),
	.C2V_2 (C2V_72_286),
	.C2V_3 (C2V_111_286),
	.C2V_4 (C2V_128_286),
	.C2V_5 (C2V_202_286),
	.C2V_6 (C2V_251_286),
	.L (L[4289:4275]),
	.V2C_1 (V2C_286_67),
	.V2C_2 (V2C_286_72),
	.V2C_3 (V2C_286_111),
	.V2C_4 (V2C_286_128),
	.V2C_5 (V2C_286_202),
	.V2C_6 (V2C_286_251),
	.V (V_286)
);

VNU_6 #(quan_width) VNU287 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_287),
	.C2V_2 (C2V_78_287),
	.C2V_3 (C2V_117_287),
	.C2V_4 (C2V_134_287),
	.C2V_5 (C2V_208_287),
	.C2V_6 (C2V_257_287),
	.L (L[4304:4290]),
	.V2C_1 (V2C_287_73),
	.V2C_2 (V2C_287_78),
	.V2C_3 (V2C_287_117),
	.V2C_4 (V2C_287_134),
	.V2C_5 (V2C_287_208),
	.V2C_6 (V2C_287_257),
	.V (V_287)
);

VNU_6 #(quan_width) VNU288 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_288),
	.C2V_2 (C2V_84_288),
	.C2V_3 (C2V_123_288),
	.C2V_4 (C2V_140_288),
	.C2V_5 (C2V_214_288),
	.C2V_6 (C2V_263_288),
	.L (L[4319:4305]),
	.V2C_1 (V2C_288_79),
	.V2C_2 (V2C_288_84),
	.V2C_3 (V2C_288_123),
	.V2C_4 (V2C_288_140),
	.V2C_5 (V2C_288_214),
	.V2C_6 (V2C_288_263),
	.V (V_288)
);

VNU_3 #(quan_width) VNU289 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_60_289),
	.C2V_2 (C2V_128_289),
	.C2V_3 (C2V_263_289),
	.L (L[4334:4320]),
	.V2C_1 (V2C_289_60),
	.V2C_2 (V2C_289_128),
	.V2C_3 (V2C_289_263),
	.V (V_289)
);

VNU_3 #(quan_width) VNU290 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_66_290),
	.C2V_2 (C2V_134_290),
	.C2V_3 (C2V_269_290),
	.L (L[4349:4335]),
	.V2C_1 (V2C_290_66),
	.V2C_2 (V2C_290_134),
	.V2C_3 (V2C_290_269),
	.V (V_290)
);

VNU_3 #(quan_width) VNU291 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_72_291),
	.C2V_2 (C2V_140_291),
	.C2V_3 (C2V_275_291),
	.L (L[4364:4350]),
	.V2C_1 (V2C_291_72),
	.V2C_2 (V2C_291_140),
	.V2C_3 (V2C_291_275),
	.V (V_291)
);

VNU_3 #(quan_width) VNU292 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_78_292),
	.C2V_2 (C2V_146_292),
	.C2V_3 (C2V_281_292),
	.L (L[4379:4365]),
	.V2C_1 (V2C_292_78),
	.V2C_2 (V2C_292_146),
	.V2C_3 (V2C_292_281),
	.V (V_292)
);

VNU_3 #(quan_width) VNU293 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_84_293),
	.C2V_2 (C2V_152_293),
	.C2V_3 (C2V_287_293),
	.L (L[4394:4380]),
	.V2C_1 (V2C_293_84),
	.V2C_2 (V2C_293_152),
	.V2C_3 (V2C_293_287),
	.V (V_293)
);

VNU_3 #(quan_width) VNU294 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_294),
	.C2V_2 (C2V_90_294),
	.C2V_3 (C2V_158_294),
	.L (L[4409:4395]),
	.V2C_1 (V2C_294_5),
	.V2C_2 (V2C_294_90),
	.V2C_3 (V2C_294_158),
	.V (V_294)
);

VNU_3 #(quan_width) VNU295 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_295),
	.C2V_2 (C2V_96_295),
	.C2V_3 (C2V_164_295),
	.L (L[4424:4410]),
	.V2C_1 (V2C_295_11),
	.V2C_2 (V2C_295_96),
	.V2C_3 (V2C_295_164),
	.V (V_295)
);

VNU_3 #(quan_width) VNU296 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_296),
	.C2V_2 (C2V_102_296),
	.C2V_3 (C2V_170_296),
	.L (L[4439:4425]),
	.V2C_1 (V2C_296_17),
	.V2C_2 (V2C_296_102),
	.V2C_3 (V2C_296_170),
	.V (V_296)
);

VNU_3 #(quan_width) VNU297 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_297),
	.C2V_2 (C2V_108_297),
	.C2V_3 (C2V_176_297),
	.L (L[4454:4440]),
	.V2C_1 (V2C_297_23),
	.V2C_2 (V2C_297_108),
	.V2C_3 (V2C_297_176),
	.V (V_297)
);

VNU_3 #(quan_width) VNU298 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_298),
	.C2V_2 (C2V_114_298),
	.C2V_3 (C2V_182_298),
	.L (L[4469:4455]),
	.V2C_1 (V2C_298_29),
	.V2C_2 (V2C_298_114),
	.V2C_3 (V2C_298_182),
	.V (V_298)
);

VNU_3 #(quan_width) VNU299 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_299),
	.C2V_2 (C2V_120_299),
	.C2V_3 (C2V_188_299),
	.L (L[4484:4470]),
	.V2C_1 (V2C_299_35),
	.V2C_2 (V2C_299_120),
	.V2C_3 (V2C_299_188),
	.V (V_299)
);

VNU_3 #(quan_width) VNU300 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_300),
	.C2V_2 (C2V_126_300),
	.C2V_3 (C2V_194_300),
	.L (L[4499:4485]),
	.V2C_1 (V2C_300_41),
	.V2C_2 (V2C_300_126),
	.V2C_3 (V2C_300_194),
	.V (V_300)
);

VNU_3 #(quan_width) VNU301 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_301),
	.C2V_2 (C2V_132_301),
	.C2V_3 (C2V_200_301),
	.L (L[4514:4500]),
	.V2C_1 (V2C_301_47),
	.V2C_2 (V2C_301_132),
	.V2C_3 (V2C_301_200),
	.V (V_301)
);

VNU_3 #(quan_width) VNU302 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_302),
	.C2V_2 (C2V_138_302),
	.C2V_3 (C2V_206_302),
	.L (L[4529:4515]),
	.V2C_1 (V2C_302_53),
	.V2C_2 (V2C_302_138),
	.V2C_3 (V2C_302_206),
	.V (V_302)
);

VNU_3 #(quan_width) VNU303 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_59_303),
	.C2V_2 (C2V_144_303),
	.C2V_3 (C2V_212_303),
	.L (L[4544:4530]),
	.V2C_1 (V2C_303_59),
	.V2C_2 (V2C_303_144),
	.V2C_3 (V2C_303_212),
	.V (V_303)
);

VNU_3 #(quan_width) VNU304 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_65_304),
	.C2V_2 (C2V_150_304),
	.C2V_3 (C2V_218_304),
	.L (L[4559:4545]),
	.V2C_1 (V2C_304_65),
	.V2C_2 (V2C_304_150),
	.V2C_3 (V2C_304_218),
	.V (V_304)
);

VNU_3 #(quan_width) VNU305 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_71_305),
	.C2V_2 (C2V_156_305),
	.C2V_3 (C2V_224_305),
	.L (L[4574:4560]),
	.V2C_1 (V2C_305_71),
	.V2C_2 (V2C_305_156),
	.V2C_3 (V2C_305_224),
	.V (V_305)
);

VNU_3 #(quan_width) VNU306 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_77_306),
	.C2V_2 (C2V_162_306),
	.C2V_3 (C2V_230_306),
	.L (L[4589:4575]),
	.V2C_1 (V2C_306_77),
	.V2C_2 (V2C_306_162),
	.V2C_3 (V2C_306_230),
	.V (V_306)
);

VNU_3 #(quan_width) VNU307 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_83_307),
	.C2V_2 (C2V_168_307),
	.C2V_3 (C2V_236_307),
	.L (L[4604:4590]),
	.V2C_1 (V2C_307_83),
	.V2C_2 (V2C_307_168),
	.V2C_3 (V2C_307_236),
	.V (V_307)
);

VNU_3 #(quan_width) VNU308 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_89_308),
	.C2V_2 (C2V_174_308),
	.C2V_3 (C2V_242_308),
	.L (L[4619:4605]),
	.V2C_1 (V2C_308_89),
	.V2C_2 (V2C_308_174),
	.V2C_3 (V2C_308_242),
	.V (V_308)
);

VNU_3 #(quan_width) VNU309 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_95_309),
	.C2V_2 (C2V_180_309),
	.C2V_3 (C2V_248_309),
	.L (L[4634:4620]),
	.V2C_1 (V2C_309_95),
	.V2C_2 (V2C_309_180),
	.V2C_3 (V2C_309_248),
	.V (V_309)
);

VNU_3 #(quan_width) VNU310 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_101_310),
	.C2V_2 (C2V_186_310),
	.C2V_3 (C2V_254_310),
	.L (L[4649:4635]),
	.V2C_1 (V2C_310_101),
	.V2C_2 (V2C_310_186),
	.V2C_3 (V2C_310_254),
	.V (V_310)
);

VNU_3 #(quan_width) VNU311 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_107_311),
	.C2V_2 (C2V_192_311),
	.C2V_3 (C2V_260_311),
	.L (L[4664:4650]),
	.V2C_1 (V2C_311_107),
	.V2C_2 (V2C_311_192),
	.V2C_3 (V2C_311_260),
	.V (V_311)
);

VNU_3 #(quan_width) VNU312 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_113_312),
	.C2V_2 (C2V_198_312),
	.C2V_3 (C2V_266_312),
	.L (L[4679:4665]),
	.V2C_1 (V2C_312_113),
	.V2C_2 (V2C_312_198),
	.V2C_3 (V2C_312_266),
	.V (V_312)
);

VNU_3 #(quan_width) VNU313 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_119_313),
	.C2V_2 (C2V_204_313),
	.C2V_3 (C2V_272_313),
	.L (L[4694:4680]),
	.V2C_1 (V2C_313_119),
	.V2C_2 (V2C_313_204),
	.V2C_3 (V2C_313_272),
	.V (V_313)
);

VNU_3 #(quan_width) VNU314 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_125_314),
	.C2V_2 (C2V_210_314),
	.C2V_3 (C2V_278_314),
	.L (L[4709:4695]),
	.V2C_1 (V2C_314_125),
	.V2C_2 (V2C_314_210),
	.V2C_3 (V2C_314_278),
	.V (V_314)
);

VNU_3 #(quan_width) VNU315 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_131_315),
	.C2V_2 (C2V_216_315),
	.C2V_3 (C2V_284_315),
	.L (L[4724:4710]),
	.V2C_1 (V2C_315_131),
	.V2C_2 (V2C_315_216),
	.V2C_3 (V2C_315_284),
	.V (V_315)
);

VNU_3 #(quan_width) VNU316 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_316),
	.C2V_2 (C2V_137_316),
	.C2V_3 (C2V_222_316),
	.L (L[4739:4725]),
	.V2C_1 (V2C_316_2),
	.V2C_2 (V2C_316_137),
	.V2C_3 (V2C_316_222),
	.V (V_316)
);

VNU_3 #(quan_width) VNU317 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_317),
	.C2V_2 (C2V_143_317),
	.C2V_3 (C2V_228_317),
	.L (L[4754:4740]),
	.V2C_1 (V2C_317_8),
	.V2C_2 (V2C_317_143),
	.V2C_3 (V2C_317_228),
	.V (V_317)
);

VNU_3 #(quan_width) VNU318 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_318),
	.C2V_2 (C2V_149_318),
	.C2V_3 (C2V_234_318),
	.L (L[4769:4755]),
	.V2C_1 (V2C_318_14),
	.V2C_2 (V2C_318_149),
	.V2C_3 (V2C_318_234),
	.V (V_318)
);

VNU_3 #(quan_width) VNU319 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_319),
	.C2V_2 (C2V_155_319),
	.C2V_3 (C2V_240_319),
	.L (L[4784:4770]),
	.V2C_1 (V2C_319_20),
	.V2C_2 (V2C_319_155),
	.V2C_3 (V2C_319_240),
	.V (V_319)
);

VNU_3 #(quan_width) VNU320 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_320),
	.C2V_2 (C2V_161_320),
	.C2V_3 (C2V_246_320),
	.L (L[4799:4785]),
	.V2C_1 (V2C_320_26),
	.V2C_2 (V2C_320_161),
	.V2C_3 (V2C_320_246),
	.V (V_320)
);

VNU_3 #(quan_width) VNU321 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_321),
	.C2V_2 (C2V_167_321),
	.C2V_3 (C2V_252_321),
	.L (L[4814:4800]),
	.V2C_1 (V2C_321_32),
	.V2C_2 (V2C_321_167),
	.V2C_3 (V2C_321_252),
	.V (V_321)
);

VNU_3 #(quan_width) VNU322 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_322),
	.C2V_2 (C2V_173_322),
	.C2V_3 (C2V_258_322),
	.L (L[4829:4815]),
	.V2C_1 (V2C_322_38),
	.V2C_2 (V2C_322_173),
	.V2C_3 (V2C_322_258),
	.V (V_322)
);

VNU_3 #(quan_width) VNU323 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_323),
	.C2V_2 (C2V_179_323),
	.C2V_3 (C2V_264_323),
	.L (L[4844:4830]),
	.V2C_1 (V2C_323_44),
	.V2C_2 (V2C_323_179),
	.V2C_3 (V2C_323_264),
	.V (V_323)
);

VNU_3 #(quan_width) VNU324 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_324),
	.C2V_2 (C2V_185_324),
	.C2V_3 (C2V_270_324),
	.L (L[4859:4845]),
	.V2C_1 (V2C_324_50),
	.V2C_2 (V2C_324_185),
	.V2C_3 (V2C_324_270),
	.V (V_324)
);

VNU_3 #(quan_width) VNU325 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_325),
	.C2V_2 (C2V_191_325),
	.C2V_3 (C2V_276_325),
	.L (L[4874:4860]),
	.V2C_1 (V2C_325_56),
	.V2C_2 (V2C_325_191),
	.V2C_3 (V2C_325_276),
	.V (V_325)
);

VNU_3 #(quan_width) VNU326 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_326),
	.C2V_2 (C2V_197_326),
	.C2V_3 (C2V_282_326),
	.L (L[4889:4875]),
	.V2C_1 (V2C_326_62),
	.V2C_2 (V2C_326_197),
	.V2C_3 (V2C_326_282),
	.V (V_326)
);

VNU_3 #(quan_width) VNU327 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_327),
	.C2V_2 (C2V_203_327),
	.C2V_3 (C2V_288_327),
	.L (L[4904:4890]),
	.V2C_1 (V2C_327_68),
	.V2C_2 (V2C_327_203),
	.V2C_3 (V2C_327_288),
	.V (V_327)
);

VNU_3 #(quan_width) VNU328 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_328),
	.C2V_2 (C2V_74_328),
	.C2V_3 (C2V_209_328),
	.L (L[4919:4905]),
	.V2C_1 (V2C_328_6),
	.V2C_2 (V2C_328_74),
	.V2C_3 (V2C_328_209),
	.V (V_328)
);

VNU_3 #(quan_width) VNU329 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_329),
	.C2V_2 (C2V_80_329),
	.C2V_3 (C2V_215_329),
	.L (L[4934:4920]),
	.V2C_1 (V2C_329_12),
	.V2C_2 (V2C_329_80),
	.V2C_3 (V2C_329_215),
	.V (V_329)
);

VNU_3 #(quan_width) VNU330 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_330),
	.C2V_2 (C2V_86_330),
	.C2V_3 (C2V_221_330),
	.L (L[4949:4935]),
	.V2C_1 (V2C_330_18),
	.V2C_2 (V2C_330_86),
	.V2C_3 (V2C_330_221),
	.V (V_330)
);

VNU_3 #(quan_width) VNU331 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_331),
	.C2V_2 (C2V_92_331),
	.C2V_3 (C2V_227_331),
	.L (L[4964:4950]),
	.V2C_1 (V2C_331_24),
	.V2C_2 (V2C_331_92),
	.V2C_3 (V2C_331_227),
	.V (V_331)
);

VNU_3 #(quan_width) VNU332 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_332),
	.C2V_2 (C2V_98_332),
	.C2V_3 (C2V_233_332),
	.L (L[4979:4965]),
	.V2C_1 (V2C_332_30),
	.V2C_2 (V2C_332_98),
	.V2C_3 (V2C_332_233),
	.V (V_332)
);

VNU_3 #(quan_width) VNU333 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_333),
	.C2V_2 (C2V_104_333),
	.C2V_3 (C2V_239_333),
	.L (L[4994:4980]),
	.V2C_1 (V2C_333_36),
	.V2C_2 (V2C_333_104),
	.V2C_3 (V2C_333_239),
	.V (V_333)
);

VNU_3 #(quan_width) VNU334 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_334),
	.C2V_2 (C2V_110_334),
	.C2V_3 (C2V_245_334),
	.L (L[5009:4995]),
	.V2C_1 (V2C_334_42),
	.V2C_2 (V2C_334_110),
	.V2C_3 (V2C_334_245),
	.V (V_334)
);

VNU_3 #(quan_width) VNU335 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_335),
	.C2V_2 (C2V_116_335),
	.C2V_3 (C2V_251_335),
	.L (L[5024:5010]),
	.V2C_1 (V2C_335_48),
	.V2C_2 (V2C_335_116),
	.V2C_3 (V2C_335_251),
	.V (V_335)
);

VNU_3 #(quan_width) VNU336 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_54_336),
	.C2V_2 (C2V_122_336),
	.C2V_3 (C2V_257_336),
	.L (L[5039:5025]),
	.V2C_1 (V2C_336_54),
	.V2C_2 (V2C_336_122),
	.V2C_3 (V2C_336_257),
	.V (V_336)
);

VNU_3 #(quan_width) VNU337 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_337),
	.C2V_2 (C2V_123_337),
	.C2V_3 (C2V_149_337),
	.L (L[5054:5040]),
	.V2C_1 (V2C_337_61),
	.V2C_2 (V2C_337_123),
	.V2C_3 (V2C_337_149),
	.V (V_337)
);

VNU_3 #(quan_width) VNU338 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_338),
	.C2V_2 (C2V_129_338),
	.C2V_3 (C2V_155_338),
	.L (L[5069:5055]),
	.V2C_1 (V2C_338_67),
	.V2C_2 (V2C_338_129),
	.V2C_3 (V2C_338_155),
	.V (V_338)
);

VNU_3 #(quan_width) VNU339 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_339),
	.C2V_2 (C2V_135_339),
	.C2V_3 (C2V_161_339),
	.L (L[5084:5070]),
	.V2C_1 (V2C_339_73),
	.V2C_2 (V2C_339_135),
	.V2C_3 (V2C_339_161),
	.V (V_339)
);

VNU_3 #(quan_width) VNU340 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_340),
	.C2V_2 (C2V_141_340),
	.C2V_3 (C2V_167_340),
	.L (L[5099:5085]),
	.V2C_1 (V2C_340_79),
	.V2C_2 (V2C_340_141),
	.V2C_3 (V2C_340_167),
	.V (V_340)
);

VNU_3 #(quan_width) VNU341 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_341),
	.C2V_2 (C2V_147_341),
	.C2V_3 (C2V_173_341),
	.L (L[5114:5100]),
	.V2C_1 (V2C_341_85),
	.V2C_2 (V2C_341_147),
	.V2C_3 (V2C_341_173),
	.V (V_341)
);

VNU_3 #(quan_width) VNU342 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_91_342),
	.C2V_2 (C2V_153_342),
	.C2V_3 (C2V_179_342),
	.L (L[5129:5115]),
	.V2C_1 (V2C_342_91),
	.V2C_2 (V2C_342_153),
	.V2C_3 (V2C_342_179),
	.V (V_342)
);

VNU_3 #(quan_width) VNU343 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_97_343),
	.C2V_2 (C2V_159_343),
	.C2V_3 (C2V_185_343),
	.L (L[5144:5130]),
	.V2C_1 (V2C_343_97),
	.V2C_2 (V2C_343_159),
	.V2C_3 (V2C_343_185),
	.V (V_343)
);

VNU_3 #(quan_width) VNU344 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_103_344),
	.C2V_2 (C2V_165_344),
	.C2V_3 (C2V_191_344),
	.L (L[5159:5145]),
	.V2C_1 (V2C_344_103),
	.V2C_2 (V2C_344_165),
	.V2C_3 (V2C_344_191),
	.V (V_344)
);

VNU_3 #(quan_width) VNU345 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_109_345),
	.C2V_2 (C2V_171_345),
	.C2V_3 (C2V_197_345),
	.L (L[5174:5160]),
	.V2C_1 (V2C_345_109),
	.V2C_2 (V2C_345_171),
	.V2C_3 (V2C_345_197),
	.V (V_345)
);

VNU_3 #(quan_width) VNU346 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_115_346),
	.C2V_2 (C2V_177_346),
	.C2V_3 (C2V_203_346),
	.L (L[5189:5175]),
	.V2C_1 (V2C_346_115),
	.V2C_2 (V2C_346_177),
	.V2C_3 (V2C_346_203),
	.V (V_346)
);

VNU_3 #(quan_width) VNU347 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_121_347),
	.C2V_2 (C2V_183_347),
	.C2V_3 (C2V_209_347),
	.L (L[5204:5190]),
	.V2C_1 (V2C_347_121),
	.V2C_2 (V2C_347_183),
	.V2C_3 (V2C_347_209),
	.V (V_347)
);

VNU_3 #(quan_width) VNU348 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_127_348),
	.C2V_2 (C2V_189_348),
	.C2V_3 (C2V_215_348),
	.L (L[5219:5205]),
	.V2C_1 (V2C_348_127),
	.V2C_2 (V2C_348_189),
	.V2C_3 (V2C_348_215),
	.V (V_348)
);

VNU_3 #(quan_width) VNU349 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_133_349),
	.C2V_2 (C2V_195_349),
	.C2V_3 (C2V_221_349),
	.L (L[5234:5220]),
	.V2C_1 (V2C_349_133),
	.V2C_2 (V2C_349_195),
	.V2C_3 (V2C_349_221),
	.V (V_349)
);

VNU_3 #(quan_width) VNU350 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_139_350),
	.C2V_2 (C2V_201_350),
	.C2V_3 (C2V_227_350),
	.L (L[5249:5235]),
	.V2C_1 (V2C_350_139),
	.V2C_2 (V2C_350_201),
	.V2C_3 (V2C_350_227),
	.V (V_350)
);

VNU_3 #(quan_width) VNU351 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_145_351),
	.C2V_2 (C2V_207_351),
	.C2V_3 (C2V_233_351),
	.L (L[5264:5250]),
	.V2C_1 (V2C_351_145),
	.V2C_2 (V2C_351_207),
	.V2C_3 (V2C_351_233),
	.V (V_351)
);

VNU_3 #(quan_width) VNU352 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_151_352),
	.C2V_2 (C2V_213_352),
	.C2V_3 (C2V_239_352),
	.L (L[5279:5265]),
	.V2C_1 (V2C_352_151),
	.V2C_2 (V2C_352_213),
	.V2C_3 (V2C_352_239),
	.V (V_352)
);

VNU_3 #(quan_width) VNU353 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_157_353),
	.C2V_2 (C2V_219_353),
	.C2V_3 (C2V_245_353),
	.L (L[5294:5280]),
	.V2C_1 (V2C_353_157),
	.V2C_2 (V2C_353_219),
	.V2C_3 (V2C_353_245),
	.V (V_353)
);

VNU_3 #(quan_width) VNU354 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_163_354),
	.C2V_2 (C2V_225_354),
	.C2V_3 (C2V_251_354),
	.L (L[5309:5295]),
	.V2C_1 (V2C_354_163),
	.V2C_2 (V2C_354_225),
	.V2C_3 (V2C_354_251),
	.V (V_354)
);

VNU_3 #(quan_width) VNU355 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_169_355),
	.C2V_2 (C2V_231_355),
	.C2V_3 (C2V_257_355),
	.L (L[5324:5310]),
	.V2C_1 (V2C_355_169),
	.V2C_2 (V2C_355_231),
	.V2C_3 (V2C_355_257),
	.V (V_355)
);

VNU_3 #(quan_width) VNU356 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_175_356),
	.C2V_2 (C2V_237_356),
	.C2V_3 (C2V_263_356),
	.L (L[5339:5325]),
	.V2C_1 (V2C_356_175),
	.V2C_2 (V2C_356_237),
	.V2C_3 (V2C_356_263),
	.V (V_356)
);

VNU_3 #(quan_width) VNU357 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_181_357),
	.C2V_2 (C2V_243_357),
	.C2V_3 (C2V_269_357),
	.L (L[5354:5340]),
	.V2C_1 (V2C_357_181),
	.V2C_2 (V2C_357_243),
	.V2C_3 (V2C_357_269),
	.V (V_357)
);

VNU_3 #(quan_width) VNU358 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_187_358),
	.C2V_2 (C2V_249_358),
	.C2V_3 (C2V_275_358),
	.L (L[5369:5355]),
	.V2C_1 (V2C_358_187),
	.V2C_2 (V2C_358_249),
	.V2C_3 (V2C_358_275),
	.V (V_358)
);

VNU_3 #(quan_width) VNU359 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_193_359),
	.C2V_2 (C2V_255_359),
	.C2V_3 (C2V_281_359),
	.L (L[5384:5370]),
	.V2C_1 (V2C_359_193),
	.V2C_2 (V2C_359_255),
	.V2C_3 (V2C_359_281),
	.V (V_359)
);

VNU_3 #(quan_width) VNU360 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_199_360),
	.C2V_2 (C2V_261_360),
	.C2V_3 (C2V_287_360),
	.L (L[5399:5385]),
	.V2C_1 (V2C_360_199),
	.V2C_2 (V2C_360_261),
	.V2C_3 (V2C_360_287),
	.V (V_360)
);

VNU_3 #(quan_width) VNU361 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_361),
	.C2V_2 (C2V_205_361),
	.C2V_3 (C2V_267_361),
	.L (L[5414:5400]),
	.V2C_1 (V2C_361_5),
	.V2C_2 (V2C_361_205),
	.V2C_3 (V2C_361_267),
	.V (V_361)
);

VNU_3 #(quan_width) VNU362 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_362),
	.C2V_2 (C2V_211_362),
	.C2V_3 (C2V_273_362),
	.L (L[5429:5415]),
	.V2C_1 (V2C_362_11),
	.V2C_2 (V2C_362_211),
	.V2C_3 (V2C_362_273),
	.V (V_362)
);

VNU_3 #(quan_width) VNU363 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_363),
	.C2V_2 (C2V_217_363),
	.C2V_3 (C2V_279_363),
	.L (L[5444:5430]),
	.V2C_1 (V2C_363_17),
	.V2C_2 (V2C_363_217),
	.V2C_3 (V2C_363_279),
	.V (V_363)
);

VNU_3 #(quan_width) VNU364 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_364),
	.C2V_2 (C2V_223_364),
	.C2V_3 (C2V_285_364),
	.L (L[5459:5445]),
	.V2C_1 (V2C_364_23),
	.V2C_2 (V2C_364_223),
	.V2C_3 (V2C_364_285),
	.V (V_364)
);

VNU_3 #(quan_width) VNU365 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_365),
	.C2V_2 (C2V_29_365),
	.C2V_3 (C2V_229_365),
	.L (L[5474:5460]),
	.V2C_1 (V2C_365_3),
	.V2C_2 (V2C_365_29),
	.V2C_3 (V2C_365_229),
	.V (V_365)
);

VNU_3 #(quan_width) VNU366 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_366),
	.C2V_2 (C2V_35_366),
	.C2V_3 (C2V_235_366),
	.L (L[5489:5475]),
	.V2C_1 (V2C_366_9),
	.V2C_2 (V2C_366_35),
	.V2C_3 (V2C_366_235),
	.V (V_366)
);

VNU_3 #(quan_width) VNU367 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_367),
	.C2V_2 (C2V_41_367),
	.C2V_3 (C2V_241_367),
	.L (L[5504:5490]),
	.V2C_1 (V2C_367_15),
	.V2C_2 (V2C_367_41),
	.V2C_3 (V2C_367_241),
	.V (V_367)
);

VNU_3 #(quan_width) VNU368 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_368),
	.C2V_2 (C2V_47_368),
	.C2V_3 (C2V_247_368),
	.L (L[5519:5505]),
	.V2C_1 (V2C_368_21),
	.V2C_2 (V2C_368_47),
	.V2C_3 (V2C_368_247),
	.V (V_368)
);

VNU_3 #(quan_width) VNU369 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_369),
	.C2V_2 (C2V_53_369),
	.C2V_3 (C2V_253_369),
	.L (L[5534:5520]),
	.V2C_1 (V2C_369_27),
	.V2C_2 (V2C_369_53),
	.V2C_3 (V2C_369_253),
	.V (V_369)
);

VNU_3 #(quan_width) VNU370 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_370),
	.C2V_2 (C2V_59_370),
	.C2V_3 (C2V_259_370),
	.L (L[5549:5535]),
	.V2C_1 (V2C_370_33),
	.V2C_2 (V2C_370_59),
	.V2C_3 (V2C_370_259),
	.V (V_370)
);

VNU_3 #(quan_width) VNU371 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_371),
	.C2V_2 (C2V_65_371),
	.C2V_3 (C2V_265_371),
	.L (L[5564:5550]),
	.V2C_1 (V2C_371_39),
	.V2C_2 (V2C_371_65),
	.V2C_3 (V2C_371_265),
	.V (V_371)
);

VNU_3 #(quan_width) VNU372 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_372),
	.C2V_2 (C2V_71_372),
	.C2V_3 (C2V_271_372),
	.L (L[5579:5565]),
	.V2C_1 (V2C_372_45),
	.V2C_2 (V2C_372_71),
	.V2C_3 (V2C_372_271),
	.V (V_372)
);

VNU_3 #(quan_width) VNU373 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_373),
	.C2V_2 (C2V_77_373),
	.C2V_3 (C2V_277_373),
	.L (L[5594:5580]),
	.V2C_1 (V2C_373_51),
	.V2C_2 (V2C_373_77),
	.V2C_3 (V2C_373_277),
	.V (V_373)
);

VNU_3 #(quan_width) VNU374 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_374),
	.C2V_2 (C2V_83_374),
	.C2V_3 (C2V_283_374),
	.L (L[5609:5595]),
	.V2C_1 (V2C_374_57),
	.V2C_2 (V2C_374_83),
	.V2C_3 (V2C_374_283),
	.V (V_374)
);

VNU_3 #(quan_width) VNU375 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_375),
	.C2V_2 (C2V_63_375),
	.C2V_3 (C2V_89_375),
	.L (L[5624:5610]),
	.V2C_1 (V2C_375_1),
	.V2C_2 (V2C_375_63),
	.V2C_3 (V2C_375_89),
	.V (V_375)
);

VNU_3 #(quan_width) VNU376 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_376),
	.C2V_2 (C2V_69_376),
	.C2V_3 (C2V_95_376),
	.L (L[5639:5625]),
	.V2C_1 (V2C_376_7),
	.V2C_2 (V2C_376_69),
	.V2C_3 (V2C_376_95),
	.V (V_376)
);

VNU_3 #(quan_width) VNU377 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_377),
	.C2V_2 (C2V_75_377),
	.C2V_3 (C2V_101_377),
	.L (L[5654:5640]),
	.V2C_1 (V2C_377_13),
	.V2C_2 (V2C_377_75),
	.V2C_3 (V2C_377_101),
	.V (V_377)
);

VNU_3 #(quan_width) VNU378 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_378),
	.C2V_2 (C2V_81_378),
	.C2V_3 (C2V_107_378),
	.L (L[5669:5655]),
	.V2C_1 (V2C_378_19),
	.V2C_2 (V2C_378_81),
	.V2C_3 (V2C_378_107),
	.V (V_378)
);

VNU_3 #(quan_width) VNU379 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_379),
	.C2V_2 (C2V_87_379),
	.C2V_3 (C2V_113_379),
	.L (L[5684:5670]),
	.V2C_1 (V2C_379_25),
	.V2C_2 (V2C_379_87),
	.V2C_3 (V2C_379_113),
	.V (V_379)
);

VNU_3 #(quan_width) VNU380 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_380),
	.C2V_2 (C2V_93_380),
	.C2V_3 (C2V_119_380),
	.L (L[5699:5685]),
	.V2C_1 (V2C_380_31),
	.V2C_2 (V2C_380_93),
	.V2C_3 (V2C_380_119),
	.V (V_380)
);

VNU_3 #(quan_width) VNU381 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_381),
	.C2V_2 (C2V_99_381),
	.C2V_3 (C2V_125_381),
	.L (L[5714:5700]),
	.V2C_1 (V2C_381_37),
	.V2C_2 (V2C_381_99),
	.V2C_3 (V2C_381_125),
	.V (V_381)
);

VNU_3 #(quan_width) VNU382 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_382),
	.C2V_2 (C2V_105_382),
	.C2V_3 (C2V_131_382),
	.L (L[5729:5715]),
	.V2C_1 (V2C_382_43),
	.V2C_2 (V2C_382_105),
	.V2C_3 (V2C_382_131),
	.V (V_382)
);

VNU_3 #(quan_width) VNU383 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_383),
	.C2V_2 (C2V_111_383),
	.C2V_3 (C2V_137_383),
	.L (L[5744:5730]),
	.V2C_1 (V2C_383_49),
	.V2C_2 (V2C_383_111),
	.V2C_3 (V2C_383_137),
	.V (V_383)
);

VNU_3 #(quan_width) VNU384 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_384),
	.C2V_2 (C2V_117_384),
	.C2V_3 (C2V_143_384),
	.L (L[5759:5745]),
	.V2C_1 (V2C_384_55),
	.V2C_2 (V2C_384_117),
	.V2C_3 (V2C_384_143),
	.V (V_384)
);

VNU_3 #(quan_width) VNU385 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_385),
	.C2V_2 (C2V_62_385),
	.C2V_3 (C2V_81_385),
	.L (L[5774:5760]),
	.V2C_1 (V2C_385_25),
	.V2C_2 (V2C_385_62),
	.V2C_3 (V2C_385_81),
	.V (V_385)
);

VNU_3 #(quan_width) VNU386 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_386),
	.C2V_2 (C2V_68_386),
	.C2V_3 (C2V_87_386),
	.L (L[5789:5775]),
	.V2C_1 (V2C_386_31),
	.V2C_2 (V2C_386_68),
	.V2C_3 (V2C_386_87),
	.V (V_386)
);

VNU_3 #(quan_width) VNU387 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_387),
	.C2V_2 (C2V_74_387),
	.C2V_3 (C2V_93_387),
	.L (L[5804:5790]),
	.V2C_1 (V2C_387_37),
	.V2C_2 (V2C_387_74),
	.V2C_3 (V2C_387_93),
	.V (V_387)
);

VNU_3 #(quan_width) VNU388 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_388),
	.C2V_2 (C2V_80_388),
	.C2V_3 (C2V_99_388),
	.L (L[5819:5805]),
	.V2C_1 (V2C_388_43),
	.V2C_2 (V2C_388_80),
	.V2C_3 (V2C_388_99),
	.V (V_388)
);

VNU_3 #(quan_width) VNU389 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_389),
	.C2V_2 (C2V_86_389),
	.C2V_3 (C2V_105_389),
	.L (L[5834:5820]),
	.V2C_1 (V2C_389_49),
	.V2C_2 (V2C_389_86),
	.V2C_3 (V2C_389_105),
	.V (V_389)
);

VNU_3 #(quan_width) VNU390 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_390),
	.C2V_2 (C2V_92_390),
	.C2V_3 (C2V_111_390),
	.L (L[5849:5835]),
	.V2C_1 (V2C_390_55),
	.V2C_2 (V2C_390_92),
	.V2C_3 (V2C_390_111),
	.V (V_390)
);

VNU_3 #(quan_width) VNU391 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_391),
	.C2V_2 (C2V_98_391),
	.C2V_3 (C2V_117_391),
	.L (L[5864:5850]),
	.V2C_1 (V2C_391_61),
	.V2C_2 (V2C_391_98),
	.V2C_3 (V2C_391_117),
	.V (V_391)
);

VNU_3 #(quan_width) VNU392 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_392),
	.C2V_2 (C2V_104_392),
	.C2V_3 (C2V_123_392),
	.L (L[5879:5865]),
	.V2C_1 (V2C_392_67),
	.V2C_2 (V2C_392_104),
	.V2C_3 (V2C_392_123),
	.V (V_392)
);

VNU_3 #(quan_width) VNU393 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_393),
	.C2V_2 (C2V_110_393),
	.C2V_3 (C2V_129_393),
	.L (L[5894:5880]),
	.V2C_1 (V2C_393_73),
	.V2C_2 (V2C_393_110),
	.V2C_3 (V2C_393_129),
	.V (V_393)
);

VNU_3 #(quan_width) VNU394 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_394),
	.C2V_2 (C2V_116_394),
	.C2V_3 (C2V_135_394),
	.L (L[5909:5895]),
	.V2C_1 (V2C_394_79),
	.V2C_2 (V2C_394_116),
	.V2C_3 (V2C_394_135),
	.V (V_394)
);

VNU_3 #(quan_width) VNU395 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_395),
	.C2V_2 (C2V_122_395),
	.C2V_3 (C2V_141_395),
	.L (L[5924:5910]),
	.V2C_1 (V2C_395_85),
	.V2C_2 (V2C_395_122),
	.V2C_3 (V2C_395_141),
	.V (V_395)
);

VNU_3 #(quan_width) VNU396 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_91_396),
	.C2V_2 (C2V_128_396),
	.C2V_3 (C2V_147_396),
	.L (L[5939:5925]),
	.V2C_1 (V2C_396_91),
	.V2C_2 (V2C_396_128),
	.V2C_3 (V2C_396_147),
	.V (V_396)
);

VNU_3 #(quan_width) VNU397 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_97_397),
	.C2V_2 (C2V_134_397),
	.C2V_3 (C2V_153_397),
	.L (L[5954:5940]),
	.V2C_1 (V2C_397_97),
	.V2C_2 (V2C_397_134),
	.V2C_3 (V2C_397_153),
	.V (V_397)
);

VNU_3 #(quan_width) VNU398 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_103_398),
	.C2V_2 (C2V_140_398),
	.C2V_3 (C2V_159_398),
	.L (L[5969:5955]),
	.V2C_1 (V2C_398_103),
	.V2C_2 (V2C_398_140),
	.V2C_3 (V2C_398_159),
	.V (V_398)
);

VNU_3 #(quan_width) VNU399 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_109_399),
	.C2V_2 (C2V_146_399),
	.C2V_3 (C2V_165_399),
	.L (L[5984:5970]),
	.V2C_1 (V2C_399_109),
	.V2C_2 (V2C_399_146),
	.V2C_3 (V2C_399_165),
	.V (V_399)
);

VNU_3 #(quan_width) VNU400 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_115_400),
	.C2V_2 (C2V_152_400),
	.C2V_3 (C2V_171_400),
	.L (L[5999:5985]),
	.V2C_1 (V2C_400_115),
	.V2C_2 (V2C_400_152),
	.V2C_3 (V2C_400_171),
	.V (V_400)
);

VNU_3 #(quan_width) VNU401 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_121_401),
	.C2V_2 (C2V_158_401),
	.C2V_3 (C2V_177_401),
	.L (L[6014:6000]),
	.V2C_1 (V2C_401_121),
	.V2C_2 (V2C_401_158),
	.V2C_3 (V2C_401_177),
	.V (V_401)
);

VNU_3 #(quan_width) VNU402 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_127_402),
	.C2V_2 (C2V_164_402),
	.C2V_3 (C2V_183_402),
	.L (L[6029:6015]),
	.V2C_1 (V2C_402_127),
	.V2C_2 (V2C_402_164),
	.V2C_3 (V2C_402_183),
	.V (V_402)
);

VNU_3 #(quan_width) VNU403 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_133_403),
	.C2V_2 (C2V_170_403),
	.C2V_3 (C2V_189_403),
	.L (L[6044:6030]),
	.V2C_1 (V2C_403_133),
	.V2C_2 (V2C_403_170),
	.V2C_3 (V2C_403_189),
	.V (V_403)
);

VNU_3 #(quan_width) VNU404 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_139_404),
	.C2V_2 (C2V_176_404),
	.C2V_3 (C2V_195_404),
	.L (L[6059:6045]),
	.V2C_1 (V2C_404_139),
	.V2C_2 (V2C_404_176),
	.V2C_3 (V2C_404_195),
	.V (V_404)
);

VNU_3 #(quan_width) VNU405 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_145_405),
	.C2V_2 (C2V_182_405),
	.C2V_3 (C2V_201_405),
	.L (L[6074:6060]),
	.V2C_1 (V2C_405_145),
	.V2C_2 (V2C_405_182),
	.V2C_3 (V2C_405_201),
	.V (V_405)
);

VNU_3 #(quan_width) VNU406 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_151_406),
	.C2V_2 (C2V_188_406),
	.C2V_3 (C2V_207_406),
	.L (L[6089:6075]),
	.V2C_1 (V2C_406_151),
	.V2C_2 (V2C_406_188),
	.V2C_3 (V2C_406_207),
	.V (V_406)
);

VNU_3 #(quan_width) VNU407 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_157_407),
	.C2V_2 (C2V_194_407),
	.C2V_3 (C2V_213_407),
	.L (L[6104:6090]),
	.V2C_1 (V2C_407_157),
	.V2C_2 (V2C_407_194),
	.V2C_3 (V2C_407_213),
	.V (V_407)
);

VNU_3 #(quan_width) VNU408 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_163_408),
	.C2V_2 (C2V_200_408),
	.C2V_3 (C2V_219_408),
	.L (L[6119:6105]),
	.V2C_1 (V2C_408_163),
	.V2C_2 (V2C_408_200),
	.V2C_3 (V2C_408_219),
	.V (V_408)
);

VNU_3 #(quan_width) VNU409 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_169_409),
	.C2V_2 (C2V_206_409),
	.C2V_3 (C2V_225_409),
	.L (L[6134:6120]),
	.V2C_1 (V2C_409_169),
	.V2C_2 (V2C_409_206),
	.V2C_3 (V2C_409_225),
	.V (V_409)
);

VNU_3 #(quan_width) VNU410 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_175_410),
	.C2V_2 (C2V_212_410),
	.C2V_3 (C2V_231_410),
	.L (L[6149:6135]),
	.V2C_1 (V2C_410_175),
	.V2C_2 (V2C_410_212),
	.V2C_3 (V2C_410_231),
	.V (V_410)
);

VNU_3 #(quan_width) VNU411 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_181_411),
	.C2V_2 (C2V_218_411),
	.C2V_3 (C2V_237_411),
	.L (L[6164:6150]),
	.V2C_1 (V2C_411_181),
	.V2C_2 (V2C_411_218),
	.V2C_3 (V2C_411_237),
	.V (V_411)
);

VNU_3 #(quan_width) VNU412 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_187_412),
	.C2V_2 (C2V_224_412),
	.C2V_3 (C2V_243_412),
	.L (L[6179:6165]),
	.V2C_1 (V2C_412_187),
	.V2C_2 (V2C_412_224),
	.V2C_3 (V2C_412_243),
	.V (V_412)
);

VNU_3 #(quan_width) VNU413 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_193_413),
	.C2V_2 (C2V_230_413),
	.C2V_3 (C2V_249_413),
	.L (L[6194:6180]),
	.V2C_1 (V2C_413_193),
	.V2C_2 (V2C_413_230),
	.V2C_3 (V2C_413_249),
	.V (V_413)
);

VNU_3 #(quan_width) VNU414 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_199_414),
	.C2V_2 (C2V_236_414),
	.C2V_3 (C2V_255_414),
	.L (L[6209:6195]),
	.V2C_1 (V2C_414_199),
	.V2C_2 (V2C_414_236),
	.V2C_3 (V2C_414_255),
	.V (V_414)
);

VNU_3 #(quan_width) VNU415 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_205_415),
	.C2V_2 (C2V_242_415),
	.C2V_3 (C2V_261_415),
	.L (L[6224:6210]),
	.V2C_1 (V2C_415_205),
	.V2C_2 (V2C_415_242),
	.V2C_3 (V2C_415_261),
	.V (V_415)
);

VNU_3 #(quan_width) VNU416 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_211_416),
	.C2V_2 (C2V_248_416),
	.C2V_3 (C2V_267_416),
	.L (L[6239:6225]),
	.V2C_1 (V2C_416_211),
	.V2C_2 (V2C_416_248),
	.V2C_3 (V2C_416_267),
	.V (V_416)
);

VNU_3 #(quan_width) VNU417 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_217_417),
	.C2V_2 (C2V_254_417),
	.C2V_3 (C2V_273_417),
	.L (L[6254:6240]),
	.V2C_1 (V2C_417_217),
	.V2C_2 (V2C_417_254),
	.V2C_3 (V2C_417_273),
	.V (V_417)
);

VNU_3 #(quan_width) VNU418 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_223_418),
	.C2V_2 (C2V_260_418),
	.C2V_3 (C2V_279_418),
	.L (L[6269:6255]),
	.V2C_1 (V2C_418_223),
	.V2C_2 (V2C_418_260),
	.V2C_3 (V2C_418_279),
	.V (V_418)
);

VNU_3 #(quan_width) VNU419 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_229_419),
	.C2V_2 (C2V_266_419),
	.C2V_3 (C2V_285_419),
	.L (L[6284:6270]),
	.V2C_1 (V2C_419_229),
	.V2C_2 (V2C_419_266),
	.V2C_3 (V2C_419_285),
	.V (V_419)
);

VNU_3 #(quan_width) VNU420 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_420),
	.C2V_2 (C2V_235_420),
	.C2V_3 (C2V_272_420),
	.L (L[6299:6285]),
	.V2C_1 (V2C_420_3),
	.V2C_2 (V2C_420_235),
	.V2C_3 (V2C_420_272),
	.V (V_420)
);

VNU_3 #(quan_width) VNU421 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_421),
	.C2V_2 (C2V_241_421),
	.C2V_3 (C2V_278_421),
	.L (L[6314:6300]),
	.V2C_1 (V2C_421_9),
	.V2C_2 (V2C_421_241),
	.V2C_3 (V2C_421_278),
	.V (V_421)
);

VNU_3 #(quan_width) VNU422 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_422),
	.C2V_2 (C2V_247_422),
	.C2V_3 (C2V_284_422),
	.L (L[6329:6315]),
	.V2C_1 (V2C_422_15),
	.V2C_2 (V2C_422_247),
	.V2C_3 (V2C_422_284),
	.V (V_422)
);

VNU_3 #(quan_width) VNU423 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_423),
	.C2V_2 (C2V_21_423),
	.C2V_3 (C2V_253_423),
	.L (L[6344:6330]),
	.V2C_1 (V2C_423_2),
	.V2C_2 (V2C_423_21),
	.V2C_3 (V2C_423_253),
	.V (V_423)
);

VNU_3 #(quan_width) VNU424 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_424),
	.C2V_2 (C2V_27_424),
	.C2V_3 (C2V_259_424),
	.L (L[6359:6345]),
	.V2C_1 (V2C_424_8),
	.V2C_2 (V2C_424_27),
	.V2C_3 (V2C_424_259),
	.V (V_424)
);

VNU_3 #(quan_width) VNU425 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_425),
	.C2V_2 (C2V_33_425),
	.C2V_3 (C2V_265_425),
	.L (L[6374:6360]),
	.V2C_1 (V2C_425_14),
	.V2C_2 (V2C_425_33),
	.V2C_3 (V2C_425_265),
	.V (V_425)
);

VNU_3 #(quan_width) VNU426 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_426),
	.C2V_2 (C2V_39_426),
	.C2V_3 (C2V_271_426),
	.L (L[6389:6375]),
	.V2C_1 (V2C_426_20),
	.V2C_2 (V2C_426_39),
	.V2C_3 (V2C_426_271),
	.V (V_426)
);

VNU_3 #(quan_width) VNU427 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_427),
	.C2V_2 (C2V_45_427),
	.C2V_3 (C2V_277_427),
	.L (L[6404:6390]),
	.V2C_1 (V2C_427_26),
	.V2C_2 (V2C_427_45),
	.V2C_3 (V2C_427_277),
	.V (V_427)
);

VNU_3 #(quan_width) VNU428 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_428),
	.C2V_2 (C2V_51_428),
	.C2V_3 (C2V_283_428),
	.L (L[6419:6405]),
	.V2C_1 (V2C_428_32),
	.V2C_2 (V2C_428_51),
	.V2C_3 (V2C_428_283),
	.V (V_428)
);

VNU_3 #(quan_width) VNU429 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_429),
	.C2V_2 (C2V_38_429),
	.C2V_3 (C2V_57_429),
	.L (L[6434:6420]),
	.V2C_1 (V2C_429_1),
	.V2C_2 (V2C_429_38),
	.V2C_3 (V2C_429_57),
	.V (V_429)
);

VNU_3 #(quan_width) VNU430 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_430),
	.C2V_2 (C2V_44_430),
	.C2V_3 (C2V_63_430),
	.L (L[6449:6435]),
	.V2C_1 (V2C_430_7),
	.V2C_2 (V2C_430_44),
	.V2C_3 (V2C_430_63),
	.V (V_430)
);

VNU_3 #(quan_width) VNU431 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_431),
	.C2V_2 (C2V_50_431),
	.C2V_3 (C2V_69_431),
	.L (L[6464:6450]),
	.V2C_1 (V2C_431_13),
	.V2C_2 (V2C_431_50),
	.V2C_3 (V2C_431_69),
	.V (V_431)
);

VNU_3 #(quan_width) VNU432 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_432),
	.C2V_2 (C2V_56_432),
	.C2V_3 (C2V_75_432),
	.L (L[6479:6465]),
	.V2C_1 (V2C_432_19),
	.V2C_2 (V2C_432_56),
	.V2C_3 (V2C_432_75),
	.V (V_432)
);

VNU_3 #(quan_width) VNU433 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_433),
	.C2V_2 (C2V_28_433),
	.C2V_3 (C2V_251_433),
	.L (L[6494:6480]),
	.V2C_1 (V2C_433_12),
	.V2C_2 (V2C_433_28),
	.V2C_3 (V2C_433_251),
	.V (V_433)
);

VNU_3 #(quan_width) VNU434 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_434),
	.C2V_2 (C2V_34_434),
	.C2V_3 (C2V_257_434),
	.L (L[6509:6495]),
	.V2C_1 (V2C_434_18),
	.V2C_2 (V2C_434_34),
	.V2C_3 (V2C_434_257),
	.V (V_434)
);

VNU_3 #(quan_width) VNU435 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_435),
	.C2V_2 (C2V_40_435),
	.C2V_3 (C2V_263_435),
	.L (L[6524:6510]),
	.V2C_1 (V2C_435_24),
	.V2C_2 (V2C_435_40),
	.V2C_3 (V2C_435_263),
	.V (V_435)
);

VNU_3 #(quan_width) VNU436 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_436),
	.C2V_2 (C2V_46_436),
	.C2V_3 (C2V_269_436),
	.L (L[6539:6525]),
	.V2C_1 (V2C_436_30),
	.V2C_2 (V2C_436_46),
	.V2C_3 (V2C_436_269),
	.V (V_436)
);

VNU_3 #(quan_width) VNU437 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_437),
	.C2V_2 (C2V_52_437),
	.C2V_3 (C2V_275_437),
	.L (L[6554:6540]),
	.V2C_1 (V2C_437_36),
	.V2C_2 (V2C_437_52),
	.V2C_3 (V2C_437_275),
	.V (V_437)
);

VNU_3 #(quan_width) VNU438 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_438),
	.C2V_2 (C2V_58_438),
	.C2V_3 (C2V_281_438),
	.L (L[6569:6555]),
	.V2C_1 (V2C_438_42),
	.V2C_2 (V2C_438_58),
	.V2C_3 (V2C_438_281),
	.V (V_438)
);

VNU_3 #(quan_width) VNU439 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_439),
	.C2V_2 (C2V_64_439),
	.C2V_3 (C2V_287_439),
	.L (L[6584:6570]),
	.V2C_1 (V2C_439_48),
	.V2C_2 (V2C_439_64),
	.V2C_3 (V2C_439_287),
	.V (V_439)
);

VNU_3 #(quan_width) VNU440 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_440),
	.C2V_2 (C2V_54_440),
	.C2V_3 (C2V_70_440),
	.L (L[6599:6585]),
	.V2C_1 (V2C_440_5),
	.V2C_2 (V2C_440_54),
	.V2C_3 (V2C_440_70),
	.V (V_440)
);

VNU_3 #(quan_width) VNU441 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_441),
	.C2V_2 (C2V_60_441),
	.C2V_3 (C2V_76_441),
	.L (L[6614:6600]),
	.V2C_1 (V2C_441_11),
	.V2C_2 (V2C_441_60),
	.V2C_3 (V2C_441_76),
	.V (V_441)
);

VNU_3 #(quan_width) VNU442 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_442),
	.C2V_2 (C2V_66_442),
	.C2V_3 (C2V_82_442),
	.L (L[6629:6615]),
	.V2C_1 (V2C_442_17),
	.V2C_2 (V2C_442_66),
	.V2C_3 (V2C_442_82),
	.V (V_442)
);

VNU_3 #(quan_width) VNU443 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_443),
	.C2V_2 (C2V_72_443),
	.C2V_3 (C2V_88_443),
	.L (L[6644:6630]),
	.V2C_1 (V2C_443_23),
	.V2C_2 (V2C_443_72),
	.V2C_3 (V2C_443_88),
	.V (V_443)
);

VNU_3 #(quan_width) VNU444 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_444),
	.C2V_2 (C2V_78_444),
	.C2V_3 (C2V_94_444),
	.L (L[6659:6645]),
	.V2C_1 (V2C_444_29),
	.V2C_2 (V2C_444_78),
	.V2C_3 (V2C_444_94),
	.V (V_444)
);

VNU_3 #(quan_width) VNU445 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_445),
	.C2V_2 (C2V_84_445),
	.C2V_3 (C2V_100_445),
	.L (L[6674:6660]),
	.V2C_1 (V2C_445_35),
	.V2C_2 (V2C_445_84),
	.V2C_3 (V2C_445_100),
	.V (V_445)
);

VNU_3 #(quan_width) VNU446 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_446),
	.C2V_2 (C2V_90_446),
	.C2V_3 (C2V_106_446),
	.L (L[6689:6675]),
	.V2C_1 (V2C_446_41),
	.V2C_2 (V2C_446_90),
	.V2C_3 (V2C_446_106),
	.V (V_446)
);

VNU_3 #(quan_width) VNU447 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_447),
	.C2V_2 (C2V_96_447),
	.C2V_3 (C2V_112_447),
	.L (L[6704:6690]),
	.V2C_1 (V2C_447_47),
	.V2C_2 (V2C_447_96),
	.V2C_3 (V2C_447_112),
	.V (V_447)
);

VNU_3 #(quan_width) VNU448 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_448),
	.C2V_2 (C2V_102_448),
	.C2V_3 (C2V_118_448),
	.L (L[6719:6705]),
	.V2C_1 (V2C_448_53),
	.V2C_2 (V2C_448_102),
	.V2C_3 (V2C_448_118),
	.V (V_448)
);

VNU_3 #(quan_width) VNU449 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_59_449),
	.C2V_2 (C2V_108_449),
	.C2V_3 (C2V_124_449),
	.L (L[6734:6720]),
	.V2C_1 (V2C_449_59),
	.V2C_2 (V2C_449_108),
	.V2C_3 (V2C_449_124),
	.V (V_449)
);

VNU_3 #(quan_width) VNU450 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_65_450),
	.C2V_2 (C2V_114_450),
	.C2V_3 (C2V_130_450),
	.L (L[6749:6735]),
	.V2C_1 (V2C_450_65),
	.V2C_2 (V2C_450_114),
	.V2C_3 (V2C_450_130),
	.V (V_450)
);

VNU_3 #(quan_width) VNU451 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_71_451),
	.C2V_2 (C2V_120_451),
	.C2V_3 (C2V_136_451),
	.L (L[6764:6750]),
	.V2C_1 (V2C_451_71),
	.V2C_2 (V2C_451_120),
	.V2C_3 (V2C_451_136),
	.V (V_451)
);

VNU_3 #(quan_width) VNU452 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_77_452),
	.C2V_2 (C2V_126_452),
	.C2V_3 (C2V_142_452),
	.L (L[6779:6765]),
	.V2C_1 (V2C_452_77),
	.V2C_2 (V2C_452_126),
	.V2C_3 (V2C_452_142),
	.V (V_452)
);

VNU_3 #(quan_width) VNU453 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_83_453),
	.C2V_2 (C2V_132_453),
	.C2V_3 (C2V_148_453),
	.L (L[6794:6780]),
	.V2C_1 (V2C_453_83),
	.V2C_2 (V2C_453_132),
	.V2C_3 (V2C_453_148),
	.V (V_453)
);

VNU_3 #(quan_width) VNU454 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_89_454),
	.C2V_2 (C2V_138_454),
	.C2V_3 (C2V_154_454),
	.L (L[6809:6795]),
	.V2C_1 (V2C_454_89),
	.V2C_2 (V2C_454_138),
	.V2C_3 (V2C_454_154),
	.V (V_454)
);

VNU_3 #(quan_width) VNU455 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_95_455),
	.C2V_2 (C2V_144_455),
	.C2V_3 (C2V_160_455),
	.L (L[6824:6810]),
	.V2C_1 (V2C_455_95),
	.V2C_2 (V2C_455_144),
	.V2C_3 (V2C_455_160),
	.V (V_455)
);

VNU_3 #(quan_width) VNU456 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_101_456),
	.C2V_2 (C2V_150_456),
	.C2V_3 (C2V_166_456),
	.L (L[6839:6825]),
	.V2C_1 (V2C_456_101),
	.V2C_2 (V2C_456_150),
	.V2C_3 (V2C_456_166),
	.V (V_456)
);

VNU_3 #(quan_width) VNU457 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_107_457),
	.C2V_2 (C2V_156_457),
	.C2V_3 (C2V_172_457),
	.L (L[6854:6840]),
	.V2C_1 (V2C_457_107),
	.V2C_2 (V2C_457_156),
	.V2C_3 (V2C_457_172),
	.V (V_457)
);

VNU_3 #(quan_width) VNU458 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_113_458),
	.C2V_2 (C2V_162_458),
	.C2V_3 (C2V_178_458),
	.L (L[6869:6855]),
	.V2C_1 (V2C_458_113),
	.V2C_2 (V2C_458_162),
	.V2C_3 (V2C_458_178),
	.V (V_458)
);

VNU_3 #(quan_width) VNU459 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_119_459),
	.C2V_2 (C2V_168_459),
	.C2V_3 (C2V_184_459),
	.L (L[6884:6870]),
	.V2C_1 (V2C_459_119),
	.V2C_2 (V2C_459_168),
	.V2C_3 (V2C_459_184),
	.V (V_459)
);

VNU_3 #(quan_width) VNU460 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_125_460),
	.C2V_2 (C2V_174_460),
	.C2V_3 (C2V_190_460),
	.L (L[6899:6885]),
	.V2C_1 (V2C_460_125),
	.V2C_2 (V2C_460_174),
	.V2C_3 (V2C_460_190),
	.V (V_460)
);

VNU_3 #(quan_width) VNU461 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_131_461),
	.C2V_2 (C2V_180_461),
	.C2V_3 (C2V_196_461),
	.L (L[6914:6900]),
	.V2C_1 (V2C_461_131),
	.V2C_2 (V2C_461_180),
	.V2C_3 (V2C_461_196),
	.V (V_461)
);

VNU_3 #(quan_width) VNU462 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_137_462),
	.C2V_2 (C2V_186_462),
	.C2V_3 (C2V_202_462),
	.L (L[6929:6915]),
	.V2C_1 (V2C_462_137),
	.V2C_2 (V2C_462_186),
	.V2C_3 (V2C_462_202),
	.V (V_462)
);

VNU_3 #(quan_width) VNU463 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_143_463),
	.C2V_2 (C2V_192_463),
	.C2V_3 (C2V_208_463),
	.L (L[6944:6930]),
	.V2C_1 (V2C_463_143),
	.V2C_2 (V2C_463_192),
	.V2C_3 (V2C_463_208),
	.V (V_463)
);

VNU_3 #(quan_width) VNU464 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_149_464),
	.C2V_2 (C2V_198_464),
	.C2V_3 (C2V_214_464),
	.L (L[6959:6945]),
	.V2C_1 (V2C_464_149),
	.V2C_2 (V2C_464_198),
	.V2C_3 (V2C_464_214),
	.V (V_464)
);

VNU_3 #(quan_width) VNU465 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_155_465),
	.C2V_2 (C2V_204_465),
	.C2V_3 (C2V_220_465),
	.L (L[6974:6960]),
	.V2C_1 (V2C_465_155),
	.V2C_2 (V2C_465_204),
	.V2C_3 (V2C_465_220),
	.V (V_465)
);

VNU_3 #(quan_width) VNU466 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_161_466),
	.C2V_2 (C2V_210_466),
	.C2V_3 (C2V_226_466),
	.L (L[6989:6975]),
	.V2C_1 (V2C_466_161),
	.V2C_2 (V2C_466_210),
	.V2C_3 (V2C_466_226),
	.V (V_466)
);

VNU_3 #(quan_width) VNU467 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_167_467),
	.C2V_2 (C2V_216_467),
	.C2V_3 (C2V_232_467),
	.L (L[7004:6990]),
	.V2C_1 (V2C_467_167),
	.V2C_2 (V2C_467_216),
	.V2C_3 (V2C_467_232),
	.V (V_467)
);

VNU_3 #(quan_width) VNU468 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_173_468),
	.C2V_2 (C2V_222_468),
	.C2V_3 (C2V_238_468),
	.L (L[7019:7005]),
	.V2C_1 (V2C_468_173),
	.V2C_2 (V2C_468_222),
	.V2C_3 (V2C_468_238),
	.V (V_468)
);

VNU_3 #(quan_width) VNU469 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_179_469),
	.C2V_2 (C2V_228_469),
	.C2V_3 (C2V_244_469),
	.L (L[7034:7020]),
	.V2C_1 (V2C_469_179),
	.V2C_2 (V2C_469_228),
	.V2C_3 (V2C_469_244),
	.V (V_469)
);

VNU_3 #(quan_width) VNU470 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_185_470),
	.C2V_2 (C2V_234_470),
	.C2V_3 (C2V_250_470),
	.L (L[7049:7035]),
	.V2C_1 (V2C_470_185),
	.V2C_2 (V2C_470_234),
	.V2C_3 (V2C_470_250),
	.V (V_470)
);

VNU_3 #(quan_width) VNU471 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_191_471),
	.C2V_2 (C2V_240_471),
	.C2V_3 (C2V_256_471),
	.L (L[7064:7050]),
	.V2C_1 (V2C_471_191),
	.V2C_2 (V2C_471_240),
	.V2C_3 (V2C_471_256),
	.V (V_471)
);

VNU_3 #(quan_width) VNU472 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_197_472),
	.C2V_2 (C2V_246_472),
	.C2V_3 (C2V_262_472),
	.L (L[7079:7065]),
	.V2C_1 (V2C_472_197),
	.V2C_2 (V2C_472_246),
	.V2C_3 (V2C_472_262),
	.V (V_472)
);

VNU_3 #(quan_width) VNU473 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_203_473),
	.C2V_2 (C2V_252_473),
	.C2V_3 (C2V_268_473),
	.L (L[7094:7080]),
	.V2C_1 (V2C_473_203),
	.V2C_2 (V2C_473_252),
	.V2C_3 (V2C_473_268),
	.V (V_473)
);

VNU_3 #(quan_width) VNU474 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_209_474),
	.C2V_2 (C2V_258_474),
	.C2V_3 (C2V_274_474),
	.L (L[7109:7095]),
	.V2C_1 (V2C_474_209),
	.V2C_2 (V2C_474_258),
	.V2C_3 (V2C_474_274),
	.V (V_474)
);

VNU_3 #(quan_width) VNU475 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_215_475),
	.C2V_2 (C2V_264_475),
	.C2V_3 (C2V_280_475),
	.L (L[7124:7110]),
	.V2C_1 (V2C_475_215),
	.V2C_2 (V2C_475_264),
	.V2C_3 (V2C_475_280),
	.V (V_475)
);

VNU_3 #(quan_width) VNU476 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_221_476),
	.C2V_2 (C2V_270_476),
	.C2V_3 (C2V_286_476),
	.L (L[7139:7125]),
	.V2C_1 (V2C_476_221),
	.V2C_2 (V2C_476_270),
	.V2C_3 (V2C_476_286),
	.V (V_476)
);

VNU_3 #(quan_width) VNU477 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_477),
	.C2V_2 (C2V_227_477),
	.C2V_3 (C2V_276_477),
	.L (L[7154:7140]),
	.V2C_1 (V2C_477_4),
	.V2C_2 (V2C_477_227),
	.V2C_3 (V2C_477_276),
	.V (V_477)
);

VNU_3 #(quan_width) VNU478 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_478),
	.C2V_2 (C2V_233_478),
	.C2V_3 (C2V_282_478),
	.L (L[7169:7155]),
	.V2C_1 (V2C_478_10),
	.V2C_2 (V2C_478_233),
	.V2C_3 (V2C_478_282),
	.V (V_478)
);

VNU_3 #(quan_width) VNU479 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_479),
	.C2V_2 (C2V_239_479),
	.C2V_3 (C2V_288_479),
	.L (L[7184:7170]),
	.V2C_1 (V2C_479_16),
	.V2C_2 (V2C_479_239),
	.V2C_3 (V2C_479_288),
	.V (V_479)
);

VNU_3 #(quan_width) VNU480 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_480),
	.C2V_2 (C2V_22_480),
	.C2V_3 (C2V_245_480),
	.L (L[7199:7185]),
	.V2C_1 (V2C_480_6),
	.V2C_2 (V2C_480_22),
	.V2C_3 (V2C_480_245),
	.V (V_480)
);

VNU_3 #(quan_width) VNU481 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_481),
	.C2V_2 (C2V_76_481),
	.C2V_3 (C2V_104_481),
	.L (L[7214:7200]),
	.V2C_1 (V2C_481_19),
	.V2C_2 (V2C_481_76),
	.V2C_3 (V2C_481_104),
	.V (V_481)
);

VNU_3 #(quan_width) VNU482 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_482),
	.C2V_2 (C2V_82_482),
	.C2V_3 (C2V_110_482),
	.L (L[7229:7215]),
	.V2C_1 (V2C_482_25),
	.V2C_2 (V2C_482_82),
	.V2C_3 (V2C_482_110),
	.V (V_482)
);

VNU_3 #(quan_width) VNU483 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_483),
	.C2V_2 (C2V_88_483),
	.C2V_3 (C2V_116_483),
	.L (L[7244:7230]),
	.V2C_1 (V2C_483_31),
	.V2C_2 (V2C_483_88),
	.V2C_3 (V2C_483_116),
	.V (V_483)
);

VNU_3 #(quan_width) VNU484 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_484),
	.C2V_2 (C2V_94_484),
	.C2V_3 (C2V_122_484),
	.L (L[7259:7245]),
	.V2C_1 (V2C_484_37),
	.V2C_2 (V2C_484_94),
	.V2C_3 (V2C_484_122),
	.V (V_484)
);

VNU_3 #(quan_width) VNU485 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_485),
	.C2V_2 (C2V_100_485),
	.C2V_3 (C2V_128_485),
	.L (L[7274:7260]),
	.V2C_1 (V2C_485_43),
	.V2C_2 (V2C_485_100),
	.V2C_3 (V2C_485_128),
	.V (V_485)
);

VNU_3 #(quan_width) VNU486 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_486),
	.C2V_2 (C2V_106_486),
	.C2V_3 (C2V_134_486),
	.L (L[7289:7275]),
	.V2C_1 (V2C_486_49),
	.V2C_2 (V2C_486_106),
	.V2C_3 (V2C_486_134),
	.V (V_486)
);

VNU_3 #(quan_width) VNU487 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_487),
	.C2V_2 (C2V_112_487),
	.C2V_3 (C2V_140_487),
	.L (L[7304:7290]),
	.V2C_1 (V2C_487_55),
	.V2C_2 (V2C_487_112),
	.V2C_3 (V2C_487_140),
	.V (V_487)
);

VNU_3 #(quan_width) VNU488 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_488),
	.C2V_2 (C2V_118_488),
	.C2V_3 (C2V_146_488),
	.L (L[7319:7305]),
	.V2C_1 (V2C_488_61),
	.V2C_2 (V2C_488_118),
	.V2C_3 (V2C_488_146),
	.V (V_488)
);

VNU_3 #(quan_width) VNU489 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_489),
	.C2V_2 (C2V_124_489),
	.C2V_3 (C2V_152_489),
	.L (L[7334:7320]),
	.V2C_1 (V2C_489_67),
	.V2C_2 (V2C_489_124),
	.V2C_3 (V2C_489_152),
	.V (V_489)
);

VNU_3 #(quan_width) VNU490 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_490),
	.C2V_2 (C2V_130_490),
	.C2V_3 (C2V_158_490),
	.L (L[7349:7335]),
	.V2C_1 (V2C_490_73),
	.V2C_2 (V2C_490_130),
	.V2C_3 (V2C_490_158),
	.V (V_490)
);

VNU_3 #(quan_width) VNU491 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_491),
	.C2V_2 (C2V_136_491),
	.C2V_3 (C2V_164_491),
	.L (L[7364:7350]),
	.V2C_1 (V2C_491_79),
	.V2C_2 (V2C_491_136),
	.V2C_3 (V2C_491_164),
	.V (V_491)
);

VNU_3 #(quan_width) VNU492 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_492),
	.C2V_2 (C2V_142_492),
	.C2V_3 (C2V_170_492),
	.L (L[7379:7365]),
	.V2C_1 (V2C_492_85),
	.V2C_2 (V2C_492_142),
	.V2C_3 (V2C_492_170),
	.V (V_492)
);

VNU_3 #(quan_width) VNU493 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_91_493),
	.C2V_2 (C2V_148_493),
	.C2V_3 (C2V_176_493),
	.L (L[7394:7380]),
	.V2C_1 (V2C_493_91),
	.V2C_2 (V2C_493_148),
	.V2C_3 (V2C_493_176),
	.V (V_493)
);

VNU_3 #(quan_width) VNU494 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_97_494),
	.C2V_2 (C2V_154_494),
	.C2V_3 (C2V_182_494),
	.L (L[7409:7395]),
	.V2C_1 (V2C_494_97),
	.V2C_2 (V2C_494_154),
	.V2C_3 (V2C_494_182),
	.V (V_494)
);

VNU_3 #(quan_width) VNU495 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_103_495),
	.C2V_2 (C2V_160_495),
	.C2V_3 (C2V_188_495),
	.L (L[7424:7410]),
	.V2C_1 (V2C_495_103),
	.V2C_2 (V2C_495_160),
	.V2C_3 (V2C_495_188),
	.V (V_495)
);

VNU_3 #(quan_width) VNU496 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_109_496),
	.C2V_2 (C2V_166_496),
	.C2V_3 (C2V_194_496),
	.L (L[7439:7425]),
	.V2C_1 (V2C_496_109),
	.V2C_2 (V2C_496_166),
	.V2C_3 (V2C_496_194),
	.V (V_496)
);

VNU_3 #(quan_width) VNU497 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_115_497),
	.C2V_2 (C2V_172_497),
	.C2V_3 (C2V_200_497),
	.L (L[7454:7440]),
	.V2C_1 (V2C_497_115),
	.V2C_2 (V2C_497_172),
	.V2C_3 (V2C_497_200),
	.V (V_497)
);

VNU_3 #(quan_width) VNU498 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_121_498),
	.C2V_2 (C2V_178_498),
	.C2V_3 (C2V_206_498),
	.L (L[7469:7455]),
	.V2C_1 (V2C_498_121),
	.V2C_2 (V2C_498_178),
	.V2C_3 (V2C_498_206),
	.V (V_498)
);

VNU_3 #(quan_width) VNU499 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_127_499),
	.C2V_2 (C2V_184_499),
	.C2V_3 (C2V_212_499),
	.L (L[7484:7470]),
	.V2C_1 (V2C_499_127),
	.V2C_2 (V2C_499_184),
	.V2C_3 (V2C_499_212),
	.V (V_499)
);

VNU_3 #(quan_width) VNU500 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_133_500),
	.C2V_2 (C2V_190_500),
	.C2V_3 (C2V_218_500),
	.L (L[7499:7485]),
	.V2C_1 (V2C_500_133),
	.V2C_2 (V2C_500_190),
	.V2C_3 (V2C_500_218),
	.V (V_500)
);

VNU_3 #(quan_width) VNU501 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_139_501),
	.C2V_2 (C2V_196_501),
	.C2V_3 (C2V_224_501),
	.L (L[7514:7500]),
	.V2C_1 (V2C_501_139),
	.V2C_2 (V2C_501_196),
	.V2C_3 (V2C_501_224),
	.V (V_501)
);

VNU_3 #(quan_width) VNU502 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_145_502),
	.C2V_2 (C2V_202_502),
	.C2V_3 (C2V_230_502),
	.L (L[7529:7515]),
	.V2C_1 (V2C_502_145),
	.V2C_2 (V2C_502_202),
	.V2C_3 (V2C_502_230),
	.V (V_502)
);

VNU_3 #(quan_width) VNU503 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_151_503),
	.C2V_2 (C2V_208_503),
	.C2V_3 (C2V_236_503),
	.L (L[7544:7530]),
	.V2C_1 (V2C_503_151),
	.V2C_2 (V2C_503_208),
	.V2C_3 (V2C_503_236),
	.V (V_503)
);

VNU_3 #(quan_width) VNU504 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_157_504),
	.C2V_2 (C2V_214_504),
	.C2V_3 (C2V_242_504),
	.L (L[7559:7545]),
	.V2C_1 (V2C_504_157),
	.V2C_2 (V2C_504_214),
	.V2C_3 (V2C_504_242),
	.V (V_504)
);

VNU_3 #(quan_width) VNU505 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_163_505),
	.C2V_2 (C2V_220_505),
	.C2V_3 (C2V_248_505),
	.L (L[7574:7560]),
	.V2C_1 (V2C_505_163),
	.V2C_2 (V2C_505_220),
	.V2C_3 (V2C_505_248),
	.V (V_505)
);

VNU_3 #(quan_width) VNU506 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_169_506),
	.C2V_2 (C2V_226_506),
	.C2V_3 (C2V_254_506),
	.L (L[7589:7575]),
	.V2C_1 (V2C_506_169),
	.V2C_2 (V2C_506_226),
	.V2C_3 (V2C_506_254),
	.V (V_506)
);

VNU_3 #(quan_width) VNU507 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_175_507),
	.C2V_2 (C2V_232_507),
	.C2V_3 (C2V_260_507),
	.L (L[7604:7590]),
	.V2C_1 (V2C_507_175),
	.V2C_2 (V2C_507_232),
	.V2C_3 (V2C_507_260),
	.V (V_507)
);

VNU_3 #(quan_width) VNU508 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_181_508),
	.C2V_2 (C2V_238_508),
	.C2V_3 (C2V_266_508),
	.L (L[7619:7605]),
	.V2C_1 (V2C_508_181),
	.V2C_2 (V2C_508_238),
	.V2C_3 (V2C_508_266),
	.V (V_508)
);

VNU_3 #(quan_width) VNU509 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_187_509),
	.C2V_2 (C2V_244_509),
	.C2V_3 (C2V_272_509),
	.L (L[7634:7620]),
	.V2C_1 (V2C_509_187),
	.V2C_2 (V2C_509_244),
	.V2C_3 (V2C_509_272),
	.V (V_509)
);

VNU_3 #(quan_width) VNU510 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_193_510),
	.C2V_2 (C2V_250_510),
	.C2V_3 (C2V_278_510),
	.L (L[7649:7635]),
	.V2C_1 (V2C_510_193),
	.V2C_2 (V2C_510_250),
	.V2C_3 (V2C_510_278),
	.V (V_510)
);

VNU_3 #(quan_width) VNU511 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_199_511),
	.C2V_2 (C2V_256_511),
	.C2V_3 (C2V_284_511),
	.L (L[7664:7650]),
	.V2C_1 (V2C_511_199),
	.V2C_2 (V2C_511_256),
	.V2C_3 (V2C_511_284),
	.V (V_511)
);

VNU_3 #(quan_width) VNU512 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_512),
	.C2V_2 (C2V_205_512),
	.C2V_3 (C2V_262_512),
	.L (L[7679:7665]),
	.V2C_1 (V2C_512_2),
	.V2C_2 (V2C_512_205),
	.V2C_3 (V2C_512_262),
	.V (V_512)
);

VNU_3 #(quan_width) VNU513 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_513),
	.C2V_2 (C2V_211_513),
	.C2V_3 (C2V_268_513),
	.L (L[7694:7680]),
	.V2C_1 (V2C_513_8),
	.V2C_2 (V2C_513_211),
	.V2C_3 (V2C_513_268),
	.V (V_513)
);

VNU_3 #(quan_width) VNU514 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_514),
	.C2V_2 (C2V_217_514),
	.C2V_3 (C2V_274_514),
	.L (L[7709:7695]),
	.V2C_1 (V2C_514_14),
	.V2C_2 (V2C_514_217),
	.V2C_3 (V2C_514_274),
	.V (V_514)
);

VNU_3 #(quan_width) VNU515 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_515),
	.C2V_2 (C2V_223_515),
	.C2V_3 (C2V_280_515),
	.L (L[7724:7710]),
	.V2C_1 (V2C_515_20),
	.V2C_2 (V2C_515_223),
	.V2C_3 (V2C_515_280),
	.V (V_515)
);

VNU_3 #(quan_width) VNU516 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_516),
	.C2V_2 (C2V_229_516),
	.C2V_3 (C2V_286_516),
	.L (L[7739:7725]),
	.V2C_1 (V2C_516_26),
	.V2C_2 (V2C_516_229),
	.V2C_3 (V2C_516_286),
	.V (V_516)
);

VNU_3 #(quan_width) VNU517 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_517),
	.C2V_2 (C2V_32_517),
	.C2V_3 (C2V_235_517),
	.L (L[7754:7740]),
	.V2C_1 (V2C_517_4),
	.V2C_2 (V2C_517_32),
	.V2C_3 (V2C_517_235),
	.V (V_517)
);

VNU_3 #(quan_width) VNU518 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_518),
	.C2V_2 (C2V_38_518),
	.C2V_3 (C2V_241_518),
	.L (L[7769:7755]),
	.V2C_1 (V2C_518_10),
	.V2C_2 (V2C_518_38),
	.V2C_3 (V2C_518_241),
	.V (V_518)
);

VNU_3 #(quan_width) VNU519 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_519),
	.C2V_2 (C2V_44_519),
	.C2V_3 (C2V_247_519),
	.L (L[7784:7770]),
	.V2C_1 (V2C_519_16),
	.V2C_2 (V2C_519_44),
	.V2C_3 (V2C_519_247),
	.V (V_519)
);

VNU_3 #(quan_width) VNU520 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_520),
	.C2V_2 (C2V_50_520),
	.C2V_3 (C2V_253_520),
	.L (L[7799:7785]),
	.V2C_1 (V2C_520_22),
	.V2C_2 (V2C_520_50),
	.V2C_3 (V2C_520_253),
	.V (V_520)
);

VNU_3 #(quan_width) VNU521 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_521),
	.C2V_2 (C2V_56_521),
	.C2V_3 (C2V_259_521),
	.L (L[7814:7800]),
	.V2C_1 (V2C_521_28),
	.V2C_2 (V2C_521_56),
	.V2C_3 (V2C_521_259),
	.V (V_521)
);

VNU_3 #(quan_width) VNU522 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_522),
	.C2V_2 (C2V_62_522),
	.C2V_3 (C2V_265_522),
	.L (L[7829:7815]),
	.V2C_1 (V2C_522_34),
	.V2C_2 (V2C_522_62),
	.V2C_3 (V2C_522_265),
	.V (V_522)
);

VNU_3 #(quan_width) VNU523 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_523),
	.C2V_2 (C2V_68_523),
	.C2V_3 (C2V_271_523),
	.L (L[7844:7830]),
	.V2C_1 (V2C_523_40),
	.V2C_2 (V2C_523_68),
	.V2C_3 (V2C_523_271),
	.V (V_523)
);

VNU_3 #(quan_width) VNU524 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_524),
	.C2V_2 (C2V_74_524),
	.C2V_3 (C2V_277_524),
	.L (L[7859:7845]),
	.V2C_1 (V2C_524_46),
	.V2C_2 (V2C_524_74),
	.V2C_3 (V2C_524_277),
	.V (V_524)
);

VNU_3 #(quan_width) VNU525 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_525),
	.C2V_2 (C2V_80_525),
	.C2V_3 (C2V_283_525),
	.L (L[7874:7860]),
	.V2C_1 (V2C_525_52),
	.V2C_2 (V2C_525_80),
	.V2C_3 (V2C_525_283),
	.V (V_525)
);

VNU_3 #(quan_width) VNU526 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_526),
	.C2V_2 (C2V_58_526),
	.C2V_3 (C2V_86_526),
	.L (L[7889:7875]),
	.V2C_1 (V2C_526_1),
	.V2C_2 (V2C_526_58),
	.V2C_3 (V2C_526_86),
	.V (V_526)
);

VNU_3 #(quan_width) VNU527 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_527),
	.C2V_2 (C2V_64_527),
	.C2V_3 (C2V_92_527),
	.L (L[7904:7890]),
	.V2C_1 (V2C_527_7),
	.V2C_2 (V2C_527_64),
	.V2C_3 (V2C_527_92),
	.V (V_527)
);

VNU_3 #(quan_width) VNU528 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_528),
	.C2V_2 (C2V_70_528),
	.C2V_3 (C2V_98_528),
	.L (L[7919:7905]),
	.V2C_1 (V2C_528_13),
	.V2C_2 (V2C_528_70),
	.V2C_3 (V2C_528_98),
	.V (V_528)
);

VNU_3 #(quan_width) VNU529 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_529),
	.C2V_2 (C2V_148_529),
	.C2V_3 (C2V_279_529),
	.L (L[7934:7920]),
	.V2C_1 (V2C_529_6),
	.V2C_2 (V2C_529_148),
	.V2C_3 (V2C_529_279),
	.V (V_529)
);

VNU_3 #(quan_width) VNU530 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_530),
	.C2V_2 (C2V_154_530),
	.C2V_3 (C2V_285_530),
	.L (L[7949:7935]),
	.V2C_1 (V2C_530_12),
	.V2C_2 (V2C_530_154),
	.V2C_3 (V2C_530_285),
	.V (V_530)
);

VNU_3 #(quan_width) VNU531 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_531),
	.C2V_2 (C2V_18_531),
	.C2V_3 (C2V_160_531),
	.L (L[7964:7950]),
	.V2C_1 (V2C_531_3),
	.V2C_2 (V2C_531_18),
	.V2C_3 (V2C_531_160),
	.V (V_531)
);

VNU_3 #(quan_width) VNU532 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_532),
	.C2V_2 (C2V_24_532),
	.C2V_3 (C2V_166_532),
	.L (L[7979:7965]),
	.V2C_1 (V2C_532_9),
	.V2C_2 (V2C_532_24),
	.V2C_3 (V2C_532_166),
	.V (V_532)
);

VNU_3 #(quan_width) VNU533 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_533),
	.C2V_2 (C2V_30_533),
	.C2V_3 (C2V_172_533),
	.L (L[7994:7980]),
	.V2C_1 (V2C_533_15),
	.V2C_2 (V2C_533_30),
	.V2C_3 (V2C_533_172),
	.V (V_533)
);

VNU_3 #(quan_width) VNU534 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_534),
	.C2V_2 (C2V_36_534),
	.C2V_3 (C2V_178_534),
	.L (L[8009:7995]),
	.V2C_1 (V2C_534_21),
	.V2C_2 (V2C_534_36),
	.V2C_3 (V2C_534_178),
	.V (V_534)
);

VNU_3 #(quan_width) VNU535 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_535),
	.C2V_2 (C2V_42_535),
	.C2V_3 (C2V_184_535),
	.L (L[8024:8010]),
	.V2C_1 (V2C_535_27),
	.V2C_2 (V2C_535_42),
	.V2C_3 (V2C_535_184),
	.V (V_535)
);

VNU_3 #(quan_width) VNU536 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_536),
	.C2V_2 (C2V_48_536),
	.C2V_3 (C2V_190_536),
	.L (L[8039:8025]),
	.V2C_1 (V2C_536_33),
	.V2C_2 (V2C_536_48),
	.V2C_3 (V2C_536_190),
	.V (V_536)
);

VNU_3 #(quan_width) VNU537 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_537),
	.C2V_2 (C2V_54_537),
	.C2V_3 (C2V_196_537),
	.L (L[8054:8040]),
	.V2C_1 (V2C_537_39),
	.V2C_2 (V2C_537_54),
	.V2C_3 (V2C_537_196),
	.V (V_537)
);

VNU_3 #(quan_width) VNU538 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_538),
	.C2V_2 (C2V_60_538),
	.C2V_3 (C2V_202_538),
	.L (L[8069:8055]),
	.V2C_1 (V2C_538_45),
	.V2C_2 (V2C_538_60),
	.V2C_3 (V2C_538_202),
	.V (V_538)
);

VNU_3 #(quan_width) VNU539 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_539),
	.C2V_2 (C2V_66_539),
	.C2V_3 (C2V_208_539),
	.L (L[8084:8070]),
	.V2C_1 (V2C_539_51),
	.V2C_2 (V2C_539_66),
	.V2C_3 (V2C_539_208),
	.V (V_539)
);

VNU_3 #(quan_width) VNU540 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_540),
	.C2V_2 (C2V_72_540),
	.C2V_3 (C2V_214_540),
	.L (L[8099:8085]),
	.V2C_1 (V2C_540_57),
	.V2C_2 (V2C_540_72),
	.V2C_3 (V2C_540_214),
	.V (V_540)
);

VNU_3 #(quan_width) VNU541 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_541),
	.C2V_2 (C2V_78_541),
	.C2V_3 (C2V_220_541),
	.L (L[8114:8100]),
	.V2C_1 (V2C_541_63),
	.V2C_2 (V2C_541_78),
	.V2C_3 (V2C_541_220),
	.V (V_541)
);

VNU_3 #(quan_width) VNU542 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_542),
	.C2V_2 (C2V_84_542),
	.C2V_3 (C2V_226_542),
	.L (L[8129:8115]),
	.V2C_1 (V2C_542_69),
	.V2C_2 (V2C_542_84),
	.V2C_3 (V2C_542_226),
	.V (V_542)
);

VNU_3 #(quan_width) VNU543 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_543),
	.C2V_2 (C2V_90_543),
	.C2V_3 (C2V_232_543),
	.L (L[8144:8130]),
	.V2C_1 (V2C_543_75),
	.V2C_2 (V2C_543_90),
	.V2C_3 (V2C_543_232),
	.V (V_543)
);

VNU_3 #(quan_width) VNU544 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_544),
	.C2V_2 (C2V_96_544),
	.C2V_3 (C2V_238_544),
	.L (L[8159:8145]),
	.V2C_1 (V2C_544_81),
	.V2C_2 (V2C_544_96),
	.V2C_3 (V2C_544_238),
	.V (V_544)
);

VNU_3 #(quan_width) VNU545 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_545),
	.C2V_2 (C2V_102_545),
	.C2V_3 (C2V_244_545),
	.L (L[8174:8160]),
	.V2C_1 (V2C_545_87),
	.V2C_2 (V2C_545_102),
	.V2C_3 (V2C_545_244),
	.V (V_545)
);

VNU_3 #(quan_width) VNU546 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_93_546),
	.C2V_2 (C2V_108_546),
	.C2V_3 (C2V_250_546),
	.L (L[8189:8175]),
	.V2C_1 (V2C_546_93),
	.V2C_2 (V2C_546_108),
	.V2C_3 (V2C_546_250),
	.V (V_546)
);

VNU_3 #(quan_width) VNU547 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_99_547),
	.C2V_2 (C2V_114_547),
	.C2V_3 (C2V_256_547),
	.L (L[8204:8190]),
	.V2C_1 (V2C_547_99),
	.V2C_2 (V2C_547_114),
	.V2C_3 (V2C_547_256),
	.V (V_547)
);

VNU_3 #(quan_width) VNU548 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_105_548),
	.C2V_2 (C2V_120_548),
	.C2V_3 (C2V_262_548),
	.L (L[8219:8205]),
	.V2C_1 (V2C_548_105),
	.V2C_2 (V2C_548_120),
	.V2C_3 (V2C_548_262),
	.V (V_548)
);

VNU_3 #(quan_width) VNU549 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_111_549),
	.C2V_2 (C2V_126_549),
	.C2V_3 (C2V_268_549),
	.L (L[8234:8220]),
	.V2C_1 (V2C_549_111),
	.V2C_2 (V2C_549_126),
	.V2C_3 (V2C_549_268),
	.V (V_549)
);

VNU_3 #(quan_width) VNU550 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_117_550),
	.C2V_2 (C2V_132_550),
	.C2V_3 (C2V_274_550),
	.L (L[8249:8235]),
	.V2C_1 (V2C_550_117),
	.V2C_2 (V2C_550_132),
	.V2C_3 (V2C_550_274),
	.V (V_550)
);

VNU_3 #(quan_width) VNU551 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_123_551),
	.C2V_2 (C2V_138_551),
	.C2V_3 (C2V_280_551),
	.L (L[8264:8250]),
	.V2C_1 (V2C_551_123),
	.V2C_2 (V2C_551_138),
	.V2C_3 (V2C_551_280),
	.V (V_551)
);

VNU_3 #(quan_width) VNU552 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_129_552),
	.C2V_2 (C2V_144_552),
	.C2V_3 (C2V_286_552),
	.L (L[8279:8265]),
	.V2C_1 (V2C_552_129),
	.V2C_2 (V2C_552_144),
	.V2C_3 (V2C_552_286),
	.V (V_552)
);

VNU_3 #(quan_width) VNU553 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_553),
	.C2V_2 (C2V_135_553),
	.C2V_3 (C2V_150_553),
	.L (L[8294:8280]),
	.V2C_1 (V2C_553_4),
	.V2C_2 (V2C_553_135),
	.V2C_3 (V2C_553_150),
	.V (V_553)
);

VNU_3 #(quan_width) VNU554 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_554),
	.C2V_2 (C2V_141_554),
	.C2V_3 (C2V_156_554),
	.L (L[8309:8295]),
	.V2C_1 (V2C_554_10),
	.V2C_2 (V2C_554_141),
	.V2C_3 (V2C_554_156),
	.V (V_554)
);

VNU_3 #(quan_width) VNU555 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_555),
	.C2V_2 (C2V_147_555),
	.C2V_3 (C2V_162_555),
	.L (L[8324:8310]),
	.V2C_1 (V2C_555_16),
	.V2C_2 (V2C_555_147),
	.V2C_3 (V2C_555_162),
	.V (V_555)
);

VNU_3 #(quan_width) VNU556 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_556),
	.C2V_2 (C2V_153_556),
	.C2V_3 (C2V_168_556),
	.L (L[8339:8325]),
	.V2C_1 (V2C_556_22),
	.V2C_2 (V2C_556_153),
	.V2C_3 (V2C_556_168),
	.V (V_556)
);

VNU_3 #(quan_width) VNU557 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_557),
	.C2V_2 (C2V_159_557),
	.C2V_3 (C2V_174_557),
	.L (L[8354:8340]),
	.V2C_1 (V2C_557_28),
	.V2C_2 (V2C_557_159),
	.V2C_3 (V2C_557_174),
	.V (V_557)
);

VNU_3 #(quan_width) VNU558 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_558),
	.C2V_2 (C2V_165_558),
	.C2V_3 (C2V_180_558),
	.L (L[8369:8355]),
	.V2C_1 (V2C_558_34),
	.V2C_2 (V2C_558_165),
	.V2C_3 (V2C_558_180),
	.V (V_558)
);

VNU_3 #(quan_width) VNU559 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_559),
	.C2V_2 (C2V_171_559),
	.C2V_3 (C2V_186_559),
	.L (L[8384:8370]),
	.V2C_1 (V2C_559_40),
	.V2C_2 (V2C_559_171),
	.V2C_3 (V2C_559_186),
	.V (V_559)
);

VNU_3 #(quan_width) VNU560 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_560),
	.C2V_2 (C2V_177_560),
	.C2V_3 (C2V_192_560),
	.L (L[8399:8385]),
	.V2C_1 (V2C_560_46),
	.V2C_2 (V2C_560_177),
	.V2C_3 (V2C_560_192),
	.V (V_560)
);

VNU_3 #(quan_width) VNU561 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_561),
	.C2V_2 (C2V_183_561),
	.C2V_3 (C2V_198_561),
	.L (L[8414:8400]),
	.V2C_1 (V2C_561_52),
	.V2C_2 (V2C_561_183),
	.V2C_3 (V2C_561_198),
	.V (V_561)
);

VNU_3 #(quan_width) VNU562 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_562),
	.C2V_2 (C2V_189_562),
	.C2V_3 (C2V_204_562),
	.L (L[8429:8415]),
	.V2C_1 (V2C_562_58),
	.V2C_2 (V2C_562_189),
	.V2C_3 (V2C_562_204),
	.V (V_562)
);

VNU_3 #(quan_width) VNU563 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_563),
	.C2V_2 (C2V_195_563),
	.C2V_3 (C2V_210_563),
	.L (L[8444:8430]),
	.V2C_1 (V2C_563_64),
	.V2C_2 (V2C_563_195),
	.V2C_3 (V2C_563_210),
	.V (V_563)
);

VNU_3 #(quan_width) VNU564 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_564),
	.C2V_2 (C2V_201_564),
	.C2V_3 (C2V_216_564),
	.L (L[8459:8445]),
	.V2C_1 (V2C_564_70),
	.V2C_2 (V2C_564_201),
	.V2C_3 (V2C_564_216),
	.V (V_564)
);

VNU_3 #(quan_width) VNU565 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_565),
	.C2V_2 (C2V_207_565),
	.C2V_3 (C2V_222_565),
	.L (L[8474:8460]),
	.V2C_1 (V2C_565_76),
	.V2C_2 (V2C_565_207),
	.V2C_3 (V2C_565_222),
	.V (V_565)
);

VNU_3 #(quan_width) VNU566 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_566),
	.C2V_2 (C2V_213_566),
	.C2V_3 (C2V_228_566),
	.L (L[8489:8475]),
	.V2C_1 (V2C_566_82),
	.V2C_2 (V2C_566_213),
	.V2C_3 (V2C_566_228),
	.V (V_566)
);

VNU_3 #(quan_width) VNU567 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_567),
	.C2V_2 (C2V_219_567),
	.C2V_3 (C2V_234_567),
	.L (L[8504:8490]),
	.V2C_1 (V2C_567_88),
	.V2C_2 (V2C_567_219),
	.V2C_3 (V2C_567_234),
	.V (V_567)
);

VNU_3 #(quan_width) VNU568 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_568),
	.C2V_2 (C2V_225_568),
	.C2V_3 (C2V_240_568),
	.L (L[8519:8505]),
	.V2C_1 (V2C_568_94),
	.V2C_2 (V2C_568_225),
	.V2C_3 (V2C_568_240),
	.V (V_568)
);

VNU_3 #(quan_width) VNU569 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_569),
	.C2V_2 (C2V_231_569),
	.C2V_3 (C2V_246_569),
	.L (L[8534:8520]),
	.V2C_1 (V2C_569_100),
	.V2C_2 (V2C_569_231),
	.V2C_3 (V2C_569_246),
	.V (V_569)
);

VNU_3 #(quan_width) VNU570 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_570),
	.C2V_2 (C2V_237_570),
	.C2V_3 (C2V_252_570),
	.L (L[8549:8535]),
	.V2C_1 (V2C_570_106),
	.V2C_2 (V2C_570_237),
	.V2C_3 (V2C_570_252),
	.V (V_570)
);

VNU_3 #(quan_width) VNU571 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_571),
	.C2V_2 (C2V_243_571),
	.C2V_3 (C2V_258_571),
	.L (L[8564:8550]),
	.V2C_1 (V2C_571_112),
	.V2C_2 (V2C_571_243),
	.V2C_3 (V2C_571_258),
	.V (V_571)
);

VNU_3 #(quan_width) VNU572 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_118_572),
	.C2V_2 (C2V_249_572),
	.C2V_3 (C2V_264_572),
	.L (L[8579:8565]),
	.V2C_1 (V2C_572_118),
	.V2C_2 (V2C_572_249),
	.V2C_3 (V2C_572_264),
	.V (V_572)
);

VNU_3 #(quan_width) VNU573 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_124_573),
	.C2V_2 (C2V_255_573),
	.C2V_3 (C2V_270_573),
	.L (L[8594:8580]),
	.V2C_1 (V2C_573_124),
	.V2C_2 (V2C_573_255),
	.V2C_3 (V2C_573_270),
	.V (V_573)
);

VNU_3 #(quan_width) VNU574 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_130_574),
	.C2V_2 (C2V_261_574),
	.C2V_3 (C2V_276_574),
	.L (L[8609:8595]),
	.V2C_1 (V2C_574_130),
	.V2C_2 (V2C_574_261),
	.V2C_3 (V2C_574_276),
	.V (V_574)
);

VNU_3 #(quan_width) VNU575 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_136_575),
	.C2V_2 (C2V_267_575),
	.C2V_3 (C2V_282_575),
	.L (L[8624:8610]),
	.V2C_1 (V2C_575_136),
	.V2C_2 (V2C_575_267),
	.V2C_3 (V2C_575_282),
	.V (V_575)
);

VNU_3 #(quan_width) VNU576 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_142_576),
	.C2V_2 (C2V_273_576),
	.C2V_3 (C2V_288_576),
	.L (L[8639:8625]),
	.V2C_1 (V2C_576_142),
	.V2C_2 (V2C_576_273),
	.V2C_3 (V2C_576_288),
	.V (V_576)
);

VNU_3 #(quan_width) VNU577 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_577),
	.C2V_2 (C2V_96_577),
	.C2V_3 (C2V_225_577),
	.L (L[8654:8640]),
	.V2C_1 (V2C_577_64),
	.V2C_2 (V2C_577_96),
	.V2C_3 (V2C_577_225),
	.V (V_577)
);

VNU_3 #(quan_width) VNU578 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_578),
	.C2V_2 (C2V_102_578),
	.C2V_3 (C2V_231_578),
	.L (L[8669:8655]),
	.V2C_1 (V2C_578_70),
	.V2C_2 (V2C_578_102),
	.V2C_3 (V2C_578_231),
	.V (V_578)
);

VNU_3 #(quan_width) VNU579 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_579),
	.C2V_2 (C2V_108_579),
	.C2V_3 (C2V_237_579),
	.L (L[8684:8670]),
	.V2C_1 (V2C_579_76),
	.V2C_2 (V2C_579_108),
	.V2C_3 (V2C_579_237),
	.V (V_579)
);

VNU_3 #(quan_width) VNU580 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_580),
	.C2V_2 (C2V_114_580),
	.C2V_3 (C2V_243_580),
	.L (L[8699:8685]),
	.V2C_1 (V2C_580_82),
	.V2C_2 (V2C_580_114),
	.V2C_3 (V2C_580_243),
	.V (V_580)
);

VNU_3 #(quan_width) VNU581 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_581),
	.C2V_2 (C2V_120_581),
	.C2V_3 (C2V_249_581),
	.L (L[8714:8700]),
	.V2C_1 (V2C_581_88),
	.V2C_2 (V2C_581_120),
	.V2C_3 (V2C_581_249),
	.V (V_581)
);

VNU_3 #(quan_width) VNU582 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_582),
	.C2V_2 (C2V_126_582),
	.C2V_3 (C2V_255_582),
	.L (L[8729:8715]),
	.V2C_1 (V2C_582_94),
	.V2C_2 (V2C_582_126),
	.V2C_3 (V2C_582_255),
	.V (V_582)
);

VNU_3 #(quan_width) VNU583 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_583),
	.C2V_2 (C2V_132_583),
	.C2V_3 (C2V_261_583),
	.L (L[8744:8730]),
	.V2C_1 (V2C_583_100),
	.V2C_2 (V2C_583_132),
	.V2C_3 (V2C_583_261),
	.V (V_583)
);

VNU_3 #(quan_width) VNU584 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_584),
	.C2V_2 (C2V_138_584),
	.C2V_3 (C2V_267_584),
	.L (L[8759:8745]),
	.V2C_1 (V2C_584_106),
	.V2C_2 (V2C_584_138),
	.V2C_3 (V2C_584_267),
	.V (V_584)
);

VNU_3 #(quan_width) VNU585 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_585),
	.C2V_2 (C2V_144_585),
	.C2V_3 (C2V_273_585),
	.L (L[8774:8760]),
	.V2C_1 (V2C_585_112),
	.V2C_2 (V2C_585_144),
	.V2C_3 (V2C_585_273),
	.V (V_585)
);

VNU_3 #(quan_width) VNU586 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_118_586),
	.C2V_2 (C2V_150_586),
	.C2V_3 (C2V_279_586),
	.L (L[8789:8775]),
	.V2C_1 (V2C_586_118),
	.V2C_2 (V2C_586_150),
	.V2C_3 (V2C_586_279),
	.V (V_586)
);

VNU_3 #(quan_width) VNU587 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_124_587),
	.C2V_2 (C2V_156_587),
	.C2V_3 (C2V_285_587),
	.L (L[8804:8790]),
	.V2C_1 (V2C_587_124),
	.V2C_2 (V2C_587_156),
	.V2C_3 (V2C_587_285),
	.V (V_587)
);

VNU_3 #(quan_width) VNU588 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_588),
	.C2V_2 (C2V_130_588),
	.C2V_3 (C2V_162_588),
	.L (L[8819:8805]),
	.V2C_1 (V2C_588_3),
	.V2C_2 (V2C_588_130),
	.V2C_3 (V2C_588_162),
	.V (V_588)
);

VNU_3 #(quan_width) VNU589 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_589),
	.C2V_2 (C2V_136_589),
	.C2V_3 (C2V_168_589),
	.L (L[8834:8820]),
	.V2C_1 (V2C_589_9),
	.V2C_2 (V2C_589_136),
	.V2C_3 (V2C_589_168),
	.V (V_589)
);

VNU_3 #(quan_width) VNU590 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_590),
	.C2V_2 (C2V_142_590),
	.C2V_3 (C2V_174_590),
	.L (L[8849:8835]),
	.V2C_1 (V2C_590_15),
	.V2C_2 (V2C_590_142),
	.V2C_3 (V2C_590_174),
	.V (V_590)
);

VNU_3 #(quan_width) VNU591 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_591),
	.C2V_2 (C2V_148_591),
	.C2V_3 (C2V_180_591),
	.L (L[8864:8850]),
	.V2C_1 (V2C_591_21),
	.V2C_2 (V2C_591_148),
	.V2C_3 (V2C_591_180),
	.V (V_591)
);

VNU_3 #(quan_width) VNU592 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_592),
	.C2V_2 (C2V_154_592),
	.C2V_3 (C2V_186_592),
	.L (L[8879:8865]),
	.V2C_1 (V2C_592_27),
	.V2C_2 (V2C_592_154),
	.V2C_3 (V2C_592_186),
	.V (V_592)
);

VNU_3 #(quan_width) VNU593 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_593),
	.C2V_2 (C2V_160_593),
	.C2V_3 (C2V_192_593),
	.L (L[8894:8880]),
	.V2C_1 (V2C_593_33),
	.V2C_2 (V2C_593_160),
	.V2C_3 (V2C_593_192),
	.V (V_593)
);

VNU_3 #(quan_width) VNU594 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_594),
	.C2V_2 (C2V_166_594),
	.C2V_3 (C2V_198_594),
	.L (L[8909:8895]),
	.V2C_1 (V2C_594_39),
	.V2C_2 (V2C_594_166),
	.V2C_3 (V2C_594_198),
	.V (V_594)
);

VNU_3 #(quan_width) VNU595 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_595),
	.C2V_2 (C2V_172_595),
	.C2V_3 (C2V_204_595),
	.L (L[8924:8910]),
	.V2C_1 (V2C_595_45),
	.V2C_2 (V2C_595_172),
	.V2C_3 (V2C_595_204),
	.V (V_595)
);

VNU_3 #(quan_width) VNU596 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_596),
	.C2V_2 (C2V_178_596),
	.C2V_3 (C2V_210_596),
	.L (L[8939:8925]),
	.V2C_1 (V2C_596_51),
	.V2C_2 (V2C_596_178),
	.V2C_3 (V2C_596_210),
	.V (V_596)
);

VNU_3 #(quan_width) VNU597 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_597),
	.C2V_2 (C2V_184_597),
	.C2V_3 (C2V_216_597),
	.L (L[8954:8940]),
	.V2C_1 (V2C_597_57),
	.V2C_2 (V2C_597_184),
	.V2C_3 (V2C_597_216),
	.V (V_597)
);

VNU_3 #(quan_width) VNU598 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_598),
	.C2V_2 (C2V_190_598),
	.C2V_3 (C2V_222_598),
	.L (L[8969:8955]),
	.V2C_1 (V2C_598_63),
	.V2C_2 (V2C_598_190),
	.V2C_3 (V2C_598_222),
	.V (V_598)
);

VNU_3 #(quan_width) VNU599 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_599),
	.C2V_2 (C2V_196_599),
	.C2V_3 (C2V_228_599),
	.L (L[8984:8970]),
	.V2C_1 (V2C_599_69),
	.V2C_2 (V2C_599_196),
	.V2C_3 (V2C_599_228),
	.V (V_599)
);

VNU_3 #(quan_width) VNU600 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_600),
	.C2V_2 (C2V_202_600),
	.C2V_3 (C2V_234_600),
	.L (L[8999:8985]),
	.V2C_1 (V2C_600_75),
	.V2C_2 (V2C_600_202),
	.V2C_3 (V2C_600_234),
	.V (V_600)
);

VNU_3 #(quan_width) VNU601 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_601),
	.C2V_2 (C2V_208_601),
	.C2V_3 (C2V_240_601),
	.L (L[9014:9000]),
	.V2C_1 (V2C_601_81),
	.V2C_2 (V2C_601_208),
	.V2C_3 (V2C_601_240),
	.V (V_601)
);

VNU_3 #(quan_width) VNU602 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_602),
	.C2V_2 (C2V_214_602),
	.C2V_3 (C2V_246_602),
	.L (L[9029:9015]),
	.V2C_1 (V2C_602_87),
	.V2C_2 (V2C_602_214),
	.V2C_3 (V2C_602_246),
	.V (V_602)
);

VNU_3 #(quan_width) VNU603 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_93_603),
	.C2V_2 (C2V_220_603),
	.C2V_3 (C2V_252_603),
	.L (L[9044:9030]),
	.V2C_1 (V2C_603_93),
	.V2C_2 (V2C_603_220),
	.V2C_3 (V2C_603_252),
	.V (V_603)
);

VNU_3 #(quan_width) VNU604 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_99_604),
	.C2V_2 (C2V_226_604),
	.C2V_3 (C2V_258_604),
	.L (L[9059:9045]),
	.V2C_1 (V2C_604_99),
	.V2C_2 (V2C_604_226),
	.V2C_3 (V2C_604_258),
	.V (V_604)
);

VNU_3 #(quan_width) VNU605 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_105_605),
	.C2V_2 (C2V_232_605),
	.C2V_3 (C2V_264_605),
	.L (L[9074:9060]),
	.V2C_1 (V2C_605_105),
	.V2C_2 (V2C_605_232),
	.V2C_3 (V2C_605_264),
	.V (V_605)
);

VNU_3 #(quan_width) VNU606 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_111_606),
	.C2V_2 (C2V_238_606),
	.C2V_3 (C2V_270_606),
	.L (L[9089:9075]),
	.V2C_1 (V2C_606_111),
	.V2C_2 (V2C_606_238),
	.V2C_3 (V2C_606_270),
	.V (V_606)
);

VNU_3 #(quan_width) VNU607 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_117_607),
	.C2V_2 (C2V_244_607),
	.C2V_3 (C2V_276_607),
	.L (L[9104:9090]),
	.V2C_1 (V2C_607_117),
	.V2C_2 (V2C_607_244),
	.V2C_3 (V2C_607_276),
	.V (V_607)
);

VNU_3 #(quan_width) VNU608 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_123_608),
	.C2V_2 (C2V_250_608),
	.C2V_3 (C2V_282_608),
	.L (L[9119:9105]),
	.V2C_1 (V2C_608_123),
	.V2C_2 (V2C_608_250),
	.V2C_3 (V2C_608_282),
	.V (V_608)
);

VNU_3 #(quan_width) VNU609 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_129_609),
	.C2V_2 (C2V_256_609),
	.C2V_3 (C2V_288_609),
	.L (L[9134:9120]),
	.V2C_1 (V2C_609_129),
	.V2C_2 (V2C_609_256),
	.V2C_3 (V2C_609_288),
	.V (V_609)
);

VNU_3 #(quan_width) VNU610 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_610),
	.C2V_2 (C2V_135_610),
	.C2V_3 (C2V_262_610),
	.L (L[9149:9135]),
	.V2C_1 (V2C_610_6),
	.V2C_2 (V2C_610_135),
	.V2C_3 (V2C_610_262),
	.V (V_610)
);

VNU_3 #(quan_width) VNU611 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_611),
	.C2V_2 (C2V_141_611),
	.C2V_3 (C2V_268_611),
	.L (L[9164:9150]),
	.V2C_1 (V2C_611_12),
	.V2C_2 (V2C_611_141),
	.V2C_3 (V2C_611_268),
	.V (V_611)
);

VNU_3 #(quan_width) VNU612 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_612),
	.C2V_2 (C2V_147_612),
	.C2V_3 (C2V_274_612),
	.L (L[9179:9165]),
	.V2C_1 (V2C_612_18),
	.V2C_2 (V2C_612_147),
	.V2C_3 (V2C_612_274),
	.V (V_612)
);

VNU_3 #(quan_width) VNU613 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_613),
	.C2V_2 (C2V_153_613),
	.C2V_3 (C2V_280_613),
	.L (L[9194:9180]),
	.V2C_1 (V2C_613_24),
	.V2C_2 (V2C_613_153),
	.V2C_3 (V2C_613_280),
	.V (V_613)
);

VNU_3 #(quan_width) VNU614 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_614),
	.C2V_2 (C2V_159_614),
	.C2V_3 (C2V_286_614),
	.L (L[9209:9195]),
	.V2C_1 (V2C_614_30),
	.V2C_2 (V2C_614_159),
	.V2C_3 (V2C_614_286),
	.V (V_614)
);

VNU_3 #(quan_width) VNU615 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_615),
	.C2V_2 (C2V_36_615),
	.C2V_3 (C2V_165_615),
	.L (L[9224:9210]),
	.V2C_1 (V2C_615_4),
	.V2C_2 (V2C_615_36),
	.V2C_3 (V2C_615_165),
	.V (V_615)
);

VNU_3 #(quan_width) VNU616 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_616),
	.C2V_2 (C2V_42_616),
	.C2V_3 (C2V_171_616),
	.L (L[9239:9225]),
	.V2C_1 (V2C_616_10),
	.V2C_2 (V2C_616_42),
	.V2C_3 (V2C_616_171),
	.V (V_616)
);

VNU_3 #(quan_width) VNU617 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_617),
	.C2V_2 (C2V_48_617),
	.C2V_3 (C2V_177_617),
	.L (L[9254:9240]),
	.V2C_1 (V2C_617_16),
	.V2C_2 (V2C_617_48),
	.V2C_3 (V2C_617_177),
	.V (V_617)
);

VNU_3 #(quan_width) VNU618 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_618),
	.C2V_2 (C2V_54_618),
	.C2V_3 (C2V_183_618),
	.L (L[9269:9255]),
	.V2C_1 (V2C_618_22),
	.V2C_2 (V2C_618_54),
	.V2C_3 (V2C_618_183),
	.V (V_618)
);

VNU_3 #(quan_width) VNU619 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_619),
	.C2V_2 (C2V_60_619),
	.C2V_3 (C2V_189_619),
	.L (L[9284:9270]),
	.V2C_1 (V2C_619_28),
	.V2C_2 (V2C_619_60),
	.V2C_3 (V2C_619_189),
	.V (V_619)
);

VNU_3 #(quan_width) VNU620 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_620),
	.C2V_2 (C2V_66_620),
	.C2V_3 (C2V_195_620),
	.L (L[9299:9285]),
	.V2C_1 (V2C_620_34),
	.V2C_2 (V2C_620_66),
	.V2C_3 (V2C_620_195),
	.V (V_620)
);

VNU_3 #(quan_width) VNU621 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_621),
	.C2V_2 (C2V_72_621),
	.C2V_3 (C2V_201_621),
	.L (L[9314:9300]),
	.V2C_1 (V2C_621_40),
	.V2C_2 (V2C_621_72),
	.V2C_3 (V2C_621_201),
	.V (V_621)
);

VNU_3 #(quan_width) VNU622 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_622),
	.C2V_2 (C2V_78_622),
	.C2V_3 (C2V_207_622),
	.L (L[9329:9315]),
	.V2C_1 (V2C_622_46),
	.V2C_2 (V2C_622_78),
	.V2C_3 (V2C_622_207),
	.V (V_622)
);

VNU_3 #(quan_width) VNU623 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_623),
	.C2V_2 (C2V_84_623),
	.C2V_3 (C2V_213_623),
	.L (L[9344:9330]),
	.V2C_1 (V2C_623_52),
	.V2C_2 (V2C_623_84),
	.V2C_3 (V2C_623_213),
	.V (V_623)
);

VNU_3 #(quan_width) VNU624 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_624),
	.C2V_2 (C2V_90_624),
	.C2V_3 (C2V_219_624),
	.L (L[9359:9345]),
	.V2C_1 (V2C_624_58),
	.V2C_2 (V2C_624_90),
	.V2C_3 (V2C_624_219),
	.V (V_624)
);

VNU_3 #(quan_width) VNU625 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_625),
	.C2V_2 (C2V_57_625),
	.C2V_3 (C2V_202_625),
	.L (L[9374:9360]),
	.V2C_1 (V2C_625_8),
	.V2C_2 (V2C_625_57),
	.V2C_3 (V2C_625_202),
	.V (V_625)
);

VNU_3 #(quan_width) VNU626 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_626),
	.C2V_2 (C2V_63_626),
	.C2V_3 (C2V_208_626),
	.L (L[9389:9375]),
	.V2C_1 (V2C_626_14),
	.V2C_2 (V2C_626_63),
	.V2C_3 (V2C_626_208),
	.V (V_626)
);

VNU_3 #(quan_width) VNU627 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_627),
	.C2V_2 (C2V_69_627),
	.C2V_3 (C2V_214_627),
	.L (L[9404:9390]),
	.V2C_1 (V2C_627_20),
	.V2C_2 (V2C_627_69),
	.V2C_3 (V2C_627_214),
	.V (V_627)
);

VNU_3 #(quan_width) VNU628 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_628),
	.C2V_2 (C2V_75_628),
	.C2V_3 (C2V_220_628),
	.L (L[9419:9405]),
	.V2C_1 (V2C_628_26),
	.V2C_2 (V2C_628_75),
	.V2C_3 (V2C_628_220),
	.V (V_628)
);

VNU_3 #(quan_width) VNU629 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_629),
	.C2V_2 (C2V_81_629),
	.C2V_3 (C2V_226_629),
	.L (L[9434:9420]),
	.V2C_1 (V2C_629_32),
	.V2C_2 (V2C_629_81),
	.V2C_3 (V2C_629_226),
	.V (V_629)
);

VNU_3 #(quan_width) VNU630 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_630),
	.C2V_2 (C2V_87_630),
	.C2V_3 (C2V_232_630),
	.L (L[9449:9435]),
	.V2C_1 (V2C_630_38),
	.V2C_2 (V2C_630_87),
	.V2C_3 (V2C_630_232),
	.V (V_630)
);

VNU_3 #(quan_width) VNU631 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_631),
	.C2V_2 (C2V_93_631),
	.C2V_3 (C2V_238_631),
	.L (L[9464:9450]),
	.V2C_1 (V2C_631_44),
	.V2C_2 (V2C_631_93),
	.V2C_3 (V2C_631_238),
	.V (V_631)
);

VNU_3 #(quan_width) VNU632 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_632),
	.C2V_2 (C2V_99_632),
	.C2V_3 (C2V_244_632),
	.L (L[9479:9465]),
	.V2C_1 (V2C_632_50),
	.V2C_2 (V2C_632_99),
	.V2C_3 (V2C_632_244),
	.V (V_632)
);

VNU_3 #(quan_width) VNU633 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_633),
	.C2V_2 (C2V_105_633),
	.C2V_3 (C2V_250_633),
	.L (L[9494:9480]),
	.V2C_1 (V2C_633_56),
	.V2C_2 (V2C_633_105),
	.V2C_3 (V2C_633_250),
	.V (V_633)
);

VNU_3 #(quan_width) VNU634 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_634),
	.C2V_2 (C2V_111_634),
	.C2V_3 (C2V_256_634),
	.L (L[9509:9495]),
	.V2C_1 (V2C_634_62),
	.V2C_2 (V2C_634_111),
	.V2C_3 (V2C_634_256),
	.V (V_634)
);

VNU_3 #(quan_width) VNU635 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_635),
	.C2V_2 (C2V_117_635),
	.C2V_3 (C2V_262_635),
	.L (L[9524:9510]),
	.V2C_1 (V2C_635_68),
	.V2C_2 (V2C_635_117),
	.V2C_3 (V2C_635_262),
	.V (V_635)
);

VNU_3 #(quan_width) VNU636 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_636),
	.C2V_2 (C2V_123_636),
	.C2V_3 (C2V_268_636),
	.L (L[9539:9525]),
	.V2C_1 (V2C_636_74),
	.V2C_2 (V2C_636_123),
	.V2C_3 (V2C_636_268),
	.V (V_636)
);

VNU_3 #(quan_width) VNU637 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_80_637),
	.C2V_2 (C2V_129_637),
	.C2V_3 (C2V_274_637),
	.L (L[9554:9540]),
	.V2C_1 (V2C_637_80),
	.V2C_2 (V2C_637_129),
	.V2C_3 (V2C_637_274),
	.V (V_637)
);

VNU_3 #(quan_width) VNU638 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_86_638),
	.C2V_2 (C2V_135_638),
	.C2V_3 (C2V_280_638),
	.L (L[9569:9555]),
	.V2C_1 (V2C_638_86),
	.V2C_2 (V2C_638_135),
	.V2C_3 (V2C_638_280),
	.V (V_638)
);

VNU_3 #(quan_width) VNU639 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_92_639),
	.C2V_2 (C2V_141_639),
	.C2V_3 (C2V_286_639),
	.L (L[9584:9570]),
	.V2C_1 (V2C_639_92),
	.V2C_2 (V2C_639_141),
	.V2C_3 (V2C_639_286),
	.V (V_639)
);

VNU_3 #(quan_width) VNU640 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_640),
	.C2V_2 (C2V_98_640),
	.C2V_3 (C2V_147_640),
	.L (L[9599:9585]),
	.V2C_1 (V2C_640_4),
	.V2C_2 (V2C_640_98),
	.V2C_3 (V2C_640_147),
	.V (V_640)
);

VNU_3 #(quan_width) VNU641 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_641),
	.C2V_2 (C2V_104_641),
	.C2V_3 (C2V_153_641),
	.L (L[9614:9600]),
	.V2C_1 (V2C_641_10),
	.V2C_2 (V2C_641_104),
	.V2C_3 (V2C_641_153),
	.V (V_641)
);

VNU_3 #(quan_width) VNU642 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_642),
	.C2V_2 (C2V_110_642),
	.C2V_3 (C2V_159_642),
	.L (L[9629:9615]),
	.V2C_1 (V2C_642_16),
	.V2C_2 (V2C_642_110),
	.V2C_3 (V2C_642_159),
	.V (V_642)
);

VNU_3 #(quan_width) VNU643 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_643),
	.C2V_2 (C2V_116_643),
	.C2V_3 (C2V_165_643),
	.L (L[9644:9630]),
	.V2C_1 (V2C_643_22),
	.V2C_2 (V2C_643_116),
	.V2C_3 (V2C_643_165),
	.V (V_643)
);

VNU_3 #(quan_width) VNU644 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_644),
	.C2V_2 (C2V_122_644),
	.C2V_3 (C2V_171_644),
	.L (L[9659:9645]),
	.V2C_1 (V2C_644_28),
	.V2C_2 (V2C_644_122),
	.V2C_3 (V2C_644_171),
	.V (V_644)
);

VNU_3 #(quan_width) VNU645 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_645),
	.C2V_2 (C2V_128_645),
	.C2V_3 (C2V_177_645),
	.L (L[9674:9660]),
	.V2C_1 (V2C_645_34),
	.V2C_2 (V2C_645_128),
	.V2C_3 (V2C_645_177),
	.V (V_645)
);

VNU_3 #(quan_width) VNU646 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_646),
	.C2V_2 (C2V_134_646),
	.C2V_3 (C2V_183_646),
	.L (L[9689:9675]),
	.V2C_1 (V2C_646_40),
	.V2C_2 (V2C_646_134),
	.V2C_3 (V2C_646_183),
	.V (V_646)
);

VNU_3 #(quan_width) VNU647 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_647),
	.C2V_2 (C2V_140_647),
	.C2V_3 (C2V_189_647),
	.L (L[9704:9690]),
	.V2C_1 (V2C_647_46),
	.V2C_2 (V2C_647_140),
	.V2C_3 (V2C_647_189),
	.V (V_647)
);

VNU_3 #(quan_width) VNU648 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_648),
	.C2V_2 (C2V_146_648),
	.C2V_3 (C2V_195_648),
	.L (L[9719:9705]),
	.V2C_1 (V2C_648_52),
	.V2C_2 (V2C_648_146),
	.V2C_3 (V2C_648_195),
	.V (V_648)
);

VNU_3 #(quan_width) VNU649 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_649),
	.C2V_2 (C2V_152_649),
	.C2V_3 (C2V_201_649),
	.L (L[9734:9720]),
	.V2C_1 (V2C_649_58),
	.V2C_2 (V2C_649_152),
	.V2C_3 (V2C_649_201),
	.V (V_649)
);

VNU_3 #(quan_width) VNU650 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_650),
	.C2V_2 (C2V_158_650),
	.C2V_3 (C2V_207_650),
	.L (L[9749:9735]),
	.V2C_1 (V2C_650_64),
	.V2C_2 (V2C_650_158),
	.V2C_3 (V2C_650_207),
	.V (V_650)
);

VNU_3 #(quan_width) VNU651 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_651),
	.C2V_2 (C2V_164_651),
	.C2V_3 (C2V_213_651),
	.L (L[9764:9750]),
	.V2C_1 (V2C_651_70),
	.V2C_2 (V2C_651_164),
	.V2C_3 (V2C_651_213),
	.V (V_651)
);

VNU_3 #(quan_width) VNU652 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_652),
	.C2V_2 (C2V_170_652),
	.C2V_3 (C2V_219_652),
	.L (L[9779:9765]),
	.V2C_1 (V2C_652_76),
	.V2C_2 (V2C_652_170),
	.V2C_3 (V2C_652_219),
	.V (V_652)
);

VNU_3 #(quan_width) VNU653 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_653),
	.C2V_2 (C2V_176_653),
	.C2V_3 (C2V_225_653),
	.L (L[9794:9780]),
	.V2C_1 (V2C_653_82),
	.V2C_2 (V2C_653_176),
	.V2C_3 (V2C_653_225),
	.V (V_653)
);

VNU_3 #(quan_width) VNU654 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_654),
	.C2V_2 (C2V_182_654),
	.C2V_3 (C2V_231_654),
	.L (L[9809:9795]),
	.V2C_1 (V2C_654_88),
	.V2C_2 (V2C_654_182),
	.V2C_3 (V2C_654_231),
	.V (V_654)
);

VNU_3 #(quan_width) VNU655 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_655),
	.C2V_2 (C2V_188_655),
	.C2V_3 (C2V_237_655),
	.L (L[9824:9810]),
	.V2C_1 (V2C_655_94),
	.V2C_2 (V2C_655_188),
	.V2C_3 (V2C_655_237),
	.V (V_655)
);

VNU_3 #(quan_width) VNU656 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_656),
	.C2V_2 (C2V_194_656),
	.C2V_3 (C2V_243_656),
	.L (L[9839:9825]),
	.V2C_1 (V2C_656_100),
	.V2C_2 (V2C_656_194),
	.V2C_3 (V2C_656_243),
	.V (V_656)
);

VNU_3 #(quan_width) VNU657 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_657),
	.C2V_2 (C2V_200_657),
	.C2V_3 (C2V_249_657),
	.L (L[9854:9840]),
	.V2C_1 (V2C_657_106),
	.V2C_2 (V2C_657_200),
	.V2C_3 (V2C_657_249),
	.V (V_657)
);

VNU_3 #(quan_width) VNU658 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_658),
	.C2V_2 (C2V_206_658),
	.C2V_3 (C2V_255_658),
	.L (L[9869:9855]),
	.V2C_1 (V2C_658_112),
	.V2C_2 (V2C_658_206),
	.V2C_3 (V2C_658_255),
	.V (V_658)
);

VNU_3 #(quan_width) VNU659 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_118_659),
	.C2V_2 (C2V_212_659),
	.C2V_3 (C2V_261_659),
	.L (L[9884:9870]),
	.V2C_1 (V2C_659_118),
	.V2C_2 (V2C_659_212),
	.V2C_3 (V2C_659_261),
	.V (V_659)
);

VNU_3 #(quan_width) VNU660 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_124_660),
	.C2V_2 (C2V_218_660),
	.C2V_3 (C2V_267_660),
	.L (L[9899:9885]),
	.V2C_1 (V2C_660_124),
	.V2C_2 (V2C_660_218),
	.V2C_3 (V2C_660_267),
	.V (V_660)
);

VNU_3 #(quan_width) VNU661 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_130_661),
	.C2V_2 (C2V_224_661),
	.C2V_3 (C2V_273_661),
	.L (L[9914:9900]),
	.V2C_1 (V2C_661_130),
	.V2C_2 (V2C_661_224),
	.V2C_3 (V2C_661_273),
	.V (V_661)
);

VNU_3 #(quan_width) VNU662 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_136_662),
	.C2V_2 (C2V_230_662),
	.C2V_3 (C2V_279_662),
	.L (L[9929:9915]),
	.V2C_1 (V2C_662_136),
	.V2C_2 (V2C_662_230),
	.V2C_3 (V2C_662_279),
	.V (V_662)
);

VNU_3 #(quan_width) VNU663 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_142_663),
	.C2V_2 (C2V_236_663),
	.C2V_3 (C2V_285_663),
	.L (L[9944:9930]),
	.V2C_1 (V2C_663_142),
	.V2C_2 (V2C_663_236),
	.V2C_3 (V2C_663_285),
	.V (V_663)
);

VNU_3 #(quan_width) VNU664 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_664),
	.C2V_2 (C2V_148_664),
	.C2V_3 (C2V_242_664),
	.L (L[9959:9945]),
	.V2C_1 (V2C_664_3),
	.V2C_2 (V2C_664_148),
	.V2C_3 (V2C_664_242),
	.V (V_664)
);

VNU_3 #(quan_width) VNU665 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_665),
	.C2V_2 (C2V_154_665),
	.C2V_3 (C2V_248_665),
	.L (L[9974:9960]),
	.V2C_1 (V2C_665_9),
	.V2C_2 (V2C_665_154),
	.V2C_3 (V2C_665_248),
	.V (V_665)
);

VNU_3 #(quan_width) VNU666 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_666),
	.C2V_2 (C2V_160_666),
	.C2V_3 (C2V_254_666),
	.L (L[9989:9975]),
	.V2C_1 (V2C_666_15),
	.V2C_2 (V2C_666_160),
	.V2C_3 (V2C_666_254),
	.V (V_666)
);

VNU_3 #(quan_width) VNU667 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_667),
	.C2V_2 (C2V_166_667),
	.C2V_3 (C2V_260_667),
	.L (L[10004:9990]),
	.V2C_1 (V2C_667_21),
	.V2C_2 (V2C_667_166),
	.V2C_3 (V2C_667_260),
	.V (V_667)
);

VNU_3 #(quan_width) VNU668 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_668),
	.C2V_2 (C2V_172_668),
	.C2V_3 (C2V_266_668),
	.L (L[10019:10005]),
	.V2C_1 (V2C_668_27),
	.V2C_2 (V2C_668_172),
	.V2C_3 (V2C_668_266),
	.V (V_668)
);

VNU_3 #(quan_width) VNU669 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_669),
	.C2V_2 (C2V_178_669),
	.C2V_3 (C2V_272_669),
	.L (L[10034:10020]),
	.V2C_1 (V2C_669_33),
	.V2C_2 (V2C_669_178),
	.V2C_3 (V2C_669_272),
	.V (V_669)
);

VNU_3 #(quan_width) VNU670 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_670),
	.C2V_2 (C2V_184_670),
	.C2V_3 (C2V_278_670),
	.L (L[10049:10035]),
	.V2C_1 (V2C_670_39),
	.V2C_2 (V2C_670_184),
	.V2C_3 (V2C_670_278),
	.V (V_670)
);

VNU_3 #(quan_width) VNU671 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_671),
	.C2V_2 (C2V_190_671),
	.C2V_3 (C2V_284_671),
	.L (L[10064:10050]),
	.V2C_1 (V2C_671_45),
	.V2C_2 (V2C_671_190),
	.V2C_3 (V2C_671_284),
	.V (V_671)
);

VNU_3 #(quan_width) VNU672 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_672),
	.C2V_2 (C2V_51_672),
	.C2V_3 (C2V_196_672),
	.L (L[10079:10065]),
	.V2C_1 (V2C_672_2),
	.V2C_2 (V2C_672_51),
	.V2C_3 (V2C_672_196),
	.V (V_672)
);

VNU_3 #(quan_width) VNU673 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_214_673),
	.C2V_2 (C2V_218_673),
	.C2V_3 (C2V_287_673),
	.L (L[10094:10080]),
	.V2C_1 (V2C_673_214),
	.V2C_2 (V2C_673_218),
	.V2C_3 (V2C_673_287),
	.V (V_673)
);

VNU_3 #(quan_width) VNU674 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_674),
	.C2V_2 (C2V_220_674),
	.C2V_3 (C2V_224_674),
	.L (L[10109:10095]),
	.V2C_1 (V2C_674_5),
	.V2C_2 (V2C_674_220),
	.V2C_3 (V2C_674_224),
	.V (V_674)
);

VNU_3 #(quan_width) VNU675 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_675),
	.C2V_2 (C2V_226_675),
	.C2V_3 (C2V_230_675),
	.L (L[10124:10110]),
	.V2C_1 (V2C_675_11),
	.V2C_2 (V2C_675_226),
	.V2C_3 (V2C_675_230),
	.V (V_675)
);

VNU_3 #(quan_width) VNU676 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_676),
	.C2V_2 (C2V_232_676),
	.C2V_3 (C2V_236_676),
	.L (L[10139:10125]),
	.V2C_1 (V2C_676_17),
	.V2C_2 (V2C_676_232),
	.V2C_3 (V2C_676_236),
	.V (V_676)
);

VNU_3 #(quan_width) VNU677 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_677),
	.C2V_2 (C2V_238_677),
	.C2V_3 (C2V_242_677),
	.L (L[10154:10140]),
	.V2C_1 (V2C_677_23),
	.V2C_2 (V2C_677_238),
	.V2C_3 (V2C_677_242),
	.V (V_677)
);

VNU_3 #(quan_width) VNU678 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_678),
	.C2V_2 (C2V_244_678),
	.C2V_3 (C2V_248_678),
	.L (L[10169:10155]),
	.V2C_1 (V2C_678_29),
	.V2C_2 (V2C_678_244),
	.V2C_3 (V2C_678_248),
	.V (V_678)
);

VNU_3 #(quan_width) VNU679 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_679),
	.C2V_2 (C2V_250_679),
	.C2V_3 (C2V_254_679),
	.L (L[10184:10170]),
	.V2C_1 (V2C_679_35),
	.V2C_2 (V2C_679_250),
	.V2C_3 (V2C_679_254),
	.V (V_679)
);

VNU_3 #(quan_width) VNU680 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_680),
	.C2V_2 (C2V_256_680),
	.C2V_3 (C2V_260_680),
	.L (L[10199:10185]),
	.V2C_1 (V2C_680_41),
	.V2C_2 (V2C_680_256),
	.V2C_3 (V2C_680_260),
	.V (V_680)
);

VNU_3 #(quan_width) VNU681 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_681),
	.C2V_2 (C2V_262_681),
	.C2V_3 (C2V_266_681),
	.L (L[10214:10200]),
	.V2C_1 (V2C_681_47),
	.V2C_2 (V2C_681_262),
	.V2C_3 (V2C_681_266),
	.V (V_681)
);

VNU_3 #(quan_width) VNU682 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_682),
	.C2V_2 (C2V_268_682),
	.C2V_3 (C2V_272_682),
	.L (L[10229:10215]),
	.V2C_1 (V2C_682_53),
	.V2C_2 (V2C_682_268),
	.V2C_3 (V2C_682_272),
	.V (V_682)
);

VNU_3 #(quan_width) VNU683 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_59_683),
	.C2V_2 (C2V_274_683),
	.C2V_3 (C2V_278_683),
	.L (L[10244:10230]),
	.V2C_1 (V2C_683_59),
	.V2C_2 (V2C_683_274),
	.V2C_3 (V2C_683_278),
	.V (V_683)
);

VNU_3 #(quan_width) VNU684 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_65_684),
	.C2V_2 (C2V_280_684),
	.C2V_3 (C2V_284_684),
	.L (L[10259:10245]),
	.V2C_1 (V2C_684_65),
	.V2C_2 (V2C_684_280),
	.V2C_3 (V2C_684_284),
	.V (V_684)
);

VNU_3 #(quan_width) VNU685 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_685),
	.C2V_2 (C2V_71_685),
	.C2V_3 (C2V_286_685),
	.L (L[10274:10260]),
	.V2C_1 (V2C_685_2),
	.V2C_2 (V2C_685_71),
	.V2C_3 (V2C_685_286),
	.V (V_685)
);

VNU_3 #(quan_width) VNU686 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_686),
	.C2V_2 (C2V_8_686),
	.C2V_3 (C2V_77_686),
	.L (L[10289:10275]),
	.V2C_1 (V2C_686_4),
	.V2C_2 (V2C_686_8),
	.V2C_3 (V2C_686_77),
	.V (V_686)
);

VNU_3 #(quan_width) VNU687 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_687),
	.C2V_2 (C2V_14_687),
	.C2V_3 (C2V_83_687),
	.L (L[10304:10290]),
	.V2C_1 (V2C_687_10),
	.V2C_2 (V2C_687_14),
	.V2C_3 (V2C_687_83),
	.V (V_687)
);

VNU_3 #(quan_width) VNU688 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_688),
	.C2V_2 (C2V_20_688),
	.C2V_3 (C2V_89_688),
	.L (L[10319:10305]),
	.V2C_1 (V2C_688_16),
	.V2C_2 (V2C_688_20),
	.V2C_3 (V2C_688_89),
	.V (V_688)
);

VNU_3 #(quan_width) VNU689 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_689),
	.C2V_2 (C2V_26_689),
	.C2V_3 (C2V_95_689),
	.L (L[10334:10320]),
	.V2C_1 (V2C_689_22),
	.V2C_2 (V2C_689_26),
	.V2C_3 (V2C_689_95),
	.V (V_689)
);

VNU_3 #(quan_width) VNU690 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_690),
	.C2V_2 (C2V_32_690),
	.C2V_3 (C2V_101_690),
	.L (L[10349:10335]),
	.V2C_1 (V2C_690_28),
	.V2C_2 (V2C_690_32),
	.V2C_3 (V2C_690_101),
	.V (V_690)
);

VNU_3 #(quan_width) VNU691 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_691),
	.C2V_2 (C2V_38_691),
	.C2V_3 (C2V_107_691),
	.L (L[10364:10350]),
	.V2C_1 (V2C_691_34),
	.V2C_2 (V2C_691_38),
	.V2C_3 (V2C_691_107),
	.V (V_691)
);

VNU_3 #(quan_width) VNU692 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_692),
	.C2V_2 (C2V_44_692),
	.C2V_3 (C2V_113_692),
	.L (L[10379:10365]),
	.V2C_1 (V2C_692_40),
	.V2C_2 (V2C_692_44),
	.V2C_3 (V2C_692_113),
	.V (V_692)
);

VNU_3 #(quan_width) VNU693 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_693),
	.C2V_2 (C2V_50_693),
	.C2V_3 (C2V_119_693),
	.L (L[10394:10380]),
	.V2C_1 (V2C_693_46),
	.V2C_2 (V2C_693_50),
	.V2C_3 (V2C_693_119),
	.V (V_693)
);

VNU_3 #(quan_width) VNU694 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_694),
	.C2V_2 (C2V_56_694),
	.C2V_3 (C2V_125_694),
	.L (L[10409:10395]),
	.V2C_1 (V2C_694_52),
	.V2C_2 (V2C_694_56),
	.V2C_3 (V2C_694_125),
	.V (V_694)
);

VNU_3 #(quan_width) VNU695 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_695),
	.C2V_2 (C2V_62_695),
	.C2V_3 (C2V_131_695),
	.L (L[10424:10410]),
	.V2C_1 (V2C_695_58),
	.V2C_2 (V2C_695_62),
	.V2C_3 (V2C_695_131),
	.V (V_695)
);

VNU_3 #(quan_width) VNU696 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_696),
	.C2V_2 (C2V_68_696),
	.C2V_3 (C2V_137_696),
	.L (L[10439:10425]),
	.V2C_1 (V2C_696_64),
	.V2C_2 (V2C_696_68),
	.V2C_3 (V2C_696_137),
	.V (V_696)
);

VNU_3 #(quan_width) VNU697 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_697),
	.C2V_2 (C2V_74_697),
	.C2V_3 (C2V_143_697),
	.L (L[10454:10440]),
	.V2C_1 (V2C_697_70),
	.V2C_2 (V2C_697_74),
	.V2C_3 (V2C_697_143),
	.V (V_697)
);

VNU_3 #(quan_width) VNU698 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_698),
	.C2V_2 (C2V_80_698),
	.C2V_3 (C2V_149_698),
	.L (L[10469:10455]),
	.V2C_1 (V2C_698_76),
	.V2C_2 (V2C_698_80),
	.V2C_3 (V2C_698_149),
	.V (V_698)
);

VNU_3 #(quan_width) VNU699 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_699),
	.C2V_2 (C2V_86_699),
	.C2V_3 (C2V_155_699),
	.L (L[10484:10470]),
	.V2C_1 (V2C_699_82),
	.V2C_2 (V2C_699_86),
	.V2C_3 (V2C_699_155),
	.V (V_699)
);

VNU_3 #(quan_width) VNU700 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_700),
	.C2V_2 (C2V_92_700),
	.C2V_3 (C2V_161_700),
	.L (L[10499:10485]),
	.V2C_1 (V2C_700_88),
	.V2C_2 (V2C_700_92),
	.V2C_3 (V2C_700_161),
	.V (V_700)
);

VNU_3 #(quan_width) VNU701 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_701),
	.C2V_2 (C2V_98_701),
	.C2V_3 (C2V_167_701),
	.L (L[10514:10500]),
	.V2C_1 (V2C_701_94),
	.V2C_2 (V2C_701_98),
	.V2C_3 (V2C_701_167),
	.V (V_701)
);

VNU_3 #(quan_width) VNU702 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_702),
	.C2V_2 (C2V_104_702),
	.C2V_3 (C2V_173_702),
	.L (L[10529:10515]),
	.V2C_1 (V2C_702_100),
	.V2C_2 (V2C_702_104),
	.V2C_3 (V2C_702_173),
	.V (V_702)
);

VNU_3 #(quan_width) VNU703 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_703),
	.C2V_2 (C2V_110_703),
	.C2V_3 (C2V_179_703),
	.L (L[10544:10530]),
	.V2C_1 (V2C_703_106),
	.V2C_2 (V2C_703_110),
	.V2C_3 (V2C_703_179),
	.V (V_703)
);

VNU_3 #(quan_width) VNU704 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_704),
	.C2V_2 (C2V_116_704),
	.C2V_3 (C2V_185_704),
	.L (L[10559:10545]),
	.V2C_1 (V2C_704_112),
	.V2C_2 (V2C_704_116),
	.V2C_3 (V2C_704_185),
	.V (V_704)
);

VNU_3 #(quan_width) VNU705 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_118_705),
	.C2V_2 (C2V_122_705),
	.C2V_3 (C2V_191_705),
	.L (L[10574:10560]),
	.V2C_1 (V2C_705_118),
	.V2C_2 (V2C_705_122),
	.V2C_3 (V2C_705_191),
	.V (V_705)
);

VNU_3 #(quan_width) VNU706 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_124_706),
	.C2V_2 (C2V_128_706),
	.C2V_3 (C2V_197_706),
	.L (L[10589:10575]),
	.V2C_1 (V2C_706_124),
	.V2C_2 (V2C_706_128),
	.V2C_3 (V2C_706_197),
	.V (V_706)
);

VNU_3 #(quan_width) VNU707 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_130_707),
	.C2V_2 (C2V_134_707),
	.C2V_3 (C2V_203_707),
	.L (L[10604:10590]),
	.V2C_1 (V2C_707_130),
	.V2C_2 (V2C_707_134),
	.V2C_3 (V2C_707_203),
	.V (V_707)
);

VNU_3 #(quan_width) VNU708 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_136_708),
	.C2V_2 (C2V_140_708),
	.C2V_3 (C2V_209_708),
	.L (L[10619:10605]),
	.V2C_1 (V2C_708_136),
	.V2C_2 (V2C_708_140),
	.V2C_3 (V2C_708_209),
	.V (V_708)
);

VNU_3 #(quan_width) VNU709 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_142_709),
	.C2V_2 (C2V_146_709),
	.C2V_3 (C2V_215_709),
	.L (L[10634:10620]),
	.V2C_1 (V2C_709_142),
	.V2C_2 (V2C_709_146),
	.V2C_3 (V2C_709_215),
	.V (V_709)
);

VNU_3 #(quan_width) VNU710 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_148_710),
	.C2V_2 (C2V_152_710),
	.C2V_3 (C2V_221_710),
	.L (L[10649:10635]),
	.V2C_1 (V2C_710_148),
	.V2C_2 (V2C_710_152),
	.V2C_3 (V2C_710_221),
	.V (V_710)
);

VNU_3 #(quan_width) VNU711 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_154_711),
	.C2V_2 (C2V_158_711),
	.C2V_3 (C2V_227_711),
	.L (L[10664:10650]),
	.V2C_1 (V2C_711_154),
	.V2C_2 (V2C_711_158),
	.V2C_3 (V2C_711_227),
	.V (V_711)
);

VNU_3 #(quan_width) VNU712 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_160_712),
	.C2V_2 (C2V_164_712),
	.C2V_3 (C2V_233_712),
	.L (L[10679:10665]),
	.V2C_1 (V2C_712_160),
	.V2C_2 (V2C_712_164),
	.V2C_3 (V2C_712_233),
	.V (V_712)
);

VNU_3 #(quan_width) VNU713 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_166_713),
	.C2V_2 (C2V_170_713),
	.C2V_3 (C2V_239_713),
	.L (L[10694:10680]),
	.V2C_1 (V2C_713_166),
	.V2C_2 (V2C_713_170),
	.V2C_3 (V2C_713_239),
	.V (V_713)
);

VNU_3 #(quan_width) VNU714 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_172_714),
	.C2V_2 (C2V_176_714),
	.C2V_3 (C2V_245_714),
	.L (L[10709:10695]),
	.V2C_1 (V2C_714_172),
	.V2C_2 (V2C_714_176),
	.V2C_3 (V2C_714_245),
	.V (V_714)
);

VNU_3 #(quan_width) VNU715 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_178_715),
	.C2V_2 (C2V_182_715),
	.C2V_3 (C2V_251_715),
	.L (L[10724:10710]),
	.V2C_1 (V2C_715_178),
	.V2C_2 (V2C_715_182),
	.V2C_3 (V2C_715_251),
	.V (V_715)
);

VNU_3 #(quan_width) VNU716 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_184_716),
	.C2V_2 (C2V_188_716),
	.C2V_3 (C2V_257_716),
	.L (L[10739:10725]),
	.V2C_1 (V2C_716_184),
	.V2C_2 (V2C_716_188),
	.V2C_3 (V2C_716_257),
	.V (V_716)
);

VNU_3 #(quan_width) VNU717 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_190_717),
	.C2V_2 (C2V_194_717),
	.C2V_3 (C2V_263_717),
	.L (L[10754:10740]),
	.V2C_1 (V2C_717_190),
	.V2C_2 (V2C_717_194),
	.V2C_3 (V2C_717_263),
	.V (V_717)
);

VNU_3 #(quan_width) VNU718 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_196_718),
	.C2V_2 (C2V_200_718),
	.C2V_3 (C2V_269_718),
	.L (L[10769:10755]),
	.V2C_1 (V2C_718_196),
	.V2C_2 (V2C_718_200),
	.V2C_3 (V2C_718_269),
	.V (V_718)
);

VNU_3 #(quan_width) VNU719 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_202_719),
	.C2V_2 (C2V_206_719),
	.C2V_3 (C2V_275_719),
	.L (L[10784:10770]),
	.V2C_1 (V2C_719_202),
	.V2C_2 (V2C_719_206),
	.V2C_3 (V2C_719_275),
	.V (V_719)
);

VNU_3 #(quan_width) VNU720 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_208_720),
	.C2V_2 (C2V_212_720),
	.C2V_3 (C2V_281_720),
	.L (L[10799:10785]),
	.V2C_1 (V2C_720_208),
	.V2C_2 (V2C_720_212),
	.V2C_3 (V2C_720_281),
	.V (V_720)
);

VNU_3 #(quan_width) VNU721 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_721),
	.C2V_2 (C2V_43_721),
	.C2V_3 (C2V_191_721),
	.L (L[10814:10800]),
	.V2C_1 (V2C_721_9),
	.V2C_2 (V2C_721_43),
	.V2C_3 (V2C_721_191),
	.V (V_721)
);

VNU_3 #(quan_width) VNU722 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_722),
	.C2V_2 (C2V_49_722),
	.C2V_3 (C2V_197_722),
	.L (L[10829:10815]),
	.V2C_1 (V2C_722_15),
	.V2C_2 (V2C_722_49),
	.V2C_3 (V2C_722_197),
	.V (V_722)
);

VNU_3 #(quan_width) VNU723 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_723),
	.C2V_2 (C2V_55_723),
	.C2V_3 (C2V_203_723),
	.L (L[10844:10830]),
	.V2C_1 (V2C_723_21),
	.V2C_2 (V2C_723_55),
	.V2C_3 (V2C_723_203),
	.V (V_723)
);

VNU_3 #(quan_width) VNU724 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_724),
	.C2V_2 (C2V_61_724),
	.C2V_3 (C2V_209_724),
	.L (L[10859:10845]),
	.V2C_1 (V2C_724_27),
	.V2C_2 (V2C_724_61),
	.V2C_3 (V2C_724_209),
	.V (V_724)
);

VNU_3 #(quan_width) VNU725 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_725),
	.C2V_2 (C2V_67_725),
	.C2V_3 (C2V_215_725),
	.L (L[10874:10860]),
	.V2C_1 (V2C_725_33),
	.V2C_2 (V2C_725_67),
	.V2C_3 (V2C_725_215),
	.V (V_725)
);

VNU_3 #(quan_width) VNU726 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_726),
	.C2V_2 (C2V_73_726),
	.C2V_3 (C2V_221_726),
	.L (L[10889:10875]),
	.V2C_1 (V2C_726_39),
	.V2C_2 (V2C_726_73),
	.V2C_3 (V2C_726_221),
	.V (V_726)
);

VNU_3 #(quan_width) VNU727 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_727),
	.C2V_2 (C2V_79_727),
	.C2V_3 (C2V_227_727),
	.L (L[10904:10890]),
	.V2C_1 (V2C_727_45),
	.V2C_2 (V2C_727_79),
	.V2C_3 (V2C_727_227),
	.V (V_727)
);

VNU_3 #(quan_width) VNU728 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_728),
	.C2V_2 (C2V_85_728),
	.C2V_3 (C2V_233_728),
	.L (L[10919:10905]),
	.V2C_1 (V2C_728_51),
	.V2C_2 (V2C_728_85),
	.V2C_3 (V2C_728_233),
	.V (V_728)
);

VNU_3 #(quan_width) VNU729 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_729),
	.C2V_2 (C2V_91_729),
	.C2V_3 (C2V_239_729),
	.L (L[10934:10920]),
	.V2C_1 (V2C_729_57),
	.V2C_2 (V2C_729_91),
	.V2C_3 (V2C_729_239),
	.V (V_729)
);

VNU_3 #(quan_width) VNU730 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_730),
	.C2V_2 (C2V_97_730),
	.C2V_3 (C2V_245_730),
	.L (L[10949:10935]),
	.V2C_1 (V2C_730_63),
	.V2C_2 (V2C_730_97),
	.V2C_3 (V2C_730_245),
	.V (V_730)
);

VNU_3 #(quan_width) VNU731 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_731),
	.C2V_2 (C2V_103_731),
	.C2V_3 (C2V_251_731),
	.L (L[10964:10950]),
	.V2C_1 (V2C_731_69),
	.V2C_2 (V2C_731_103),
	.V2C_3 (V2C_731_251),
	.V (V_731)
);

VNU_3 #(quan_width) VNU732 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_732),
	.C2V_2 (C2V_109_732),
	.C2V_3 (C2V_257_732),
	.L (L[10979:10965]),
	.V2C_1 (V2C_732_75),
	.V2C_2 (V2C_732_109),
	.V2C_3 (V2C_732_257),
	.V (V_732)
);

VNU_3 #(quan_width) VNU733 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_733),
	.C2V_2 (C2V_115_733),
	.C2V_3 (C2V_263_733),
	.L (L[10994:10980]),
	.V2C_1 (V2C_733_81),
	.V2C_2 (V2C_733_115),
	.V2C_3 (V2C_733_263),
	.V (V_733)
);

VNU_3 #(quan_width) VNU734 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_734),
	.C2V_2 (C2V_121_734),
	.C2V_3 (C2V_269_734),
	.L (L[11009:10995]),
	.V2C_1 (V2C_734_87),
	.V2C_2 (V2C_734_121),
	.V2C_3 (V2C_734_269),
	.V (V_734)
);

VNU_3 #(quan_width) VNU735 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_93_735),
	.C2V_2 (C2V_127_735),
	.C2V_3 (C2V_275_735),
	.L (L[11024:11010]),
	.V2C_1 (V2C_735_93),
	.V2C_2 (V2C_735_127),
	.V2C_3 (V2C_735_275),
	.V (V_735)
);

VNU_3 #(quan_width) VNU736 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_99_736),
	.C2V_2 (C2V_133_736),
	.C2V_3 (C2V_281_736),
	.L (L[11039:11025]),
	.V2C_1 (V2C_736_99),
	.V2C_2 (V2C_736_133),
	.V2C_3 (V2C_736_281),
	.V (V_736)
);

VNU_3 #(quan_width) VNU737 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_105_737),
	.C2V_2 (C2V_139_737),
	.C2V_3 (C2V_287_737),
	.L (L[11054:11040]),
	.V2C_1 (V2C_737_105),
	.V2C_2 (V2C_737_139),
	.V2C_3 (V2C_737_287),
	.V (V_737)
);

VNU_3 #(quan_width) VNU738 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_738),
	.C2V_2 (C2V_111_738),
	.C2V_3 (C2V_145_738),
	.L (L[11069:11055]),
	.V2C_1 (V2C_738_5),
	.V2C_2 (V2C_738_111),
	.V2C_3 (V2C_738_145),
	.V (V_738)
);

VNU_3 #(quan_width) VNU739 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_739),
	.C2V_2 (C2V_117_739),
	.C2V_3 (C2V_151_739),
	.L (L[11084:11070]),
	.V2C_1 (V2C_739_11),
	.V2C_2 (V2C_739_117),
	.V2C_3 (V2C_739_151),
	.V (V_739)
);

VNU_3 #(quan_width) VNU740 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_740),
	.C2V_2 (C2V_123_740),
	.C2V_3 (C2V_157_740),
	.L (L[11099:11085]),
	.V2C_1 (V2C_740_17),
	.V2C_2 (V2C_740_123),
	.V2C_3 (V2C_740_157),
	.V (V_740)
);

VNU_3 #(quan_width) VNU741 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_741),
	.C2V_2 (C2V_129_741),
	.C2V_3 (C2V_163_741),
	.L (L[11114:11100]),
	.V2C_1 (V2C_741_23),
	.V2C_2 (V2C_741_129),
	.V2C_3 (V2C_741_163),
	.V (V_741)
);

VNU_3 #(quan_width) VNU742 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_742),
	.C2V_2 (C2V_135_742),
	.C2V_3 (C2V_169_742),
	.L (L[11129:11115]),
	.V2C_1 (V2C_742_29),
	.V2C_2 (V2C_742_135),
	.V2C_3 (V2C_742_169),
	.V (V_742)
);

VNU_3 #(quan_width) VNU743 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_743),
	.C2V_2 (C2V_141_743),
	.C2V_3 (C2V_175_743),
	.L (L[11144:11130]),
	.V2C_1 (V2C_743_35),
	.V2C_2 (V2C_743_141),
	.V2C_3 (V2C_743_175),
	.V (V_743)
);

VNU_3 #(quan_width) VNU744 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_744),
	.C2V_2 (C2V_147_744),
	.C2V_3 (C2V_181_744),
	.L (L[11159:11145]),
	.V2C_1 (V2C_744_41),
	.V2C_2 (V2C_744_147),
	.V2C_3 (V2C_744_181),
	.V (V_744)
);

VNU_3 #(quan_width) VNU745 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_745),
	.C2V_2 (C2V_153_745),
	.C2V_3 (C2V_187_745),
	.L (L[11174:11160]),
	.V2C_1 (V2C_745_47),
	.V2C_2 (V2C_745_153),
	.V2C_3 (V2C_745_187),
	.V (V_745)
);

VNU_3 #(quan_width) VNU746 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_746),
	.C2V_2 (C2V_159_746),
	.C2V_3 (C2V_193_746),
	.L (L[11189:11175]),
	.V2C_1 (V2C_746_53),
	.V2C_2 (V2C_746_159),
	.V2C_3 (V2C_746_193),
	.V (V_746)
);

VNU_3 #(quan_width) VNU747 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_59_747),
	.C2V_2 (C2V_165_747),
	.C2V_3 (C2V_199_747),
	.L (L[11204:11190]),
	.V2C_1 (V2C_747_59),
	.V2C_2 (V2C_747_165),
	.V2C_3 (V2C_747_199),
	.V (V_747)
);

VNU_3 #(quan_width) VNU748 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_65_748),
	.C2V_2 (C2V_171_748),
	.C2V_3 (C2V_205_748),
	.L (L[11219:11205]),
	.V2C_1 (V2C_748_65),
	.V2C_2 (V2C_748_171),
	.V2C_3 (V2C_748_205),
	.V (V_748)
);

VNU_3 #(quan_width) VNU749 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_71_749),
	.C2V_2 (C2V_177_749),
	.C2V_3 (C2V_211_749),
	.L (L[11234:11220]),
	.V2C_1 (V2C_749_71),
	.V2C_2 (V2C_749_177),
	.V2C_3 (V2C_749_211),
	.V (V_749)
);

VNU_3 #(quan_width) VNU750 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_77_750),
	.C2V_2 (C2V_183_750),
	.C2V_3 (C2V_217_750),
	.L (L[11249:11235]),
	.V2C_1 (V2C_750_77),
	.V2C_2 (V2C_750_183),
	.V2C_3 (V2C_750_217),
	.V (V_750)
);

VNU_3 #(quan_width) VNU751 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_83_751),
	.C2V_2 (C2V_189_751),
	.C2V_3 (C2V_223_751),
	.L (L[11264:11250]),
	.V2C_1 (V2C_751_83),
	.V2C_2 (V2C_751_189),
	.V2C_3 (V2C_751_223),
	.V (V_751)
);

VNU_3 #(quan_width) VNU752 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_89_752),
	.C2V_2 (C2V_195_752),
	.C2V_3 (C2V_229_752),
	.L (L[11279:11265]),
	.V2C_1 (V2C_752_89),
	.V2C_2 (V2C_752_195),
	.V2C_3 (V2C_752_229),
	.V (V_752)
);

VNU_3 #(quan_width) VNU753 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_95_753),
	.C2V_2 (C2V_201_753),
	.C2V_3 (C2V_235_753),
	.L (L[11294:11280]),
	.V2C_1 (V2C_753_95),
	.V2C_2 (V2C_753_201),
	.V2C_3 (V2C_753_235),
	.V (V_753)
);

VNU_3 #(quan_width) VNU754 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_101_754),
	.C2V_2 (C2V_207_754),
	.C2V_3 (C2V_241_754),
	.L (L[11309:11295]),
	.V2C_1 (V2C_754_101),
	.V2C_2 (V2C_754_207),
	.V2C_3 (V2C_754_241),
	.V (V_754)
);

VNU_3 #(quan_width) VNU755 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_107_755),
	.C2V_2 (C2V_213_755),
	.C2V_3 (C2V_247_755),
	.L (L[11324:11310]),
	.V2C_1 (V2C_755_107),
	.V2C_2 (V2C_755_213),
	.V2C_3 (V2C_755_247),
	.V (V_755)
);

VNU_3 #(quan_width) VNU756 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_113_756),
	.C2V_2 (C2V_219_756),
	.C2V_3 (C2V_253_756),
	.L (L[11339:11325]),
	.V2C_1 (V2C_756_113),
	.V2C_2 (V2C_756_219),
	.V2C_3 (V2C_756_253),
	.V (V_756)
);

VNU_3 #(quan_width) VNU757 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_119_757),
	.C2V_2 (C2V_225_757),
	.C2V_3 (C2V_259_757),
	.L (L[11354:11340]),
	.V2C_1 (V2C_757_119),
	.V2C_2 (V2C_757_225),
	.V2C_3 (V2C_757_259),
	.V (V_757)
);

VNU_3 #(quan_width) VNU758 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_125_758),
	.C2V_2 (C2V_231_758),
	.C2V_3 (C2V_265_758),
	.L (L[11369:11355]),
	.V2C_1 (V2C_758_125),
	.V2C_2 (V2C_758_231),
	.V2C_3 (V2C_758_265),
	.V (V_758)
);

VNU_3 #(quan_width) VNU759 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_131_759),
	.C2V_2 (C2V_237_759),
	.C2V_3 (C2V_271_759),
	.L (L[11384:11370]),
	.V2C_1 (V2C_759_131),
	.V2C_2 (V2C_759_237),
	.V2C_3 (V2C_759_271),
	.V (V_759)
);

VNU_3 #(quan_width) VNU760 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_137_760),
	.C2V_2 (C2V_243_760),
	.C2V_3 (C2V_277_760),
	.L (L[11399:11385]),
	.V2C_1 (V2C_760_137),
	.V2C_2 (V2C_760_243),
	.V2C_3 (V2C_760_277),
	.V (V_760)
);

VNU_3 #(quan_width) VNU761 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_143_761),
	.C2V_2 (C2V_249_761),
	.C2V_3 (C2V_283_761),
	.L (L[11414:11400]),
	.V2C_1 (V2C_761_143),
	.V2C_2 (V2C_761_249),
	.V2C_3 (V2C_761_283),
	.V (V_761)
);

VNU_3 #(quan_width) VNU762 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_762),
	.C2V_2 (C2V_149_762),
	.C2V_3 (C2V_255_762),
	.L (L[11429:11415]),
	.V2C_1 (V2C_762_1),
	.V2C_2 (V2C_762_149),
	.V2C_3 (V2C_762_255),
	.V (V_762)
);

VNU_3 #(quan_width) VNU763 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_763),
	.C2V_2 (C2V_155_763),
	.C2V_3 (C2V_261_763),
	.L (L[11444:11430]),
	.V2C_1 (V2C_763_7),
	.V2C_2 (V2C_763_155),
	.V2C_3 (V2C_763_261),
	.V (V_763)
);

VNU_3 #(quan_width) VNU764 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_764),
	.C2V_2 (C2V_161_764),
	.C2V_3 (C2V_267_764),
	.L (L[11459:11445]),
	.V2C_1 (V2C_764_13),
	.V2C_2 (V2C_764_161),
	.V2C_3 (V2C_764_267),
	.V (V_764)
);

VNU_3 #(quan_width) VNU765 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_765),
	.C2V_2 (C2V_167_765),
	.C2V_3 (C2V_273_765),
	.L (L[11474:11460]),
	.V2C_1 (V2C_765_19),
	.V2C_2 (V2C_765_167),
	.V2C_3 (V2C_765_273),
	.V (V_765)
);

VNU_3 #(quan_width) VNU766 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_766),
	.C2V_2 (C2V_173_766),
	.C2V_3 (C2V_279_766),
	.L (L[11489:11475]),
	.V2C_1 (V2C_766_25),
	.V2C_2 (V2C_766_173),
	.V2C_3 (V2C_766_279),
	.V (V_766)
);

VNU_3 #(quan_width) VNU767 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_767),
	.C2V_2 (C2V_179_767),
	.C2V_3 (C2V_285_767),
	.L (L[11504:11490]),
	.V2C_1 (V2C_767_31),
	.V2C_2 (V2C_767_179),
	.V2C_3 (V2C_767_285),
	.V (V_767)
);

VNU_3 #(quan_width) VNU768 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_768),
	.C2V_2 (C2V_37_768),
	.C2V_3 (C2V_185_768),
	.L (L[11519:11505]),
	.V2C_1 (V2C_768_3),
	.V2C_2 (V2C_768_37),
	.V2C_3 (V2C_768_185),
	.V (V_768)
);

VNU_3 #(quan_width) VNU769 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_769),
	.C2V_2 (C2V_43_769),
	.C2V_3 (C2V_155_769),
	.L (L[11534:11520]),
	.V2C_1 (V2C_769_24),
	.V2C_2 (V2C_769_43),
	.V2C_3 (V2C_769_155),
	.V (V_769)
);

VNU_3 #(quan_width) VNU770 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_770),
	.C2V_2 (C2V_49_770),
	.C2V_3 (C2V_161_770),
	.L (L[11549:11535]),
	.V2C_1 (V2C_770_30),
	.V2C_2 (V2C_770_49),
	.V2C_3 (V2C_770_161),
	.V (V_770)
);

VNU_3 #(quan_width) VNU771 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_771),
	.C2V_2 (C2V_55_771),
	.C2V_3 (C2V_167_771),
	.L (L[11564:11550]),
	.V2C_1 (V2C_771_36),
	.V2C_2 (V2C_771_55),
	.V2C_3 (V2C_771_167),
	.V (V_771)
);

VNU_3 #(quan_width) VNU772 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_772),
	.C2V_2 (C2V_61_772),
	.C2V_3 (C2V_173_772),
	.L (L[11579:11565]),
	.V2C_1 (V2C_772_42),
	.V2C_2 (V2C_772_61),
	.V2C_3 (V2C_772_173),
	.V (V_772)
);

VNU_3 #(quan_width) VNU773 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_773),
	.C2V_2 (C2V_67_773),
	.C2V_3 (C2V_179_773),
	.L (L[11594:11580]),
	.V2C_1 (V2C_773_48),
	.V2C_2 (V2C_773_67),
	.V2C_3 (V2C_773_179),
	.V (V_773)
);

VNU_3 #(quan_width) VNU774 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_54_774),
	.C2V_2 (C2V_73_774),
	.C2V_3 (C2V_185_774),
	.L (L[11609:11595]),
	.V2C_1 (V2C_774_54),
	.V2C_2 (V2C_774_73),
	.V2C_3 (V2C_774_185),
	.V (V_774)
);

VNU_3 #(quan_width) VNU775 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_60_775),
	.C2V_2 (C2V_79_775),
	.C2V_3 (C2V_191_775),
	.L (L[11624:11610]),
	.V2C_1 (V2C_775_60),
	.V2C_2 (V2C_775_79),
	.V2C_3 (V2C_775_191),
	.V (V_775)
);

VNU_3 #(quan_width) VNU776 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_66_776),
	.C2V_2 (C2V_85_776),
	.C2V_3 (C2V_197_776),
	.L (L[11639:11625]),
	.V2C_1 (V2C_776_66),
	.V2C_2 (V2C_776_85),
	.V2C_3 (V2C_776_197),
	.V (V_776)
);

VNU_3 #(quan_width) VNU777 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_72_777),
	.C2V_2 (C2V_91_777),
	.C2V_3 (C2V_203_777),
	.L (L[11654:11640]),
	.V2C_1 (V2C_777_72),
	.V2C_2 (V2C_777_91),
	.V2C_3 (V2C_777_203),
	.V (V_777)
);

VNU_3 #(quan_width) VNU778 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_78_778),
	.C2V_2 (C2V_97_778),
	.C2V_3 (C2V_209_778),
	.L (L[11669:11655]),
	.V2C_1 (V2C_778_78),
	.V2C_2 (V2C_778_97),
	.V2C_3 (V2C_778_209),
	.V (V_778)
);

VNU_3 #(quan_width) VNU779 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_84_779),
	.C2V_2 (C2V_103_779),
	.C2V_3 (C2V_215_779),
	.L (L[11684:11670]),
	.V2C_1 (V2C_779_84),
	.V2C_2 (V2C_779_103),
	.V2C_3 (V2C_779_215),
	.V (V_779)
);

VNU_3 #(quan_width) VNU780 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_90_780),
	.C2V_2 (C2V_109_780),
	.C2V_3 (C2V_221_780),
	.L (L[11699:11685]),
	.V2C_1 (V2C_780_90),
	.V2C_2 (V2C_780_109),
	.V2C_3 (V2C_780_221),
	.V (V_780)
);

VNU_3 #(quan_width) VNU781 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_96_781),
	.C2V_2 (C2V_115_781),
	.C2V_3 (C2V_227_781),
	.L (L[11714:11700]),
	.V2C_1 (V2C_781_96),
	.V2C_2 (V2C_781_115),
	.V2C_3 (V2C_781_227),
	.V (V_781)
);

VNU_3 #(quan_width) VNU782 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_102_782),
	.C2V_2 (C2V_121_782),
	.C2V_3 (C2V_233_782),
	.L (L[11729:11715]),
	.V2C_1 (V2C_782_102),
	.V2C_2 (V2C_782_121),
	.V2C_3 (V2C_782_233),
	.V (V_782)
);

VNU_3 #(quan_width) VNU783 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_108_783),
	.C2V_2 (C2V_127_783),
	.C2V_3 (C2V_239_783),
	.L (L[11744:11730]),
	.V2C_1 (V2C_783_108),
	.V2C_2 (V2C_783_127),
	.V2C_3 (V2C_783_239),
	.V (V_783)
);

VNU_3 #(quan_width) VNU784 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_114_784),
	.C2V_2 (C2V_133_784),
	.C2V_3 (C2V_245_784),
	.L (L[11759:11745]),
	.V2C_1 (V2C_784_114),
	.V2C_2 (V2C_784_133),
	.V2C_3 (V2C_784_245),
	.V (V_784)
);

VNU_3 #(quan_width) VNU785 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_120_785),
	.C2V_2 (C2V_139_785),
	.C2V_3 (C2V_251_785),
	.L (L[11774:11760]),
	.V2C_1 (V2C_785_120),
	.V2C_2 (V2C_785_139),
	.V2C_3 (V2C_785_251),
	.V (V_785)
);

VNU_3 #(quan_width) VNU786 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_126_786),
	.C2V_2 (C2V_145_786),
	.C2V_3 (C2V_257_786),
	.L (L[11789:11775]),
	.V2C_1 (V2C_786_126),
	.V2C_2 (V2C_786_145),
	.V2C_3 (V2C_786_257),
	.V (V_786)
);

VNU_3 #(quan_width) VNU787 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_132_787),
	.C2V_2 (C2V_151_787),
	.C2V_3 (C2V_263_787),
	.L (L[11804:11790]),
	.V2C_1 (V2C_787_132),
	.V2C_2 (V2C_787_151),
	.V2C_3 (V2C_787_263),
	.V (V_787)
);

VNU_3 #(quan_width) VNU788 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_138_788),
	.C2V_2 (C2V_157_788),
	.C2V_3 (C2V_269_788),
	.L (L[11819:11805]),
	.V2C_1 (V2C_788_138),
	.V2C_2 (V2C_788_157),
	.V2C_3 (V2C_788_269),
	.V (V_788)
);

VNU_3 #(quan_width) VNU789 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_144_789),
	.C2V_2 (C2V_163_789),
	.C2V_3 (C2V_275_789),
	.L (L[11834:11820]),
	.V2C_1 (V2C_789_144),
	.V2C_2 (V2C_789_163),
	.V2C_3 (V2C_789_275),
	.V (V_789)
);

VNU_3 #(quan_width) VNU790 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_150_790),
	.C2V_2 (C2V_169_790),
	.C2V_3 (C2V_281_790),
	.L (L[11849:11835]),
	.V2C_1 (V2C_790_150),
	.V2C_2 (V2C_790_169),
	.V2C_3 (V2C_790_281),
	.V (V_790)
);

VNU_3 #(quan_width) VNU791 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_156_791),
	.C2V_2 (C2V_175_791),
	.C2V_3 (C2V_287_791),
	.L (L[11864:11850]),
	.V2C_1 (V2C_791_156),
	.V2C_2 (V2C_791_175),
	.V2C_3 (V2C_791_287),
	.V (V_791)
);

VNU_3 #(quan_width) VNU792 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_792),
	.C2V_2 (C2V_162_792),
	.C2V_3 (C2V_181_792),
	.L (L[11879:11865]),
	.V2C_1 (V2C_792_5),
	.V2C_2 (V2C_792_162),
	.V2C_3 (V2C_792_181),
	.V (V_792)
);

VNU_3 #(quan_width) VNU793 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_793),
	.C2V_2 (C2V_168_793),
	.C2V_3 (C2V_187_793),
	.L (L[11894:11880]),
	.V2C_1 (V2C_793_11),
	.V2C_2 (V2C_793_168),
	.V2C_3 (V2C_793_187),
	.V (V_793)
);

VNU_3 #(quan_width) VNU794 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_794),
	.C2V_2 (C2V_174_794),
	.C2V_3 (C2V_193_794),
	.L (L[11909:11895]),
	.V2C_1 (V2C_794_17),
	.V2C_2 (V2C_794_174),
	.V2C_3 (V2C_794_193),
	.V (V_794)
);

VNU_3 #(quan_width) VNU795 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_795),
	.C2V_2 (C2V_180_795),
	.C2V_3 (C2V_199_795),
	.L (L[11924:11910]),
	.V2C_1 (V2C_795_23),
	.V2C_2 (V2C_795_180),
	.V2C_3 (V2C_795_199),
	.V (V_795)
);

VNU_3 #(quan_width) VNU796 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_796),
	.C2V_2 (C2V_186_796),
	.C2V_3 (C2V_205_796),
	.L (L[11939:11925]),
	.V2C_1 (V2C_796_29),
	.V2C_2 (V2C_796_186),
	.V2C_3 (V2C_796_205),
	.V (V_796)
);

VNU_3 #(quan_width) VNU797 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_797),
	.C2V_2 (C2V_192_797),
	.C2V_3 (C2V_211_797),
	.L (L[11954:11940]),
	.V2C_1 (V2C_797_35),
	.V2C_2 (V2C_797_192),
	.V2C_3 (V2C_797_211),
	.V (V_797)
);

VNU_3 #(quan_width) VNU798 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_798),
	.C2V_2 (C2V_198_798),
	.C2V_3 (C2V_217_798),
	.L (L[11969:11955]),
	.V2C_1 (V2C_798_41),
	.V2C_2 (V2C_798_198),
	.V2C_3 (V2C_798_217),
	.V (V_798)
);

VNU_3 #(quan_width) VNU799 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_799),
	.C2V_2 (C2V_204_799),
	.C2V_3 (C2V_223_799),
	.L (L[11984:11970]),
	.V2C_1 (V2C_799_47),
	.V2C_2 (V2C_799_204),
	.V2C_3 (V2C_799_223),
	.V (V_799)
);

VNU_3 #(quan_width) VNU800 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_800),
	.C2V_2 (C2V_210_800),
	.C2V_3 (C2V_229_800),
	.L (L[11999:11985]),
	.V2C_1 (V2C_800_53),
	.V2C_2 (V2C_800_210),
	.V2C_3 (V2C_800_229),
	.V (V_800)
);

VNU_3 #(quan_width) VNU801 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_59_801),
	.C2V_2 (C2V_216_801),
	.C2V_3 (C2V_235_801),
	.L (L[12014:12000]),
	.V2C_1 (V2C_801_59),
	.V2C_2 (V2C_801_216),
	.V2C_3 (V2C_801_235),
	.V (V_801)
);

VNU_3 #(quan_width) VNU802 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_65_802),
	.C2V_2 (C2V_222_802),
	.C2V_3 (C2V_241_802),
	.L (L[12029:12015]),
	.V2C_1 (V2C_802_65),
	.V2C_2 (V2C_802_222),
	.V2C_3 (V2C_802_241),
	.V (V_802)
);

VNU_3 #(quan_width) VNU803 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_71_803),
	.C2V_2 (C2V_228_803),
	.C2V_3 (C2V_247_803),
	.L (L[12044:12030]),
	.V2C_1 (V2C_803_71),
	.V2C_2 (V2C_803_228),
	.V2C_3 (V2C_803_247),
	.V (V_803)
);

VNU_3 #(quan_width) VNU804 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_77_804),
	.C2V_2 (C2V_234_804),
	.C2V_3 (C2V_253_804),
	.L (L[12059:12045]),
	.V2C_1 (V2C_804_77),
	.V2C_2 (V2C_804_234),
	.V2C_3 (V2C_804_253),
	.V (V_804)
);

VNU_3 #(quan_width) VNU805 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_83_805),
	.C2V_2 (C2V_240_805),
	.C2V_3 (C2V_259_805),
	.L (L[12074:12060]),
	.V2C_1 (V2C_805_83),
	.V2C_2 (V2C_805_240),
	.V2C_3 (V2C_805_259),
	.V (V_805)
);

VNU_3 #(quan_width) VNU806 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_89_806),
	.C2V_2 (C2V_246_806),
	.C2V_3 (C2V_265_806),
	.L (L[12089:12075]),
	.V2C_1 (V2C_806_89),
	.V2C_2 (V2C_806_246),
	.V2C_3 (V2C_806_265),
	.V (V_806)
);

VNU_3 #(quan_width) VNU807 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_95_807),
	.C2V_2 (C2V_252_807),
	.C2V_3 (C2V_271_807),
	.L (L[12104:12090]),
	.V2C_1 (V2C_807_95),
	.V2C_2 (V2C_807_252),
	.V2C_3 (V2C_807_271),
	.V (V_807)
);

VNU_3 #(quan_width) VNU808 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_101_808),
	.C2V_2 (C2V_258_808),
	.C2V_3 (C2V_277_808),
	.L (L[12119:12105]),
	.V2C_1 (V2C_808_101),
	.V2C_2 (V2C_808_258),
	.V2C_3 (V2C_808_277),
	.V (V_808)
);

VNU_3 #(quan_width) VNU809 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_107_809),
	.C2V_2 (C2V_264_809),
	.C2V_3 (C2V_283_809),
	.L (L[12134:12120]),
	.V2C_1 (V2C_809_107),
	.V2C_2 (V2C_809_264),
	.V2C_3 (V2C_809_283),
	.V (V_809)
);

VNU_3 #(quan_width) VNU810 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_810),
	.C2V_2 (C2V_113_810),
	.C2V_3 (C2V_270_810),
	.L (L[12149:12135]),
	.V2C_1 (V2C_810_1),
	.V2C_2 (V2C_810_113),
	.V2C_3 (V2C_810_270),
	.V (V_810)
);

VNU_3 #(quan_width) VNU811 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_811),
	.C2V_2 (C2V_119_811),
	.C2V_3 (C2V_276_811),
	.L (L[12164:12150]),
	.V2C_1 (V2C_811_7),
	.V2C_2 (V2C_811_119),
	.V2C_3 (V2C_811_276),
	.V (V_811)
);

VNU_3 #(quan_width) VNU812 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_812),
	.C2V_2 (C2V_125_812),
	.C2V_3 (C2V_282_812),
	.L (L[12179:12165]),
	.V2C_1 (V2C_812_13),
	.V2C_2 (V2C_812_125),
	.V2C_3 (V2C_812_282),
	.V (V_812)
);

VNU_3 #(quan_width) VNU813 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_813),
	.C2V_2 (C2V_131_813),
	.C2V_3 (C2V_288_813),
	.L (L[12194:12180]),
	.V2C_1 (V2C_813_19),
	.V2C_2 (V2C_813_131),
	.V2C_3 (V2C_813_288),
	.V (V_813)
);

VNU_3 #(quan_width) VNU814 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_814),
	.C2V_2 (C2V_25_814),
	.C2V_3 (C2V_137_814),
	.L (L[12209:12195]),
	.V2C_1 (V2C_814_6),
	.V2C_2 (V2C_814_25),
	.V2C_3 (V2C_814_137),
	.V (V_814)
);

VNU_3 #(quan_width) VNU815 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_815),
	.C2V_2 (C2V_31_815),
	.C2V_3 (C2V_143_815),
	.L (L[12224:12210]),
	.V2C_1 (V2C_815_12),
	.V2C_2 (V2C_815_31),
	.V2C_3 (V2C_815_143),
	.V (V_815)
);

VNU_3 #(quan_width) VNU816 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_816),
	.C2V_2 (C2V_37_816),
	.C2V_3 (C2V_149_816),
	.L (L[12239:12225]),
	.V2C_1 (V2C_816_18),
	.V2C_2 (V2C_816_37),
	.V2C_3 (V2C_816_149),
	.V (V_816)
);

VNU_3 #(quan_width) VNU817 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_817),
	.C2V_2 (C2V_74_817),
	.C2V_3 (C2V_144_817),
	.L (L[12254:12240]),
	.V2C_1 (V2C_817_43),
	.V2C_2 (V2C_817_74),
	.V2C_3 (V2C_817_144),
	.V (V_817)
);

VNU_3 #(quan_width) VNU818 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_818),
	.C2V_2 (C2V_80_818),
	.C2V_3 (C2V_150_818),
	.L (L[12269:12255]),
	.V2C_1 (V2C_818_49),
	.V2C_2 (V2C_818_80),
	.V2C_3 (V2C_818_150),
	.V (V_818)
);

VNU_3 #(quan_width) VNU819 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_819),
	.C2V_2 (C2V_86_819),
	.C2V_3 (C2V_156_819),
	.L (L[12284:12270]),
	.V2C_1 (V2C_819_55),
	.V2C_2 (V2C_819_86),
	.V2C_3 (V2C_819_156),
	.V (V_819)
);

VNU_3 #(quan_width) VNU820 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_820),
	.C2V_2 (C2V_92_820),
	.C2V_3 (C2V_162_820),
	.L (L[12299:12285]),
	.V2C_1 (V2C_820_61),
	.V2C_2 (V2C_820_92),
	.V2C_3 (V2C_820_162),
	.V (V_820)
);

VNU_3 #(quan_width) VNU821 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_821),
	.C2V_2 (C2V_98_821),
	.C2V_3 (C2V_168_821),
	.L (L[12314:12300]),
	.V2C_1 (V2C_821_67),
	.V2C_2 (V2C_821_98),
	.V2C_3 (V2C_821_168),
	.V (V_821)
);

VNU_3 #(quan_width) VNU822 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_822),
	.C2V_2 (C2V_104_822),
	.C2V_3 (C2V_174_822),
	.L (L[12329:12315]),
	.V2C_1 (V2C_822_73),
	.V2C_2 (V2C_822_104),
	.V2C_3 (V2C_822_174),
	.V (V_822)
);

VNU_3 #(quan_width) VNU823 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_823),
	.C2V_2 (C2V_110_823),
	.C2V_3 (C2V_180_823),
	.L (L[12344:12330]),
	.V2C_1 (V2C_823_79),
	.V2C_2 (V2C_823_110),
	.V2C_3 (V2C_823_180),
	.V (V_823)
);

VNU_3 #(quan_width) VNU824 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_824),
	.C2V_2 (C2V_116_824),
	.C2V_3 (C2V_186_824),
	.L (L[12359:12345]),
	.V2C_1 (V2C_824_85),
	.V2C_2 (V2C_824_116),
	.V2C_3 (V2C_824_186),
	.V (V_824)
);

VNU_3 #(quan_width) VNU825 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_91_825),
	.C2V_2 (C2V_122_825),
	.C2V_3 (C2V_192_825),
	.L (L[12374:12360]),
	.V2C_1 (V2C_825_91),
	.V2C_2 (V2C_825_122),
	.V2C_3 (V2C_825_192),
	.V (V_825)
);

VNU_3 #(quan_width) VNU826 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_97_826),
	.C2V_2 (C2V_128_826),
	.C2V_3 (C2V_198_826),
	.L (L[12389:12375]),
	.V2C_1 (V2C_826_97),
	.V2C_2 (V2C_826_128),
	.V2C_3 (V2C_826_198),
	.V (V_826)
);

VNU_3 #(quan_width) VNU827 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_103_827),
	.C2V_2 (C2V_134_827),
	.C2V_3 (C2V_204_827),
	.L (L[12404:12390]),
	.V2C_1 (V2C_827_103),
	.V2C_2 (V2C_827_134),
	.V2C_3 (V2C_827_204),
	.V (V_827)
);

VNU_3 #(quan_width) VNU828 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_109_828),
	.C2V_2 (C2V_140_828),
	.C2V_3 (C2V_210_828),
	.L (L[12419:12405]),
	.V2C_1 (V2C_828_109),
	.V2C_2 (V2C_828_140),
	.V2C_3 (V2C_828_210),
	.V (V_828)
);

VNU_3 #(quan_width) VNU829 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_115_829),
	.C2V_2 (C2V_146_829),
	.C2V_3 (C2V_216_829),
	.L (L[12434:12420]),
	.V2C_1 (V2C_829_115),
	.V2C_2 (V2C_829_146),
	.V2C_3 (V2C_829_216),
	.V (V_829)
);

VNU_3 #(quan_width) VNU830 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_121_830),
	.C2V_2 (C2V_152_830),
	.C2V_3 (C2V_222_830),
	.L (L[12449:12435]),
	.V2C_1 (V2C_830_121),
	.V2C_2 (V2C_830_152),
	.V2C_3 (V2C_830_222),
	.V (V_830)
);

VNU_3 #(quan_width) VNU831 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_127_831),
	.C2V_2 (C2V_158_831),
	.C2V_3 (C2V_228_831),
	.L (L[12464:12450]),
	.V2C_1 (V2C_831_127),
	.V2C_2 (V2C_831_158),
	.V2C_3 (V2C_831_228),
	.V (V_831)
);

VNU_3 #(quan_width) VNU832 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_133_832),
	.C2V_2 (C2V_164_832),
	.C2V_3 (C2V_234_832),
	.L (L[12479:12465]),
	.V2C_1 (V2C_832_133),
	.V2C_2 (V2C_832_164),
	.V2C_3 (V2C_832_234),
	.V (V_832)
);

VNU_3 #(quan_width) VNU833 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_139_833),
	.C2V_2 (C2V_170_833),
	.C2V_3 (C2V_240_833),
	.L (L[12494:12480]),
	.V2C_1 (V2C_833_139),
	.V2C_2 (V2C_833_170),
	.V2C_3 (V2C_833_240),
	.V (V_833)
);

VNU_3 #(quan_width) VNU834 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_145_834),
	.C2V_2 (C2V_176_834),
	.C2V_3 (C2V_246_834),
	.L (L[12509:12495]),
	.V2C_1 (V2C_834_145),
	.V2C_2 (V2C_834_176),
	.V2C_3 (V2C_834_246),
	.V (V_834)
);

VNU_3 #(quan_width) VNU835 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_151_835),
	.C2V_2 (C2V_182_835),
	.C2V_3 (C2V_252_835),
	.L (L[12524:12510]),
	.V2C_1 (V2C_835_151),
	.V2C_2 (V2C_835_182),
	.V2C_3 (V2C_835_252),
	.V (V_835)
);

VNU_3 #(quan_width) VNU836 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_157_836),
	.C2V_2 (C2V_188_836),
	.C2V_3 (C2V_258_836),
	.L (L[12539:12525]),
	.V2C_1 (V2C_836_157),
	.V2C_2 (V2C_836_188),
	.V2C_3 (V2C_836_258),
	.V (V_836)
);

VNU_3 #(quan_width) VNU837 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_163_837),
	.C2V_2 (C2V_194_837),
	.C2V_3 (C2V_264_837),
	.L (L[12554:12540]),
	.V2C_1 (V2C_837_163),
	.V2C_2 (V2C_837_194),
	.V2C_3 (V2C_837_264),
	.V (V_837)
);

VNU_3 #(quan_width) VNU838 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_169_838),
	.C2V_2 (C2V_200_838),
	.C2V_3 (C2V_270_838),
	.L (L[12569:12555]),
	.V2C_1 (V2C_838_169),
	.V2C_2 (V2C_838_200),
	.V2C_3 (V2C_838_270),
	.V (V_838)
);

VNU_3 #(quan_width) VNU839 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_175_839),
	.C2V_2 (C2V_206_839),
	.C2V_3 (C2V_276_839),
	.L (L[12584:12570]),
	.V2C_1 (V2C_839_175),
	.V2C_2 (V2C_839_206),
	.V2C_3 (V2C_839_276),
	.V (V_839)
);

VNU_3 #(quan_width) VNU840 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_181_840),
	.C2V_2 (C2V_212_840),
	.C2V_3 (C2V_282_840),
	.L (L[12599:12585]),
	.V2C_1 (V2C_840_181),
	.V2C_2 (V2C_840_212),
	.V2C_3 (V2C_840_282),
	.V (V_840)
);

VNU_3 #(quan_width) VNU841 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_187_841),
	.C2V_2 (C2V_218_841),
	.C2V_3 (C2V_288_841),
	.L (L[12614:12600]),
	.V2C_1 (V2C_841_187),
	.V2C_2 (V2C_841_218),
	.V2C_3 (V2C_841_288),
	.V (V_841)
);

VNU_3 #(quan_width) VNU842 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_842),
	.C2V_2 (C2V_193_842),
	.C2V_3 (C2V_224_842),
	.L (L[12629:12615]),
	.V2C_1 (V2C_842_6),
	.V2C_2 (V2C_842_193),
	.V2C_3 (V2C_842_224),
	.V (V_842)
);

VNU_3 #(quan_width) VNU843 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_843),
	.C2V_2 (C2V_199_843),
	.C2V_3 (C2V_230_843),
	.L (L[12644:12630]),
	.V2C_1 (V2C_843_12),
	.V2C_2 (V2C_843_199),
	.V2C_3 (V2C_843_230),
	.V (V_843)
);

VNU_3 #(quan_width) VNU844 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_844),
	.C2V_2 (C2V_205_844),
	.C2V_3 (C2V_236_844),
	.L (L[12659:12645]),
	.V2C_1 (V2C_844_18),
	.V2C_2 (V2C_844_205),
	.V2C_3 (V2C_844_236),
	.V (V_844)
);

VNU_3 #(quan_width) VNU845 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_845),
	.C2V_2 (C2V_211_845),
	.C2V_3 (C2V_242_845),
	.L (L[12674:12660]),
	.V2C_1 (V2C_845_24),
	.V2C_2 (V2C_845_211),
	.V2C_3 (V2C_845_242),
	.V (V_845)
);

VNU_3 #(quan_width) VNU846 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_846),
	.C2V_2 (C2V_217_846),
	.C2V_3 (C2V_248_846),
	.L (L[12689:12675]),
	.V2C_1 (V2C_846_30),
	.V2C_2 (V2C_846_217),
	.V2C_3 (V2C_846_248),
	.V (V_846)
);

VNU_3 #(quan_width) VNU847 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_847),
	.C2V_2 (C2V_223_847),
	.C2V_3 (C2V_254_847),
	.L (L[12704:12690]),
	.V2C_1 (V2C_847_36),
	.V2C_2 (V2C_847_223),
	.V2C_3 (V2C_847_254),
	.V (V_847)
);

VNU_3 #(quan_width) VNU848 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_848),
	.C2V_2 (C2V_229_848),
	.C2V_3 (C2V_260_848),
	.L (L[12719:12705]),
	.V2C_1 (V2C_848_42),
	.V2C_2 (V2C_848_229),
	.V2C_3 (V2C_848_260),
	.V (V_848)
);

VNU_3 #(quan_width) VNU849 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_849),
	.C2V_2 (C2V_235_849),
	.C2V_3 (C2V_266_849),
	.L (L[12734:12720]),
	.V2C_1 (V2C_849_48),
	.V2C_2 (V2C_849_235),
	.V2C_3 (V2C_849_266),
	.V (V_849)
);

VNU_3 #(quan_width) VNU850 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_54_850),
	.C2V_2 (C2V_241_850),
	.C2V_3 (C2V_272_850),
	.L (L[12749:12735]),
	.V2C_1 (V2C_850_54),
	.V2C_2 (V2C_850_241),
	.V2C_3 (V2C_850_272),
	.V (V_850)
);

VNU_3 #(quan_width) VNU851 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_60_851),
	.C2V_2 (C2V_247_851),
	.C2V_3 (C2V_278_851),
	.L (L[12764:12750]),
	.V2C_1 (V2C_851_60),
	.V2C_2 (V2C_851_247),
	.V2C_3 (V2C_851_278),
	.V (V_851)
);

VNU_3 #(quan_width) VNU852 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_66_852),
	.C2V_2 (C2V_253_852),
	.C2V_3 (C2V_284_852),
	.L (L[12779:12765]),
	.V2C_1 (V2C_852_66),
	.V2C_2 (V2C_852_253),
	.V2C_3 (V2C_852_284),
	.V (V_852)
);

VNU_3 #(quan_width) VNU853 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_853),
	.C2V_2 (C2V_72_853),
	.C2V_3 (C2V_259_853),
	.L (L[12794:12780]),
	.V2C_1 (V2C_853_2),
	.V2C_2 (V2C_853_72),
	.V2C_3 (V2C_853_259),
	.V (V_853)
);

VNU_3 #(quan_width) VNU854 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_854),
	.C2V_2 (C2V_78_854),
	.C2V_3 (C2V_265_854),
	.L (L[12809:12795]),
	.V2C_1 (V2C_854_8),
	.V2C_2 (V2C_854_78),
	.V2C_3 (V2C_854_265),
	.V (V_854)
);

VNU_3 #(quan_width) VNU855 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_855),
	.C2V_2 (C2V_84_855),
	.C2V_3 (C2V_271_855),
	.L (L[12824:12810]),
	.V2C_1 (V2C_855_14),
	.V2C_2 (V2C_855_84),
	.V2C_3 (V2C_855_271),
	.V (V_855)
);

VNU_3 #(quan_width) VNU856 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_856),
	.C2V_2 (C2V_90_856),
	.C2V_3 (C2V_277_856),
	.L (L[12839:12825]),
	.V2C_1 (V2C_856_20),
	.V2C_2 (V2C_856_90),
	.V2C_3 (V2C_856_277),
	.V (V_856)
);

VNU_3 #(quan_width) VNU857 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_857),
	.C2V_2 (C2V_96_857),
	.C2V_3 (C2V_283_857),
	.L (L[12854:12840]),
	.V2C_1 (V2C_857_26),
	.V2C_2 (V2C_857_96),
	.V2C_3 (V2C_857_283),
	.V (V_857)
);

VNU_3 #(quan_width) VNU858 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_858),
	.C2V_2 (C2V_32_858),
	.C2V_3 (C2V_102_858),
	.L (L[12869:12855]),
	.V2C_1 (V2C_858_1),
	.V2C_2 (V2C_858_32),
	.V2C_3 (V2C_858_102),
	.V (V_858)
);

VNU_3 #(quan_width) VNU859 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_859),
	.C2V_2 (C2V_38_859),
	.C2V_3 (C2V_108_859),
	.L (L[12884:12870]),
	.V2C_1 (V2C_859_7),
	.V2C_2 (V2C_859_38),
	.V2C_3 (V2C_859_108),
	.V (V_859)
);

VNU_3 #(quan_width) VNU860 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_860),
	.C2V_2 (C2V_44_860),
	.C2V_3 (C2V_114_860),
	.L (L[12899:12885]),
	.V2C_1 (V2C_860_13),
	.V2C_2 (V2C_860_44),
	.V2C_3 (V2C_860_114),
	.V (V_860)
);

VNU_3 #(quan_width) VNU861 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_861),
	.C2V_2 (C2V_50_861),
	.C2V_3 (C2V_120_861),
	.L (L[12914:12900]),
	.V2C_1 (V2C_861_19),
	.V2C_2 (V2C_861_50),
	.V2C_3 (V2C_861_120),
	.V (V_861)
);

VNU_3 #(quan_width) VNU862 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_862),
	.C2V_2 (C2V_56_862),
	.C2V_3 (C2V_126_862),
	.L (L[12929:12915]),
	.V2C_1 (V2C_862_25),
	.V2C_2 (V2C_862_56),
	.V2C_3 (V2C_862_126),
	.V (V_862)
);

VNU_3 #(quan_width) VNU863 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_863),
	.C2V_2 (C2V_62_863),
	.C2V_3 (C2V_132_863),
	.L (L[12944:12930]),
	.V2C_1 (V2C_863_31),
	.V2C_2 (V2C_863_62),
	.V2C_3 (V2C_863_132),
	.V (V_863)
);

VNU_3 #(quan_width) VNU864 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_864),
	.C2V_2 (C2V_68_864),
	.C2V_3 (C2V_138_864),
	.L (L[12959:12945]),
	.V2C_1 (V2C_864_37),
	.V2C_2 (V2C_864_68),
	.V2C_3 (V2C_864_138),
	.V (V_864)
);

VNU_6 #(quan_width) VNU865 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_865),
	.C2V_2 (C2V_85_865),
	.C2V_3 (C2V_87_865),
	.C2V_4 (C2V_110_865),
	.C2V_5 (C2V_234_865),
	.C2V_6 (C2V_263_865),
	.L (L[12974:12960]),
	.V2C_1 (V2C_865_64),
	.V2C_2 (V2C_865_85),
	.V2C_3 (V2C_865_87),
	.V2C_4 (V2C_865_110),
	.V2C_5 (V2C_865_234),
	.V2C_6 (V2C_865_263),
	.V (V_865)
);

VNU_6 #(quan_width) VNU866 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_866),
	.C2V_2 (C2V_91_866),
	.C2V_3 (C2V_93_866),
	.C2V_4 (C2V_116_866),
	.C2V_5 (C2V_240_866),
	.C2V_6 (C2V_269_866),
	.L (L[12989:12975]),
	.V2C_1 (V2C_866_70),
	.V2C_2 (V2C_866_91),
	.V2C_3 (V2C_866_93),
	.V2C_4 (V2C_866_116),
	.V2C_5 (V2C_866_240),
	.V2C_6 (V2C_866_269),
	.V (V_866)
);

VNU_6 #(quan_width) VNU867 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_867),
	.C2V_2 (C2V_97_867),
	.C2V_3 (C2V_99_867),
	.C2V_4 (C2V_122_867),
	.C2V_5 (C2V_246_867),
	.C2V_6 (C2V_275_867),
	.L (L[13004:12990]),
	.V2C_1 (V2C_867_76),
	.V2C_2 (V2C_867_97),
	.V2C_3 (V2C_867_99),
	.V2C_4 (V2C_867_122),
	.V2C_5 (V2C_867_246),
	.V2C_6 (V2C_867_275),
	.V (V_867)
);

VNU_6 #(quan_width) VNU868 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_868),
	.C2V_2 (C2V_103_868),
	.C2V_3 (C2V_105_868),
	.C2V_4 (C2V_128_868),
	.C2V_5 (C2V_252_868),
	.C2V_6 (C2V_281_868),
	.L (L[13019:13005]),
	.V2C_1 (V2C_868_82),
	.V2C_2 (V2C_868_103),
	.V2C_3 (V2C_868_105),
	.V2C_4 (V2C_868_128),
	.V2C_5 (V2C_868_252),
	.V2C_6 (V2C_868_281),
	.V (V_868)
);

VNU_6 #(quan_width) VNU869 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_869),
	.C2V_2 (C2V_109_869),
	.C2V_3 (C2V_111_869),
	.C2V_4 (C2V_134_869),
	.C2V_5 (C2V_258_869),
	.C2V_6 (C2V_287_869),
	.L (L[13034:13020]),
	.V2C_1 (V2C_869_88),
	.V2C_2 (V2C_869_109),
	.V2C_3 (V2C_869_111),
	.V2C_4 (V2C_869_134),
	.V2C_5 (V2C_869_258),
	.V2C_6 (V2C_869_287),
	.V (V_869)
);

VNU_6 #(quan_width) VNU870 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_870),
	.C2V_2 (C2V_94_870),
	.C2V_3 (C2V_115_870),
	.C2V_4 (C2V_117_870),
	.C2V_5 (C2V_140_870),
	.C2V_6 (C2V_264_870),
	.L (L[13049:13035]),
	.V2C_1 (V2C_870_5),
	.V2C_2 (V2C_870_94),
	.V2C_3 (V2C_870_115),
	.V2C_4 (V2C_870_117),
	.V2C_5 (V2C_870_140),
	.V2C_6 (V2C_870_264),
	.V (V_870)
);

VNU_6 #(quan_width) VNU871 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_871),
	.C2V_2 (C2V_100_871),
	.C2V_3 (C2V_121_871),
	.C2V_4 (C2V_123_871),
	.C2V_5 (C2V_146_871),
	.C2V_6 (C2V_270_871),
	.L (L[13064:13050]),
	.V2C_1 (V2C_871_11),
	.V2C_2 (V2C_871_100),
	.V2C_3 (V2C_871_121),
	.V2C_4 (V2C_871_123),
	.V2C_5 (V2C_871_146),
	.V2C_6 (V2C_871_270),
	.V (V_871)
);

VNU_6 #(quan_width) VNU872 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_872),
	.C2V_2 (C2V_106_872),
	.C2V_3 (C2V_127_872),
	.C2V_4 (C2V_129_872),
	.C2V_5 (C2V_152_872),
	.C2V_6 (C2V_276_872),
	.L (L[13079:13065]),
	.V2C_1 (V2C_872_17),
	.V2C_2 (V2C_872_106),
	.V2C_3 (V2C_872_127),
	.V2C_4 (V2C_872_129),
	.V2C_5 (V2C_872_152),
	.V2C_6 (V2C_872_276),
	.V (V_872)
);

VNU_6 #(quan_width) VNU873 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_873),
	.C2V_2 (C2V_112_873),
	.C2V_3 (C2V_133_873),
	.C2V_4 (C2V_135_873),
	.C2V_5 (C2V_158_873),
	.C2V_6 (C2V_282_873),
	.L (L[13094:13080]),
	.V2C_1 (V2C_873_23),
	.V2C_2 (V2C_873_112),
	.V2C_3 (V2C_873_133),
	.V2C_4 (V2C_873_135),
	.V2C_5 (V2C_873_158),
	.V2C_6 (V2C_873_282),
	.V (V_873)
);

VNU_6 #(quan_width) VNU874 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_874),
	.C2V_2 (C2V_118_874),
	.C2V_3 (C2V_139_874),
	.C2V_4 (C2V_141_874),
	.C2V_5 (C2V_164_874),
	.C2V_6 (C2V_288_874),
	.L (L[13109:13095]),
	.V2C_1 (V2C_874_29),
	.V2C_2 (V2C_874_118),
	.V2C_3 (V2C_874_139),
	.V2C_4 (V2C_874_141),
	.V2C_5 (V2C_874_164),
	.V2C_6 (V2C_874_288),
	.V (V_874)
);

VNU_6 #(quan_width) VNU875 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_875),
	.C2V_2 (C2V_35_875),
	.C2V_3 (C2V_124_875),
	.C2V_4 (C2V_145_875),
	.C2V_5 (C2V_147_875),
	.C2V_6 (C2V_170_875),
	.L (L[13124:13110]),
	.V2C_1 (V2C_875_6),
	.V2C_2 (V2C_875_35),
	.V2C_3 (V2C_875_124),
	.V2C_4 (V2C_875_145),
	.V2C_5 (V2C_875_147),
	.V2C_6 (V2C_875_170),
	.V (V_875)
);

VNU_6 #(quan_width) VNU876 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_876),
	.C2V_2 (C2V_41_876),
	.C2V_3 (C2V_130_876),
	.C2V_4 (C2V_151_876),
	.C2V_5 (C2V_153_876),
	.C2V_6 (C2V_176_876),
	.L (L[13139:13125]),
	.V2C_1 (V2C_876_12),
	.V2C_2 (V2C_876_41),
	.V2C_3 (V2C_876_130),
	.V2C_4 (V2C_876_151),
	.V2C_5 (V2C_876_153),
	.V2C_6 (V2C_876_176),
	.V (V_876)
);

VNU_6 #(quan_width) VNU877 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_877),
	.C2V_2 (C2V_47_877),
	.C2V_3 (C2V_136_877),
	.C2V_4 (C2V_157_877),
	.C2V_5 (C2V_159_877),
	.C2V_6 (C2V_182_877),
	.L (L[13154:13140]),
	.V2C_1 (V2C_877_18),
	.V2C_2 (V2C_877_47),
	.V2C_3 (V2C_877_136),
	.V2C_4 (V2C_877_157),
	.V2C_5 (V2C_877_159),
	.V2C_6 (V2C_877_182),
	.V (V_877)
);

VNU_6 #(quan_width) VNU878 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_878),
	.C2V_2 (C2V_53_878),
	.C2V_3 (C2V_142_878),
	.C2V_4 (C2V_163_878),
	.C2V_5 (C2V_165_878),
	.C2V_6 (C2V_188_878),
	.L (L[13169:13155]),
	.V2C_1 (V2C_878_24),
	.V2C_2 (V2C_878_53),
	.V2C_3 (V2C_878_142),
	.V2C_4 (V2C_878_163),
	.V2C_5 (V2C_878_165),
	.V2C_6 (V2C_878_188),
	.V (V_878)
);

VNU_6 #(quan_width) VNU879 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_879),
	.C2V_2 (C2V_59_879),
	.C2V_3 (C2V_148_879),
	.C2V_4 (C2V_169_879),
	.C2V_5 (C2V_171_879),
	.C2V_6 (C2V_194_879),
	.L (L[13184:13170]),
	.V2C_1 (V2C_879_30),
	.V2C_2 (V2C_879_59),
	.V2C_3 (V2C_879_148),
	.V2C_4 (V2C_879_169),
	.V2C_5 (V2C_879_171),
	.V2C_6 (V2C_879_194),
	.V (V_879)
);

VNU_6 #(quan_width) VNU880 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_880),
	.C2V_2 (C2V_65_880),
	.C2V_3 (C2V_154_880),
	.C2V_4 (C2V_175_880),
	.C2V_5 (C2V_177_880),
	.C2V_6 (C2V_200_880),
	.L (L[13199:13185]),
	.V2C_1 (V2C_880_36),
	.V2C_2 (V2C_880_65),
	.V2C_3 (V2C_880_154),
	.V2C_4 (V2C_880_175),
	.V2C_5 (V2C_880_177),
	.V2C_6 (V2C_880_200),
	.V (V_880)
);

VNU_6 #(quan_width) VNU881 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_881),
	.C2V_2 (C2V_71_881),
	.C2V_3 (C2V_160_881),
	.C2V_4 (C2V_181_881),
	.C2V_5 (C2V_183_881),
	.C2V_6 (C2V_206_881),
	.L (L[13214:13200]),
	.V2C_1 (V2C_881_42),
	.V2C_2 (V2C_881_71),
	.V2C_3 (V2C_881_160),
	.V2C_4 (V2C_881_181),
	.V2C_5 (V2C_881_183),
	.V2C_6 (V2C_881_206),
	.V (V_881)
);

VNU_6 #(quan_width) VNU882 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_882),
	.C2V_2 (C2V_77_882),
	.C2V_3 (C2V_166_882),
	.C2V_4 (C2V_187_882),
	.C2V_5 (C2V_189_882),
	.C2V_6 (C2V_212_882),
	.L (L[13229:13215]),
	.V2C_1 (V2C_882_48),
	.V2C_2 (V2C_882_77),
	.V2C_3 (V2C_882_166),
	.V2C_4 (V2C_882_187),
	.V2C_5 (V2C_882_189),
	.V2C_6 (V2C_882_212),
	.V (V_882)
);

VNU_6 #(quan_width) VNU883 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_54_883),
	.C2V_2 (C2V_83_883),
	.C2V_3 (C2V_172_883),
	.C2V_4 (C2V_193_883),
	.C2V_5 (C2V_195_883),
	.C2V_6 (C2V_218_883),
	.L (L[13244:13230]),
	.V2C_1 (V2C_883_54),
	.V2C_2 (V2C_883_83),
	.V2C_3 (V2C_883_172),
	.V2C_4 (V2C_883_193),
	.V2C_5 (V2C_883_195),
	.V2C_6 (V2C_883_218),
	.V (V_883)
);

VNU_6 #(quan_width) VNU884 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_60_884),
	.C2V_2 (C2V_89_884),
	.C2V_3 (C2V_178_884),
	.C2V_4 (C2V_199_884),
	.C2V_5 (C2V_201_884),
	.C2V_6 (C2V_224_884),
	.L (L[13259:13245]),
	.V2C_1 (V2C_884_60),
	.V2C_2 (V2C_884_89),
	.V2C_3 (V2C_884_178),
	.V2C_4 (V2C_884_199),
	.V2C_5 (V2C_884_201),
	.V2C_6 (V2C_884_224),
	.V (V_884)
);

VNU_6 #(quan_width) VNU885 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_66_885),
	.C2V_2 (C2V_95_885),
	.C2V_3 (C2V_184_885),
	.C2V_4 (C2V_205_885),
	.C2V_5 (C2V_207_885),
	.C2V_6 (C2V_230_885),
	.L (L[13274:13260]),
	.V2C_1 (V2C_885_66),
	.V2C_2 (V2C_885_95),
	.V2C_3 (V2C_885_184),
	.V2C_4 (V2C_885_205),
	.V2C_5 (V2C_885_207),
	.V2C_6 (V2C_885_230),
	.V (V_885)
);

VNU_6 #(quan_width) VNU886 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_72_886),
	.C2V_2 (C2V_101_886),
	.C2V_3 (C2V_190_886),
	.C2V_4 (C2V_211_886),
	.C2V_5 (C2V_213_886),
	.C2V_6 (C2V_236_886),
	.L (L[13289:13275]),
	.V2C_1 (V2C_886_72),
	.V2C_2 (V2C_886_101),
	.V2C_3 (V2C_886_190),
	.V2C_4 (V2C_886_211),
	.V2C_5 (V2C_886_213),
	.V2C_6 (V2C_886_236),
	.V (V_886)
);

VNU_6 #(quan_width) VNU887 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_78_887),
	.C2V_2 (C2V_107_887),
	.C2V_3 (C2V_196_887),
	.C2V_4 (C2V_217_887),
	.C2V_5 (C2V_219_887),
	.C2V_6 (C2V_242_887),
	.L (L[13304:13290]),
	.V2C_1 (V2C_887_78),
	.V2C_2 (V2C_887_107),
	.V2C_3 (V2C_887_196),
	.V2C_4 (V2C_887_217),
	.V2C_5 (V2C_887_219),
	.V2C_6 (V2C_887_242),
	.V (V_887)
);

VNU_6 #(quan_width) VNU888 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_84_888),
	.C2V_2 (C2V_113_888),
	.C2V_3 (C2V_202_888),
	.C2V_4 (C2V_223_888),
	.C2V_5 (C2V_225_888),
	.C2V_6 (C2V_248_888),
	.L (L[13319:13305]),
	.V2C_1 (V2C_888_84),
	.V2C_2 (V2C_888_113),
	.V2C_3 (V2C_888_202),
	.V2C_4 (V2C_888_223),
	.V2C_5 (V2C_888_225),
	.V2C_6 (V2C_888_248),
	.V (V_888)
);

VNU_6 #(quan_width) VNU889 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_90_889),
	.C2V_2 (C2V_119_889),
	.C2V_3 (C2V_208_889),
	.C2V_4 (C2V_229_889),
	.C2V_5 (C2V_231_889),
	.C2V_6 (C2V_254_889),
	.L (L[13334:13320]),
	.V2C_1 (V2C_889_90),
	.V2C_2 (V2C_889_119),
	.V2C_3 (V2C_889_208),
	.V2C_4 (V2C_889_229),
	.V2C_5 (V2C_889_231),
	.V2C_6 (V2C_889_254),
	.V (V_889)
);

VNU_6 #(quan_width) VNU890 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_96_890),
	.C2V_2 (C2V_125_890),
	.C2V_3 (C2V_214_890),
	.C2V_4 (C2V_235_890),
	.C2V_5 (C2V_237_890),
	.C2V_6 (C2V_260_890),
	.L (L[13349:13335]),
	.V2C_1 (V2C_890_96),
	.V2C_2 (V2C_890_125),
	.V2C_3 (V2C_890_214),
	.V2C_4 (V2C_890_235),
	.V2C_5 (V2C_890_237),
	.V2C_6 (V2C_890_260),
	.V (V_890)
);

VNU_6 #(quan_width) VNU891 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_102_891),
	.C2V_2 (C2V_131_891),
	.C2V_3 (C2V_220_891),
	.C2V_4 (C2V_241_891),
	.C2V_5 (C2V_243_891),
	.C2V_6 (C2V_266_891),
	.L (L[13364:13350]),
	.V2C_1 (V2C_891_102),
	.V2C_2 (V2C_891_131),
	.V2C_3 (V2C_891_220),
	.V2C_4 (V2C_891_241),
	.V2C_5 (V2C_891_243),
	.V2C_6 (V2C_891_266),
	.V (V_891)
);

VNU_6 #(quan_width) VNU892 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_108_892),
	.C2V_2 (C2V_137_892),
	.C2V_3 (C2V_226_892),
	.C2V_4 (C2V_247_892),
	.C2V_5 (C2V_249_892),
	.C2V_6 (C2V_272_892),
	.L (L[13379:13365]),
	.V2C_1 (V2C_892_108),
	.V2C_2 (V2C_892_137),
	.V2C_3 (V2C_892_226),
	.V2C_4 (V2C_892_247),
	.V2C_5 (V2C_892_249),
	.V2C_6 (V2C_892_272),
	.V (V_892)
);

VNU_6 #(quan_width) VNU893 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_114_893),
	.C2V_2 (C2V_143_893),
	.C2V_3 (C2V_232_893),
	.C2V_4 (C2V_253_893),
	.C2V_5 (C2V_255_893),
	.C2V_6 (C2V_278_893),
	.L (L[13394:13380]),
	.V2C_1 (V2C_893_114),
	.V2C_2 (V2C_893_143),
	.V2C_3 (V2C_893_232),
	.V2C_4 (V2C_893_253),
	.V2C_5 (V2C_893_255),
	.V2C_6 (V2C_893_278),
	.V (V_893)
);

VNU_6 #(quan_width) VNU894 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_120_894),
	.C2V_2 (C2V_149_894),
	.C2V_3 (C2V_238_894),
	.C2V_4 (C2V_259_894),
	.C2V_5 (C2V_261_894),
	.C2V_6 (C2V_284_894),
	.L (L[13409:13395]),
	.V2C_1 (V2C_894_120),
	.V2C_2 (V2C_894_149),
	.V2C_3 (V2C_894_238),
	.V2C_4 (V2C_894_259),
	.V2C_5 (V2C_894_261),
	.V2C_6 (V2C_894_284),
	.V (V_894)
);

VNU_6 #(quan_width) VNU895 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_895),
	.C2V_2 (C2V_126_895),
	.C2V_3 (C2V_155_895),
	.C2V_4 (C2V_244_895),
	.C2V_5 (C2V_265_895),
	.C2V_6 (C2V_267_895),
	.L (L[13424:13410]),
	.V2C_1 (V2C_895_2),
	.V2C_2 (V2C_895_126),
	.V2C_3 (V2C_895_155),
	.V2C_4 (V2C_895_244),
	.V2C_5 (V2C_895_265),
	.V2C_6 (V2C_895_267),
	.V (V_895)
);

VNU_6 #(quan_width) VNU896 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_896),
	.C2V_2 (C2V_132_896),
	.C2V_3 (C2V_161_896),
	.C2V_4 (C2V_250_896),
	.C2V_5 (C2V_271_896),
	.C2V_6 (C2V_273_896),
	.L (L[13439:13425]),
	.V2C_1 (V2C_896_8),
	.V2C_2 (V2C_896_132),
	.V2C_3 (V2C_896_161),
	.V2C_4 (V2C_896_250),
	.V2C_5 (V2C_896_271),
	.V2C_6 (V2C_896_273),
	.V (V_896)
);

VNU_6 #(quan_width) VNU897 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_897),
	.C2V_2 (C2V_138_897),
	.C2V_3 (C2V_167_897),
	.C2V_4 (C2V_256_897),
	.C2V_5 (C2V_277_897),
	.C2V_6 (C2V_279_897),
	.L (L[13454:13440]),
	.V2C_1 (V2C_897_14),
	.V2C_2 (V2C_897_138),
	.V2C_3 (V2C_897_167),
	.V2C_4 (V2C_897_256),
	.V2C_5 (V2C_897_277),
	.V2C_6 (V2C_897_279),
	.V (V_897)
);

VNU_6 #(quan_width) VNU898 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_898),
	.C2V_2 (C2V_144_898),
	.C2V_3 (C2V_173_898),
	.C2V_4 (C2V_262_898),
	.C2V_5 (C2V_283_898),
	.C2V_6 (C2V_285_898),
	.L (L[13469:13455]),
	.V2C_1 (V2C_898_20),
	.V2C_2 (V2C_898_144),
	.V2C_3 (V2C_898_173),
	.V2C_4 (V2C_898_262),
	.V2C_5 (V2C_898_283),
	.V2C_6 (V2C_898_285),
	.V (V_898)
);

VNU_6 #(quan_width) VNU899 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_899),
	.C2V_2 (C2V_3_899),
	.C2V_3 (C2V_26_899),
	.C2V_4 (C2V_150_899),
	.C2V_5 (C2V_179_899),
	.C2V_6 (C2V_268_899),
	.L (L[13484:13470]),
	.V2C_1 (V2C_899_1),
	.V2C_2 (V2C_899_3),
	.V2C_3 (V2C_899_26),
	.V2C_4 (V2C_899_150),
	.V2C_5 (V2C_899_179),
	.V2C_6 (V2C_899_268),
	.V (V_899)
);

VNU_6 #(quan_width) VNU900 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_900),
	.C2V_2 (C2V_9_900),
	.C2V_3 (C2V_32_900),
	.C2V_4 (C2V_156_900),
	.C2V_5 (C2V_185_900),
	.C2V_6 (C2V_274_900),
	.L (L[13499:13485]),
	.V2C_1 (V2C_900_7),
	.V2C_2 (V2C_900_9),
	.V2C_3 (V2C_900_32),
	.V2C_4 (V2C_900_156),
	.V2C_5 (V2C_900_185),
	.V2C_6 (V2C_900_274),
	.V (V_900)
);

VNU_6 #(quan_width) VNU901 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_901),
	.C2V_2 (C2V_15_901),
	.C2V_3 (C2V_38_901),
	.C2V_4 (C2V_162_901),
	.C2V_5 (C2V_191_901),
	.C2V_6 (C2V_280_901),
	.L (L[13514:13500]),
	.V2C_1 (V2C_901_13),
	.V2C_2 (V2C_901_15),
	.V2C_3 (V2C_901_38),
	.V2C_4 (V2C_901_162),
	.V2C_5 (V2C_901_191),
	.V2C_6 (V2C_901_280),
	.V (V_901)
);

VNU_6 #(quan_width) VNU902 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_902),
	.C2V_2 (C2V_21_902),
	.C2V_3 (C2V_44_902),
	.C2V_4 (C2V_168_902),
	.C2V_5 (C2V_197_902),
	.C2V_6 (C2V_286_902),
	.L (L[13529:13515]),
	.V2C_1 (V2C_902_19),
	.V2C_2 (V2C_902_21),
	.V2C_3 (V2C_902_44),
	.V2C_4 (V2C_902_168),
	.V2C_5 (V2C_902_197),
	.V2C_6 (V2C_902_286),
	.V (V_902)
);

VNU_6 #(quan_width) VNU903 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_903),
	.C2V_2 (C2V_25_903),
	.C2V_3 (C2V_27_903),
	.C2V_4 (C2V_50_903),
	.C2V_5 (C2V_174_903),
	.C2V_6 (C2V_203_903),
	.L (L[13544:13530]),
	.V2C_1 (V2C_903_4),
	.V2C_2 (V2C_903_25),
	.V2C_3 (V2C_903_27),
	.V2C_4 (V2C_903_50),
	.V2C_5 (V2C_903_174),
	.V2C_6 (V2C_903_203),
	.V (V_903)
);

VNU_6 #(quan_width) VNU904 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_904),
	.C2V_2 (C2V_31_904),
	.C2V_3 (C2V_33_904),
	.C2V_4 (C2V_56_904),
	.C2V_5 (C2V_180_904),
	.C2V_6 (C2V_209_904),
	.L (L[13559:13545]),
	.V2C_1 (V2C_904_10),
	.V2C_2 (V2C_904_31),
	.V2C_3 (V2C_904_33),
	.V2C_4 (V2C_904_56),
	.V2C_5 (V2C_904_180),
	.V2C_6 (V2C_904_209),
	.V (V_904)
);

VNU_6 #(quan_width) VNU905 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_905),
	.C2V_2 (C2V_37_905),
	.C2V_3 (C2V_39_905),
	.C2V_4 (C2V_62_905),
	.C2V_5 (C2V_186_905),
	.C2V_6 (C2V_215_905),
	.L (L[13574:13560]),
	.V2C_1 (V2C_905_16),
	.V2C_2 (V2C_905_37),
	.V2C_3 (V2C_905_39),
	.V2C_4 (V2C_905_62),
	.V2C_5 (V2C_905_186),
	.V2C_6 (V2C_905_215),
	.V (V_905)
);

VNU_6 #(quan_width) VNU906 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_906),
	.C2V_2 (C2V_43_906),
	.C2V_3 (C2V_45_906),
	.C2V_4 (C2V_68_906),
	.C2V_5 (C2V_192_906),
	.C2V_6 (C2V_221_906),
	.L (L[13589:13575]),
	.V2C_1 (V2C_906_22),
	.V2C_2 (V2C_906_43),
	.V2C_3 (V2C_906_45),
	.V2C_4 (V2C_906_68),
	.V2C_5 (V2C_906_192),
	.V2C_6 (V2C_906_221),
	.V (V_906)
);

VNU_6 #(quan_width) VNU907 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_907),
	.C2V_2 (C2V_49_907),
	.C2V_3 (C2V_51_907),
	.C2V_4 (C2V_74_907),
	.C2V_5 (C2V_198_907),
	.C2V_6 (C2V_227_907),
	.L (L[13604:13590]),
	.V2C_1 (V2C_907_28),
	.V2C_2 (V2C_907_49),
	.V2C_3 (V2C_907_51),
	.V2C_4 (V2C_907_74),
	.V2C_5 (V2C_907_198),
	.V2C_6 (V2C_907_227),
	.V (V_907)
);

VNU_6 #(quan_width) VNU908 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_908),
	.C2V_2 (C2V_55_908),
	.C2V_3 (C2V_57_908),
	.C2V_4 (C2V_80_908),
	.C2V_5 (C2V_204_908),
	.C2V_6 (C2V_233_908),
	.L (L[13619:13605]),
	.V2C_1 (V2C_908_34),
	.V2C_2 (V2C_908_55),
	.V2C_3 (V2C_908_57),
	.V2C_4 (V2C_908_80),
	.V2C_5 (V2C_908_204),
	.V2C_6 (V2C_908_233),
	.V (V_908)
);

VNU_6 #(quan_width) VNU909 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_909),
	.C2V_2 (C2V_61_909),
	.C2V_3 (C2V_63_909),
	.C2V_4 (C2V_86_909),
	.C2V_5 (C2V_210_909),
	.C2V_6 (C2V_239_909),
	.L (L[13634:13620]),
	.V2C_1 (V2C_909_40),
	.V2C_2 (V2C_909_61),
	.V2C_3 (V2C_909_63),
	.V2C_4 (V2C_909_86),
	.V2C_5 (V2C_909_210),
	.V2C_6 (V2C_909_239),
	.V (V_909)
);

VNU_6 #(quan_width) VNU910 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_910),
	.C2V_2 (C2V_67_910),
	.C2V_3 (C2V_69_910),
	.C2V_4 (C2V_92_910),
	.C2V_5 (C2V_216_910),
	.C2V_6 (C2V_245_910),
	.L (L[13649:13635]),
	.V2C_1 (V2C_910_46),
	.V2C_2 (V2C_910_67),
	.V2C_3 (V2C_910_69),
	.V2C_4 (V2C_910_92),
	.V2C_5 (V2C_910_216),
	.V2C_6 (V2C_910_245),
	.V (V_910)
);

VNU_6 #(quan_width) VNU911 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_911),
	.C2V_2 (C2V_73_911),
	.C2V_3 (C2V_75_911),
	.C2V_4 (C2V_98_911),
	.C2V_5 (C2V_222_911),
	.C2V_6 (C2V_251_911),
	.L (L[13664:13650]),
	.V2C_1 (V2C_911_52),
	.V2C_2 (V2C_911_73),
	.V2C_3 (V2C_911_75),
	.V2C_4 (V2C_911_98),
	.V2C_5 (V2C_911_222),
	.V2C_6 (V2C_911_251),
	.V (V_911)
);

VNU_6 #(quan_width) VNU912 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_912),
	.C2V_2 (C2V_79_912),
	.C2V_3 (C2V_81_912),
	.C2V_4 (C2V_104_912),
	.C2V_5 (C2V_228_912),
	.C2V_6 (C2V_257_912),
	.L (L[13679:13665]),
	.V2C_1 (V2C_912_58),
	.V2C_2 (V2C_912_79),
	.V2C_3 (V2C_912_81),
	.V2C_4 (V2C_912_104),
	.V2C_5 (V2C_912_228),
	.V2C_6 (V2C_912_257),
	.V (V_912)
);

VNU_6 #(quan_width) VNU913 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_913),
	.C2V_2 (C2V_111_913),
	.C2V_3 (C2V_127_913),
	.C2V_4 (C2V_150_913),
	.C2V_5 (C2V_208_913),
	.C2V_6 (C2V_263_913),
	.L (L[13694:13680]),
	.V2C_1 (V2C_913_20),
	.V2C_2 (V2C_913_111),
	.V2C_3 (V2C_913_127),
	.V2C_4 (V2C_913_150),
	.V2C_5 (V2C_913_208),
	.V2C_6 (V2C_913_263),
	.V (V_913)
);

VNU_6 #(quan_width) VNU914 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_914),
	.C2V_2 (C2V_117_914),
	.C2V_3 (C2V_133_914),
	.C2V_4 (C2V_156_914),
	.C2V_5 (C2V_214_914),
	.C2V_6 (C2V_269_914),
	.L (L[13709:13695]),
	.V2C_1 (V2C_914_26),
	.V2C_2 (V2C_914_117),
	.V2C_3 (V2C_914_133),
	.V2C_4 (V2C_914_156),
	.V2C_5 (V2C_914_214),
	.V2C_6 (V2C_914_269),
	.V (V_914)
);

VNU_6 #(quan_width) VNU915 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_915),
	.C2V_2 (C2V_123_915),
	.C2V_3 (C2V_139_915),
	.C2V_4 (C2V_162_915),
	.C2V_5 (C2V_220_915),
	.C2V_6 (C2V_275_915),
	.L (L[13724:13710]),
	.V2C_1 (V2C_915_32),
	.V2C_2 (V2C_915_123),
	.V2C_3 (V2C_915_139),
	.V2C_4 (V2C_915_162),
	.V2C_5 (V2C_915_220),
	.V2C_6 (V2C_915_275),
	.V (V_915)
);

VNU_6 #(quan_width) VNU916 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_916),
	.C2V_2 (C2V_129_916),
	.C2V_3 (C2V_145_916),
	.C2V_4 (C2V_168_916),
	.C2V_5 (C2V_226_916),
	.C2V_6 (C2V_281_916),
	.L (L[13739:13725]),
	.V2C_1 (V2C_916_38),
	.V2C_2 (V2C_916_129),
	.V2C_3 (V2C_916_145),
	.V2C_4 (V2C_916_168),
	.V2C_5 (V2C_916_226),
	.V2C_6 (V2C_916_281),
	.V (V_916)
);

VNU_6 #(quan_width) VNU917 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_917),
	.C2V_2 (C2V_135_917),
	.C2V_3 (C2V_151_917),
	.C2V_4 (C2V_174_917),
	.C2V_5 (C2V_232_917),
	.C2V_6 (C2V_287_917),
	.L (L[13754:13740]),
	.V2C_1 (V2C_917_44),
	.V2C_2 (V2C_917_135),
	.V2C_3 (V2C_917_151),
	.V2C_4 (V2C_917_174),
	.V2C_5 (V2C_917_232),
	.V2C_6 (V2C_917_287),
	.V (V_917)
);

VNU_6 #(quan_width) VNU918 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_918),
	.C2V_2 (C2V_50_918),
	.C2V_3 (C2V_141_918),
	.C2V_4 (C2V_157_918),
	.C2V_5 (C2V_180_918),
	.C2V_6 (C2V_238_918),
	.L (L[13769:13755]),
	.V2C_1 (V2C_918_5),
	.V2C_2 (V2C_918_50),
	.V2C_3 (V2C_918_141),
	.V2C_4 (V2C_918_157),
	.V2C_5 (V2C_918_180),
	.V2C_6 (V2C_918_238),
	.V (V_918)
);

VNU_6 #(quan_width) VNU919 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_919),
	.C2V_2 (C2V_56_919),
	.C2V_3 (C2V_147_919),
	.C2V_4 (C2V_163_919),
	.C2V_5 (C2V_186_919),
	.C2V_6 (C2V_244_919),
	.L (L[13784:13770]),
	.V2C_1 (V2C_919_11),
	.V2C_2 (V2C_919_56),
	.V2C_3 (V2C_919_147),
	.V2C_4 (V2C_919_163),
	.V2C_5 (V2C_919_186),
	.V2C_6 (V2C_919_244),
	.V (V_919)
);

VNU_6 #(quan_width) VNU920 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_920),
	.C2V_2 (C2V_62_920),
	.C2V_3 (C2V_153_920),
	.C2V_4 (C2V_169_920),
	.C2V_5 (C2V_192_920),
	.C2V_6 (C2V_250_920),
	.L (L[13799:13785]),
	.V2C_1 (V2C_920_17),
	.V2C_2 (V2C_920_62),
	.V2C_3 (V2C_920_153),
	.V2C_4 (V2C_920_169),
	.V2C_5 (V2C_920_192),
	.V2C_6 (V2C_920_250),
	.V (V_920)
);

VNU_6 #(quan_width) VNU921 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_921),
	.C2V_2 (C2V_68_921),
	.C2V_3 (C2V_159_921),
	.C2V_4 (C2V_175_921),
	.C2V_5 (C2V_198_921),
	.C2V_6 (C2V_256_921),
	.L (L[13814:13800]),
	.V2C_1 (V2C_921_23),
	.V2C_2 (V2C_921_68),
	.V2C_3 (V2C_921_159),
	.V2C_4 (V2C_921_175),
	.V2C_5 (V2C_921_198),
	.V2C_6 (V2C_921_256),
	.V (V_921)
);

VNU_6 #(quan_width) VNU922 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_922),
	.C2V_2 (C2V_74_922),
	.C2V_3 (C2V_165_922),
	.C2V_4 (C2V_181_922),
	.C2V_5 (C2V_204_922),
	.C2V_6 (C2V_262_922),
	.L (L[13829:13815]),
	.V2C_1 (V2C_922_29),
	.V2C_2 (V2C_922_74),
	.V2C_3 (V2C_922_165),
	.V2C_4 (V2C_922_181),
	.V2C_5 (V2C_922_204),
	.V2C_6 (V2C_922_262),
	.V (V_922)
);

VNU_6 #(quan_width) VNU923 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_923),
	.C2V_2 (C2V_80_923),
	.C2V_3 (C2V_171_923),
	.C2V_4 (C2V_187_923),
	.C2V_5 (C2V_210_923),
	.C2V_6 (C2V_268_923),
	.L (L[13844:13830]),
	.V2C_1 (V2C_923_35),
	.V2C_2 (V2C_923_80),
	.V2C_3 (V2C_923_171),
	.V2C_4 (V2C_923_187),
	.V2C_5 (V2C_923_210),
	.V2C_6 (V2C_923_268),
	.V (V_923)
);

VNU_6 #(quan_width) VNU924 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_924),
	.C2V_2 (C2V_86_924),
	.C2V_3 (C2V_177_924),
	.C2V_4 (C2V_193_924),
	.C2V_5 (C2V_216_924),
	.C2V_6 (C2V_274_924),
	.L (L[13859:13845]),
	.V2C_1 (V2C_924_41),
	.V2C_2 (V2C_924_86),
	.V2C_3 (V2C_924_177),
	.V2C_4 (V2C_924_193),
	.V2C_5 (V2C_924_216),
	.V2C_6 (V2C_924_274),
	.V (V_924)
);

VNU_6 #(quan_width) VNU925 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_925),
	.C2V_2 (C2V_92_925),
	.C2V_3 (C2V_183_925),
	.C2V_4 (C2V_199_925),
	.C2V_5 (C2V_222_925),
	.C2V_6 (C2V_280_925),
	.L (L[13874:13860]),
	.V2C_1 (V2C_925_47),
	.V2C_2 (V2C_925_92),
	.V2C_3 (V2C_925_183),
	.V2C_4 (V2C_925_199),
	.V2C_5 (V2C_925_222),
	.V2C_6 (V2C_925_280),
	.V (V_925)
);

VNU_6 #(quan_width) VNU926 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_926),
	.C2V_2 (C2V_98_926),
	.C2V_3 (C2V_189_926),
	.C2V_4 (C2V_205_926),
	.C2V_5 (C2V_228_926),
	.C2V_6 (C2V_286_926),
	.L (L[13889:13875]),
	.V2C_1 (V2C_926_53),
	.V2C_2 (V2C_926_98),
	.V2C_3 (V2C_926_189),
	.V2C_4 (V2C_926_205),
	.V2C_5 (V2C_926_228),
	.V2C_6 (V2C_926_286),
	.V (V_926)
);

VNU_6 #(quan_width) VNU927 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_927),
	.C2V_2 (C2V_59_927),
	.C2V_3 (C2V_104_927),
	.C2V_4 (C2V_195_927),
	.C2V_5 (C2V_211_927),
	.C2V_6 (C2V_234_927),
	.L (L[13904:13890]),
	.V2C_1 (V2C_927_4),
	.V2C_2 (V2C_927_59),
	.V2C_3 (V2C_927_104),
	.V2C_4 (V2C_927_195),
	.V2C_5 (V2C_927_211),
	.V2C_6 (V2C_927_234),
	.V (V_927)
);

VNU_6 #(quan_width) VNU928 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_928),
	.C2V_2 (C2V_65_928),
	.C2V_3 (C2V_110_928),
	.C2V_4 (C2V_201_928),
	.C2V_5 (C2V_217_928),
	.C2V_6 (C2V_240_928),
	.L (L[13919:13905]),
	.V2C_1 (V2C_928_10),
	.V2C_2 (V2C_928_65),
	.V2C_3 (V2C_928_110),
	.V2C_4 (V2C_928_201),
	.V2C_5 (V2C_928_217),
	.V2C_6 (V2C_928_240),
	.V (V_928)
);

VNU_6 #(quan_width) VNU929 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_929),
	.C2V_2 (C2V_71_929),
	.C2V_3 (C2V_116_929),
	.C2V_4 (C2V_207_929),
	.C2V_5 (C2V_223_929),
	.C2V_6 (C2V_246_929),
	.L (L[13934:13920]),
	.V2C_1 (V2C_929_16),
	.V2C_2 (V2C_929_71),
	.V2C_3 (V2C_929_116),
	.V2C_4 (V2C_929_207),
	.V2C_5 (V2C_929_223),
	.V2C_6 (V2C_929_246),
	.V (V_929)
);

VNU_6 #(quan_width) VNU930 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_930),
	.C2V_2 (C2V_77_930),
	.C2V_3 (C2V_122_930),
	.C2V_4 (C2V_213_930),
	.C2V_5 (C2V_229_930),
	.C2V_6 (C2V_252_930),
	.L (L[13949:13935]),
	.V2C_1 (V2C_930_22),
	.V2C_2 (V2C_930_77),
	.V2C_3 (V2C_930_122),
	.V2C_4 (V2C_930_213),
	.V2C_5 (V2C_930_229),
	.V2C_6 (V2C_930_252),
	.V (V_930)
);

VNU_6 #(quan_width) VNU931 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_931),
	.C2V_2 (C2V_83_931),
	.C2V_3 (C2V_128_931),
	.C2V_4 (C2V_219_931),
	.C2V_5 (C2V_235_931),
	.C2V_6 (C2V_258_931),
	.L (L[13964:13950]),
	.V2C_1 (V2C_931_28),
	.V2C_2 (V2C_931_83),
	.V2C_3 (V2C_931_128),
	.V2C_4 (V2C_931_219),
	.V2C_5 (V2C_931_235),
	.V2C_6 (V2C_931_258),
	.V (V_931)
);

VNU_6 #(quan_width) VNU932 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_932),
	.C2V_2 (C2V_89_932),
	.C2V_3 (C2V_134_932),
	.C2V_4 (C2V_225_932),
	.C2V_5 (C2V_241_932),
	.C2V_6 (C2V_264_932),
	.L (L[13979:13965]),
	.V2C_1 (V2C_932_34),
	.V2C_2 (V2C_932_89),
	.V2C_3 (V2C_932_134),
	.V2C_4 (V2C_932_225),
	.V2C_5 (V2C_932_241),
	.V2C_6 (V2C_932_264),
	.V (V_932)
);

VNU_6 #(quan_width) VNU933 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_933),
	.C2V_2 (C2V_95_933),
	.C2V_3 (C2V_140_933),
	.C2V_4 (C2V_231_933),
	.C2V_5 (C2V_247_933),
	.C2V_6 (C2V_270_933),
	.L (L[13994:13980]),
	.V2C_1 (V2C_933_40),
	.V2C_2 (V2C_933_95),
	.V2C_3 (V2C_933_140),
	.V2C_4 (V2C_933_231),
	.V2C_5 (V2C_933_247),
	.V2C_6 (V2C_933_270),
	.V (V_933)
);

VNU_6 #(quan_width) VNU934 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_934),
	.C2V_2 (C2V_101_934),
	.C2V_3 (C2V_146_934),
	.C2V_4 (C2V_237_934),
	.C2V_5 (C2V_253_934),
	.C2V_6 (C2V_276_934),
	.L (L[14009:13995]),
	.V2C_1 (V2C_934_46),
	.V2C_2 (V2C_934_101),
	.V2C_3 (V2C_934_146),
	.V2C_4 (V2C_934_237),
	.V2C_5 (V2C_934_253),
	.V2C_6 (V2C_934_276),
	.V (V_934)
);

VNU_6 #(quan_width) VNU935 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_935),
	.C2V_2 (C2V_107_935),
	.C2V_3 (C2V_152_935),
	.C2V_4 (C2V_243_935),
	.C2V_5 (C2V_259_935),
	.C2V_6 (C2V_282_935),
	.L (L[14024:14010]),
	.V2C_1 (V2C_935_52),
	.V2C_2 (V2C_935_107),
	.V2C_3 (V2C_935_152),
	.V2C_4 (V2C_935_243),
	.V2C_5 (V2C_935_259),
	.V2C_6 (V2C_935_282),
	.V (V_935)
);

VNU_6 #(quan_width) VNU936 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_936),
	.C2V_2 (C2V_113_936),
	.C2V_3 (C2V_158_936),
	.C2V_4 (C2V_249_936),
	.C2V_5 (C2V_265_936),
	.C2V_6 (C2V_288_936),
	.L (L[14039:14025]),
	.V2C_1 (V2C_936_58),
	.V2C_2 (V2C_936_113),
	.V2C_3 (V2C_936_158),
	.V2C_4 (V2C_936_249),
	.V2C_5 (V2C_936_265),
	.V2C_6 (V2C_936_288),
	.V (V_936)
);

VNU_6 #(quan_width) VNU937 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_937),
	.C2V_2 (C2V_64_937),
	.C2V_3 (C2V_119_937),
	.C2V_4 (C2V_164_937),
	.C2V_5 (C2V_255_937),
	.C2V_6 (C2V_271_937),
	.L (L[14054:14040]),
	.V2C_1 (V2C_937_6),
	.V2C_2 (V2C_937_64),
	.V2C_3 (V2C_937_119),
	.V2C_4 (V2C_937_164),
	.V2C_5 (V2C_937_255),
	.V2C_6 (V2C_937_271),
	.V (V_937)
);

VNU_6 #(quan_width) VNU938 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_938),
	.C2V_2 (C2V_70_938),
	.C2V_3 (C2V_125_938),
	.C2V_4 (C2V_170_938),
	.C2V_5 (C2V_261_938),
	.C2V_6 (C2V_277_938),
	.L (L[14069:14055]),
	.V2C_1 (V2C_938_12),
	.V2C_2 (V2C_938_70),
	.V2C_3 (V2C_938_125),
	.V2C_4 (V2C_938_170),
	.V2C_5 (V2C_938_261),
	.V2C_6 (V2C_938_277),
	.V (V_938)
);

VNU_6 #(quan_width) VNU939 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_939),
	.C2V_2 (C2V_76_939),
	.C2V_3 (C2V_131_939),
	.C2V_4 (C2V_176_939),
	.C2V_5 (C2V_267_939),
	.C2V_6 (C2V_283_939),
	.L (L[14084:14070]),
	.V2C_1 (V2C_939_18),
	.V2C_2 (V2C_939_76),
	.V2C_3 (V2C_939_131),
	.V2C_4 (V2C_939_176),
	.V2C_5 (V2C_939_267),
	.V2C_6 (V2C_939_283),
	.V (V_939)
);

VNU_6 #(quan_width) VNU940 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_940),
	.C2V_2 (C2V_24_940),
	.C2V_3 (C2V_82_940),
	.C2V_4 (C2V_137_940),
	.C2V_5 (C2V_182_940),
	.C2V_6 (C2V_273_940),
	.L (L[14099:14085]),
	.V2C_1 (V2C_940_1),
	.V2C_2 (V2C_940_24),
	.V2C_3 (V2C_940_82),
	.V2C_4 (V2C_940_137),
	.V2C_5 (V2C_940_182),
	.V2C_6 (V2C_940_273),
	.V (V_940)
);

VNU_6 #(quan_width) VNU941 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_941),
	.C2V_2 (C2V_30_941),
	.C2V_3 (C2V_88_941),
	.C2V_4 (C2V_143_941),
	.C2V_5 (C2V_188_941),
	.C2V_6 (C2V_279_941),
	.L (L[14114:14100]),
	.V2C_1 (V2C_941_7),
	.V2C_2 (V2C_941_30),
	.V2C_3 (V2C_941_88),
	.V2C_4 (V2C_941_143),
	.V2C_5 (V2C_941_188),
	.V2C_6 (V2C_941_279),
	.V (V_941)
);

VNU_6 #(quan_width) VNU942 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_942),
	.C2V_2 (C2V_36_942),
	.C2V_3 (C2V_94_942),
	.C2V_4 (C2V_149_942),
	.C2V_5 (C2V_194_942),
	.C2V_6 (C2V_285_942),
	.L (L[14129:14115]),
	.V2C_1 (V2C_942_13),
	.V2C_2 (V2C_942_36),
	.V2C_3 (V2C_942_94),
	.V2C_4 (V2C_942_149),
	.V2C_5 (V2C_942_194),
	.V2C_6 (V2C_942_285),
	.V (V_942)
);

VNU_6 #(quan_width) VNU943 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_943),
	.C2V_2 (C2V_19_943),
	.C2V_3 (C2V_42_943),
	.C2V_4 (C2V_100_943),
	.C2V_5 (C2V_155_943),
	.C2V_6 (C2V_200_943),
	.L (L[14144:14130]),
	.V2C_1 (V2C_943_3),
	.V2C_2 (V2C_943_19),
	.V2C_3 (V2C_943_42),
	.V2C_4 (V2C_943_100),
	.V2C_5 (V2C_943_155),
	.V2C_6 (V2C_943_200),
	.V (V_943)
);

VNU_6 #(quan_width) VNU944 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_944),
	.C2V_2 (C2V_25_944),
	.C2V_3 (C2V_48_944),
	.C2V_4 (C2V_106_944),
	.C2V_5 (C2V_161_944),
	.C2V_6 (C2V_206_944),
	.L (L[14159:14145]),
	.V2C_1 (V2C_944_9),
	.V2C_2 (V2C_944_25),
	.V2C_3 (V2C_944_48),
	.V2C_4 (V2C_944_106),
	.V2C_5 (V2C_944_161),
	.V2C_6 (V2C_944_206),
	.V (V_944)
);

VNU_6 #(quan_width) VNU945 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_945),
	.C2V_2 (C2V_31_945),
	.C2V_3 (C2V_54_945),
	.C2V_4 (C2V_112_945),
	.C2V_5 (C2V_167_945),
	.C2V_6 (C2V_212_945),
	.L (L[14174:14160]),
	.V2C_1 (V2C_945_15),
	.V2C_2 (V2C_945_31),
	.V2C_3 (V2C_945_54),
	.V2C_4 (V2C_945_112),
	.V2C_5 (V2C_945_167),
	.V2C_6 (V2C_945_212),
	.V (V_945)
);

VNU_6 #(quan_width) VNU946 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_946),
	.C2V_2 (C2V_37_946),
	.C2V_3 (C2V_60_946),
	.C2V_4 (C2V_118_946),
	.C2V_5 (C2V_173_946),
	.C2V_6 (C2V_218_946),
	.L (L[14189:14175]),
	.V2C_1 (V2C_946_21),
	.V2C_2 (V2C_946_37),
	.V2C_3 (V2C_946_60),
	.V2C_4 (V2C_946_118),
	.V2C_5 (V2C_946_173),
	.V2C_6 (V2C_946_218),
	.V (V_946)
);

VNU_6 #(quan_width) VNU947 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_947),
	.C2V_2 (C2V_43_947),
	.C2V_3 (C2V_66_947),
	.C2V_4 (C2V_124_947),
	.C2V_5 (C2V_179_947),
	.C2V_6 (C2V_224_947),
	.L (L[14204:14190]),
	.V2C_1 (V2C_947_27),
	.V2C_2 (V2C_947_43),
	.V2C_3 (V2C_947_66),
	.V2C_4 (V2C_947_124),
	.V2C_5 (V2C_947_179),
	.V2C_6 (V2C_947_224),
	.V (V_947)
);

VNU_6 #(quan_width) VNU948 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_948),
	.C2V_2 (C2V_49_948),
	.C2V_3 (C2V_72_948),
	.C2V_4 (C2V_130_948),
	.C2V_5 (C2V_185_948),
	.C2V_6 (C2V_230_948),
	.L (L[14219:14205]),
	.V2C_1 (V2C_948_33),
	.V2C_2 (V2C_948_49),
	.V2C_3 (V2C_948_72),
	.V2C_4 (V2C_948_130),
	.V2C_5 (V2C_948_185),
	.V2C_6 (V2C_948_230),
	.V (V_948)
);

VNU_6 #(quan_width) VNU949 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_949),
	.C2V_2 (C2V_55_949),
	.C2V_3 (C2V_78_949),
	.C2V_4 (C2V_136_949),
	.C2V_5 (C2V_191_949),
	.C2V_6 (C2V_236_949),
	.L (L[14234:14220]),
	.V2C_1 (V2C_949_39),
	.V2C_2 (V2C_949_55),
	.V2C_3 (V2C_949_78),
	.V2C_4 (V2C_949_136),
	.V2C_5 (V2C_949_191),
	.V2C_6 (V2C_949_236),
	.V (V_949)
);

VNU_6 #(quan_width) VNU950 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_950),
	.C2V_2 (C2V_61_950),
	.C2V_3 (C2V_84_950),
	.C2V_4 (C2V_142_950),
	.C2V_5 (C2V_197_950),
	.C2V_6 (C2V_242_950),
	.L (L[14249:14235]),
	.V2C_1 (V2C_950_45),
	.V2C_2 (V2C_950_61),
	.V2C_3 (V2C_950_84),
	.V2C_4 (V2C_950_142),
	.V2C_5 (V2C_950_197),
	.V2C_6 (V2C_950_242),
	.V (V_950)
);

VNU_6 #(quan_width) VNU951 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_951),
	.C2V_2 (C2V_67_951),
	.C2V_3 (C2V_90_951),
	.C2V_4 (C2V_148_951),
	.C2V_5 (C2V_203_951),
	.C2V_6 (C2V_248_951),
	.L (L[14264:14250]),
	.V2C_1 (V2C_951_51),
	.V2C_2 (V2C_951_67),
	.V2C_3 (V2C_951_90),
	.V2C_4 (V2C_951_148),
	.V2C_5 (V2C_951_203),
	.V2C_6 (V2C_951_248),
	.V (V_951)
);

VNU_6 #(quan_width) VNU952 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_952),
	.C2V_2 (C2V_73_952),
	.C2V_3 (C2V_96_952),
	.C2V_4 (C2V_154_952),
	.C2V_5 (C2V_209_952),
	.C2V_6 (C2V_254_952),
	.L (L[14279:14265]),
	.V2C_1 (V2C_952_57),
	.V2C_2 (V2C_952_73),
	.V2C_3 (V2C_952_96),
	.V2C_4 (V2C_952_154),
	.V2C_5 (V2C_952_209),
	.V2C_6 (V2C_952_254),
	.V (V_952)
);

VNU_6 #(quan_width) VNU953 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_953),
	.C2V_2 (C2V_79_953),
	.C2V_3 (C2V_102_953),
	.C2V_4 (C2V_160_953),
	.C2V_5 (C2V_215_953),
	.C2V_6 (C2V_260_953),
	.L (L[14294:14280]),
	.V2C_1 (V2C_953_63),
	.V2C_2 (V2C_953_79),
	.V2C_3 (V2C_953_102),
	.V2C_4 (V2C_953_160),
	.V2C_5 (V2C_953_215),
	.V2C_6 (V2C_953_260),
	.V (V_953)
);

VNU_6 #(quan_width) VNU954 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_954),
	.C2V_2 (C2V_85_954),
	.C2V_3 (C2V_108_954),
	.C2V_4 (C2V_166_954),
	.C2V_5 (C2V_221_954),
	.C2V_6 (C2V_266_954),
	.L (L[14309:14295]),
	.V2C_1 (V2C_954_69),
	.V2C_2 (V2C_954_85),
	.V2C_3 (V2C_954_108),
	.V2C_4 (V2C_954_166),
	.V2C_5 (V2C_954_221),
	.V2C_6 (V2C_954_266),
	.V (V_954)
);

VNU_6 #(quan_width) VNU955 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_955),
	.C2V_2 (C2V_91_955),
	.C2V_3 (C2V_114_955),
	.C2V_4 (C2V_172_955),
	.C2V_5 (C2V_227_955),
	.C2V_6 (C2V_272_955),
	.L (L[14324:14310]),
	.V2C_1 (V2C_955_75),
	.V2C_2 (V2C_955_91),
	.V2C_3 (V2C_955_114),
	.V2C_4 (V2C_955_172),
	.V2C_5 (V2C_955_227),
	.V2C_6 (V2C_955_272),
	.V (V_955)
);

VNU_6 #(quan_width) VNU956 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_956),
	.C2V_2 (C2V_97_956),
	.C2V_3 (C2V_120_956),
	.C2V_4 (C2V_178_956),
	.C2V_5 (C2V_233_956),
	.C2V_6 (C2V_278_956),
	.L (L[14339:14325]),
	.V2C_1 (V2C_956_81),
	.V2C_2 (V2C_956_97),
	.V2C_3 (V2C_956_120),
	.V2C_4 (V2C_956_178),
	.V2C_5 (V2C_956_233),
	.V2C_6 (V2C_956_278),
	.V (V_956)
);

VNU_6 #(quan_width) VNU957 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_957),
	.C2V_2 (C2V_103_957),
	.C2V_3 (C2V_126_957),
	.C2V_4 (C2V_184_957),
	.C2V_5 (C2V_239_957),
	.C2V_6 (C2V_284_957),
	.L (L[14354:14340]),
	.V2C_1 (V2C_957_87),
	.V2C_2 (V2C_957_103),
	.V2C_3 (V2C_957_126),
	.V2C_4 (V2C_957_184),
	.V2C_5 (V2C_957_239),
	.V2C_6 (V2C_957_284),
	.V (V_957)
);

VNU_6 #(quan_width) VNU958 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_958),
	.C2V_2 (C2V_93_958),
	.C2V_3 (C2V_109_958),
	.C2V_4 (C2V_132_958),
	.C2V_5 (C2V_190_958),
	.C2V_6 (C2V_245_958),
	.L (L[14369:14355]),
	.V2C_1 (V2C_958_2),
	.V2C_2 (V2C_958_93),
	.V2C_3 (V2C_958_109),
	.V2C_4 (V2C_958_132),
	.V2C_5 (V2C_958_190),
	.V2C_6 (V2C_958_245),
	.V (V_958)
);

VNU_6 #(quan_width) VNU959 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_959),
	.C2V_2 (C2V_99_959),
	.C2V_3 (C2V_115_959),
	.C2V_4 (C2V_138_959),
	.C2V_5 (C2V_196_959),
	.C2V_6 (C2V_251_959),
	.L (L[14384:14370]),
	.V2C_1 (V2C_959_8),
	.V2C_2 (V2C_959_99),
	.V2C_3 (V2C_959_115),
	.V2C_4 (V2C_959_138),
	.V2C_5 (V2C_959_196),
	.V2C_6 (V2C_959_251),
	.V (V_959)
);

VNU_6 #(quan_width) VNU960 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_960),
	.C2V_2 (C2V_105_960),
	.C2V_3 (C2V_121_960),
	.C2V_4 (C2V_144_960),
	.C2V_5 (C2V_202_960),
	.C2V_6 (C2V_257_960),
	.L (L[14399:14385]),
	.V2C_1 (V2C_960_14),
	.V2C_2 (V2C_960_105),
	.V2C_3 (V2C_960_121),
	.V2C_4 (V2C_960_144),
	.V2C_5 (V2C_960_202),
	.V2C_6 (V2C_960_257),
	.V (V_960)
);

VNU_6 #(quan_width) VNU961 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_961),
	.C2V_2 (C2V_122_961),
	.C2V_3 (C2V_211_961),
	.C2V_4 (C2V_228_961),
	.C2V_5 (C2V_249_961),
	.C2V_6 (C2V_280_961),
	.L (L[14414:14400]),
	.V2C_1 (V2C_961_5),
	.V2C_2 (V2C_961_122),
	.V2C_3 (V2C_961_211),
	.V2C_4 (V2C_961_228),
	.V2C_5 (V2C_961_249),
	.V2C_6 (V2C_961_280),
	.V (V_961)
);

VNU_6 #(quan_width) VNU962 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_962),
	.C2V_2 (C2V_128_962),
	.C2V_3 (C2V_217_962),
	.C2V_4 (C2V_234_962),
	.C2V_5 (C2V_255_962),
	.C2V_6 (C2V_286_962),
	.L (L[14429:14415]),
	.V2C_1 (V2C_962_11),
	.V2C_2 (V2C_962_128),
	.V2C_3 (V2C_962_217),
	.V2C_4 (V2C_962_234),
	.V2C_5 (V2C_962_255),
	.V2C_6 (V2C_962_286),
	.V (V_962)
);

VNU_6 #(quan_width) VNU963 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_963),
	.C2V_2 (C2V_17_963),
	.C2V_3 (C2V_134_963),
	.C2V_4 (C2V_223_963),
	.C2V_5 (C2V_240_963),
	.C2V_6 (C2V_261_963),
	.L (L[14444:14430]),
	.V2C_1 (V2C_963_4),
	.V2C_2 (V2C_963_17),
	.V2C_3 (V2C_963_134),
	.V2C_4 (V2C_963_223),
	.V2C_5 (V2C_963_240),
	.V2C_6 (V2C_963_261),
	.V (V_963)
);

VNU_6 #(quan_width) VNU964 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_964),
	.C2V_2 (C2V_23_964),
	.C2V_3 (C2V_140_964),
	.C2V_4 (C2V_229_964),
	.C2V_5 (C2V_246_964),
	.C2V_6 (C2V_267_964),
	.L (L[14459:14445]),
	.V2C_1 (V2C_964_10),
	.V2C_2 (V2C_964_23),
	.V2C_3 (V2C_964_140),
	.V2C_4 (V2C_964_229),
	.V2C_5 (V2C_964_246),
	.V2C_6 (V2C_964_267),
	.V (V_964)
);

VNU_6 #(quan_width) VNU965 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_965),
	.C2V_2 (C2V_29_965),
	.C2V_3 (C2V_146_965),
	.C2V_4 (C2V_235_965),
	.C2V_5 (C2V_252_965),
	.C2V_6 (C2V_273_965),
	.L (L[14474:14460]),
	.V2C_1 (V2C_965_16),
	.V2C_2 (V2C_965_29),
	.V2C_3 (V2C_965_146),
	.V2C_4 (V2C_965_235),
	.V2C_5 (V2C_965_252),
	.V2C_6 (V2C_965_273),
	.V (V_965)
);

VNU_6 #(quan_width) VNU966 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_966),
	.C2V_2 (C2V_35_966),
	.C2V_3 (C2V_152_966),
	.C2V_4 (C2V_241_966),
	.C2V_5 (C2V_258_966),
	.C2V_6 (C2V_279_966),
	.L (L[14489:14475]),
	.V2C_1 (V2C_966_22),
	.V2C_2 (V2C_966_35),
	.V2C_3 (V2C_966_152),
	.V2C_4 (V2C_966_241),
	.V2C_5 (V2C_966_258),
	.V2C_6 (V2C_966_279),
	.V (V_966)
);

VNU_6 #(quan_width) VNU967 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_967),
	.C2V_2 (C2V_41_967),
	.C2V_3 (C2V_158_967),
	.C2V_4 (C2V_247_967),
	.C2V_5 (C2V_264_967),
	.C2V_6 (C2V_285_967),
	.L (L[14504:14490]),
	.V2C_1 (V2C_967_28),
	.V2C_2 (V2C_967_41),
	.V2C_3 (V2C_967_158),
	.V2C_4 (V2C_967_247),
	.V2C_5 (V2C_967_264),
	.V2C_6 (V2C_967_285),
	.V (V_967)
);

VNU_6 #(quan_width) VNU968 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_968),
	.C2V_2 (C2V_34_968),
	.C2V_3 (C2V_47_968),
	.C2V_4 (C2V_164_968),
	.C2V_5 (C2V_253_968),
	.C2V_6 (C2V_270_968),
	.L (L[14519:14505]),
	.V2C_1 (V2C_968_3),
	.V2C_2 (V2C_968_34),
	.V2C_3 (V2C_968_47),
	.V2C_4 (V2C_968_164),
	.V2C_5 (V2C_968_253),
	.V2C_6 (V2C_968_270),
	.V (V_968)
);

VNU_6 #(quan_width) VNU969 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_969),
	.C2V_2 (C2V_40_969),
	.C2V_3 (C2V_53_969),
	.C2V_4 (C2V_170_969),
	.C2V_5 (C2V_259_969),
	.C2V_6 (C2V_276_969),
	.L (L[14534:14520]),
	.V2C_1 (V2C_969_9),
	.V2C_2 (V2C_969_40),
	.V2C_3 (V2C_969_53),
	.V2C_4 (V2C_969_170),
	.V2C_5 (V2C_969_259),
	.V2C_6 (V2C_969_276),
	.V (V_969)
);

VNU_6 #(quan_width) VNU970 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_970),
	.C2V_2 (C2V_46_970),
	.C2V_3 (C2V_59_970),
	.C2V_4 (C2V_176_970),
	.C2V_5 (C2V_265_970),
	.C2V_6 (C2V_282_970),
	.L (L[14549:14535]),
	.V2C_1 (V2C_970_15),
	.V2C_2 (V2C_970_46),
	.V2C_3 (V2C_970_59),
	.V2C_4 (V2C_970_176),
	.V2C_5 (V2C_970_265),
	.V2C_6 (V2C_970_282),
	.V (V_970)
);

VNU_6 #(quan_width) VNU971 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_971),
	.C2V_2 (C2V_52_971),
	.C2V_3 (C2V_65_971),
	.C2V_4 (C2V_182_971),
	.C2V_5 (C2V_271_971),
	.C2V_6 (C2V_288_971),
	.L (L[14564:14550]),
	.V2C_1 (V2C_971_21),
	.V2C_2 (V2C_971_52),
	.V2C_3 (V2C_971_65),
	.V2C_4 (V2C_971_182),
	.V2C_5 (V2C_971_271),
	.V2C_6 (V2C_971_288),
	.V (V_971)
);

VNU_6 #(quan_width) VNU972 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_972),
	.C2V_2 (C2V_27_972),
	.C2V_3 (C2V_58_972),
	.C2V_4 (C2V_71_972),
	.C2V_5 (C2V_188_972),
	.C2V_6 (C2V_277_972),
	.L (L[14579:14565]),
	.V2C_1 (V2C_972_6),
	.V2C_2 (V2C_972_27),
	.V2C_3 (V2C_972_58),
	.V2C_4 (V2C_972_71),
	.V2C_5 (V2C_972_188),
	.V2C_6 (V2C_972_277),
	.V (V_972)
);

VNU_6 #(quan_width) VNU973 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_973),
	.C2V_2 (C2V_33_973),
	.C2V_3 (C2V_64_973),
	.C2V_4 (C2V_77_973),
	.C2V_5 (C2V_194_973),
	.C2V_6 (C2V_283_973),
	.L (L[14594:14580]),
	.V2C_1 (V2C_973_12),
	.V2C_2 (V2C_973_33),
	.V2C_3 (V2C_973_64),
	.V2C_4 (V2C_973_77),
	.V2C_5 (V2C_973_194),
	.V2C_6 (V2C_973_283),
	.V (V_973)
);

VNU_6 #(quan_width) VNU974 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_974),
	.C2V_2 (C2V_18_974),
	.C2V_3 (C2V_39_974),
	.C2V_4 (C2V_70_974),
	.C2V_5 (C2V_83_974),
	.C2V_6 (C2V_200_974),
	.L (L[14609:14595]),
	.V2C_1 (V2C_974_1),
	.V2C_2 (V2C_974_18),
	.V2C_3 (V2C_974_39),
	.V2C_4 (V2C_974_70),
	.V2C_5 (V2C_974_83),
	.V2C_6 (V2C_974_200),
	.V (V_974)
);

VNU_6 #(quan_width) VNU975 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_975),
	.C2V_2 (C2V_24_975),
	.C2V_3 (C2V_45_975),
	.C2V_4 (C2V_76_975),
	.C2V_5 (C2V_89_975),
	.C2V_6 (C2V_206_975),
	.L (L[14624:14610]),
	.V2C_1 (V2C_975_7),
	.V2C_2 (V2C_975_24),
	.V2C_3 (V2C_975_45),
	.V2C_4 (V2C_975_76),
	.V2C_5 (V2C_975_89),
	.V2C_6 (V2C_975_206),
	.V (V_975)
);

VNU_6 #(quan_width) VNU976 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_976),
	.C2V_2 (C2V_30_976),
	.C2V_3 (C2V_51_976),
	.C2V_4 (C2V_82_976),
	.C2V_5 (C2V_95_976),
	.C2V_6 (C2V_212_976),
	.L (L[14639:14625]),
	.V2C_1 (V2C_976_13),
	.V2C_2 (V2C_976_30),
	.V2C_3 (V2C_976_51),
	.V2C_4 (V2C_976_82),
	.V2C_5 (V2C_976_95),
	.V2C_6 (V2C_976_212),
	.V (V_976)
);

VNU_6 #(quan_width) VNU977 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_977),
	.C2V_2 (C2V_36_977),
	.C2V_3 (C2V_57_977),
	.C2V_4 (C2V_88_977),
	.C2V_5 (C2V_101_977),
	.C2V_6 (C2V_218_977),
	.L (L[14654:14640]),
	.V2C_1 (V2C_977_19),
	.V2C_2 (V2C_977_36),
	.V2C_3 (V2C_977_57),
	.V2C_4 (V2C_977_88),
	.V2C_5 (V2C_977_101),
	.V2C_6 (V2C_977_218),
	.V (V_977)
);

VNU_6 #(quan_width) VNU978 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_978),
	.C2V_2 (C2V_42_978),
	.C2V_3 (C2V_63_978),
	.C2V_4 (C2V_94_978),
	.C2V_5 (C2V_107_978),
	.C2V_6 (C2V_224_978),
	.L (L[14669:14655]),
	.V2C_1 (V2C_978_25),
	.V2C_2 (V2C_978_42),
	.V2C_3 (V2C_978_63),
	.V2C_4 (V2C_978_94),
	.V2C_5 (V2C_978_107),
	.V2C_6 (V2C_978_224),
	.V (V_978)
);

VNU_6 #(quan_width) VNU979 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_979),
	.C2V_2 (C2V_48_979),
	.C2V_3 (C2V_69_979),
	.C2V_4 (C2V_100_979),
	.C2V_5 (C2V_113_979),
	.C2V_6 (C2V_230_979),
	.L (L[14684:14670]),
	.V2C_1 (V2C_979_31),
	.V2C_2 (V2C_979_48),
	.V2C_3 (V2C_979_69),
	.V2C_4 (V2C_979_100),
	.V2C_5 (V2C_979_113),
	.V2C_6 (V2C_979_230),
	.V (V_979)
);

VNU_6 #(quan_width) VNU980 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_980),
	.C2V_2 (C2V_54_980),
	.C2V_3 (C2V_75_980),
	.C2V_4 (C2V_106_980),
	.C2V_5 (C2V_119_980),
	.C2V_6 (C2V_236_980),
	.L (L[14699:14685]),
	.V2C_1 (V2C_980_37),
	.V2C_2 (V2C_980_54),
	.V2C_3 (V2C_980_75),
	.V2C_4 (V2C_980_106),
	.V2C_5 (V2C_980_119),
	.V2C_6 (V2C_980_236),
	.V (V_980)
);

VNU_6 #(quan_width) VNU981 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_981),
	.C2V_2 (C2V_60_981),
	.C2V_3 (C2V_81_981),
	.C2V_4 (C2V_112_981),
	.C2V_5 (C2V_125_981),
	.C2V_6 (C2V_242_981),
	.L (L[14714:14700]),
	.V2C_1 (V2C_981_43),
	.V2C_2 (V2C_981_60),
	.V2C_3 (V2C_981_81),
	.V2C_4 (V2C_981_112),
	.V2C_5 (V2C_981_125),
	.V2C_6 (V2C_981_242),
	.V (V_981)
);

VNU_6 #(quan_width) VNU982 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_982),
	.C2V_2 (C2V_66_982),
	.C2V_3 (C2V_87_982),
	.C2V_4 (C2V_118_982),
	.C2V_5 (C2V_131_982),
	.C2V_6 (C2V_248_982),
	.L (L[14729:14715]),
	.V2C_1 (V2C_982_49),
	.V2C_2 (V2C_982_66),
	.V2C_3 (V2C_982_87),
	.V2C_4 (V2C_982_118),
	.V2C_5 (V2C_982_131),
	.V2C_6 (V2C_982_248),
	.V (V_982)
);

VNU_6 #(quan_width) VNU983 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_983),
	.C2V_2 (C2V_72_983),
	.C2V_3 (C2V_93_983),
	.C2V_4 (C2V_124_983),
	.C2V_5 (C2V_137_983),
	.C2V_6 (C2V_254_983),
	.L (L[14744:14730]),
	.V2C_1 (V2C_983_55),
	.V2C_2 (V2C_983_72),
	.V2C_3 (V2C_983_93),
	.V2C_4 (V2C_983_124),
	.V2C_5 (V2C_983_137),
	.V2C_6 (V2C_983_254),
	.V (V_983)
);

VNU_6 #(quan_width) VNU984 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_984),
	.C2V_2 (C2V_78_984),
	.C2V_3 (C2V_99_984),
	.C2V_4 (C2V_130_984),
	.C2V_5 (C2V_143_984),
	.C2V_6 (C2V_260_984),
	.L (L[14759:14745]),
	.V2C_1 (V2C_984_61),
	.V2C_2 (V2C_984_78),
	.V2C_3 (V2C_984_99),
	.V2C_4 (V2C_984_130),
	.V2C_5 (V2C_984_143),
	.V2C_6 (V2C_984_260),
	.V (V_984)
);

VNU_6 #(quan_width) VNU985 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_985),
	.C2V_2 (C2V_84_985),
	.C2V_3 (C2V_105_985),
	.C2V_4 (C2V_136_985),
	.C2V_5 (C2V_149_985),
	.C2V_6 (C2V_266_985),
	.L (L[14774:14760]),
	.V2C_1 (V2C_985_67),
	.V2C_2 (V2C_985_84),
	.V2C_3 (V2C_985_105),
	.V2C_4 (V2C_985_136),
	.V2C_5 (V2C_985_149),
	.V2C_6 (V2C_985_266),
	.V (V_985)
);

VNU_6 #(quan_width) VNU986 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_986),
	.C2V_2 (C2V_90_986),
	.C2V_3 (C2V_111_986),
	.C2V_4 (C2V_142_986),
	.C2V_5 (C2V_155_986),
	.C2V_6 (C2V_272_986),
	.L (L[14789:14775]),
	.V2C_1 (V2C_986_73),
	.V2C_2 (V2C_986_90),
	.V2C_3 (V2C_986_111),
	.V2C_4 (V2C_986_142),
	.V2C_5 (V2C_986_155),
	.V2C_6 (V2C_986_272),
	.V (V_986)
);

VNU_6 #(quan_width) VNU987 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_987),
	.C2V_2 (C2V_96_987),
	.C2V_3 (C2V_117_987),
	.C2V_4 (C2V_148_987),
	.C2V_5 (C2V_161_987),
	.C2V_6 (C2V_278_987),
	.L (L[14804:14790]),
	.V2C_1 (V2C_987_79),
	.V2C_2 (V2C_987_96),
	.V2C_3 (V2C_987_117),
	.V2C_4 (V2C_987_148),
	.V2C_5 (V2C_987_161),
	.V2C_6 (V2C_987_278),
	.V (V_987)
);

VNU_6 #(quan_width) VNU988 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_988),
	.C2V_2 (C2V_102_988),
	.C2V_3 (C2V_123_988),
	.C2V_4 (C2V_154_988),
	.C2V_5 (C2V_167_988),
	.C2V_6 (C2V_284_988),
	.L (L[14819:14805]),
	.V2C_1 (V2C_988_85),
	.V2C_2 (V2C_988_102),
	.V2C_3 (V2C_988_123),
	.V2C_4 (V2C_988_154),
	.V2C_5 (V2C_988_167),
	.V2C_6 (V2C_988_284),
	.V (V_988)
);

VNU_6 #(quan_width) VNU989 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_989),
	.C2V_2 (C2V_91_989),
	.C2V_3 (C2V_108_989),
	.C2V_4 (C2V_129_989),
	.C2V_5 (C2V_160_989),
	.C2V_6 (C2V_173_989),
	.L (L[14834:14820]),
	.V2C_1 (V2C_989_2),
	.V2C_2 (V2C_989_91),
	.V2C_3 (V2C_989_108),
	.V2C_4 (V2C_989_129),
	.V2C_5 (V2C_989_160),
	.V2C_6 (V2C_989_173),
	.V (V_989)
);

VNU_6 #(quan_width) VNU990 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_990),
	.C2V_2 (C2V_97_990),
	.C2V_3 (C2V_114_990),
	.C2V_4 (C2V_135_990),
	.C2V_5 (C2V_166_990),
	.C2V_6 (C2V_179_990),
	.L (L[14849:14835]),
	.V2C_1 (V2C_990_8),
	.V2C_2 (V2C_990_97),
	.V2C_3 (V2C_990_114),
	.V2C_4 (V2C_990_135),
	.V2C_5 (V2C_990_166),
	.V2C_6 (V2C_990_179),
	.V (V_990)
);

VNU_6 #(quan_width) VNU991 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_991),
	.C2V_2 (C2V_103_991),
	.C2V_3 (C2V_120_991),
	.C2V_4 (C2V_141_991),
	.C2V_5 (C2V_172_991),
	.C2V_6 (C2V_185_991),
	.L (L[14864:14850]),
	.V2C_1 (V2C_991_14),
	.V2C_2 (V2C_991_103),
	.V2C_3 (V2C_991_120),
	.V2C_4 (V2C_991_141),
	.V2C_5 (V2C_991_172),
	.V2C_6 (V2C_991_185),
	.V (V_991)
);

VNU_6 #(quan_width) VNU992 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_992),
	.C2V_2 (C2V_109_992),
	.C2V_3 (C2V_126_992),
	.C2V_4 (C2V_147_992),
	.C2V_5 (C2V_178_992),
	.C2V_6 (C2V_191_992),
	.L (L[14879:14865]),
	.V2C_1 (V2C_992_20),
	.V2C_2 (V2C_992_109),
	.V2C_3 (V2C_992_126),
	.V2C_4 (V2C_992_147),
	.V2C_5 (V2C_992_178),
	.V2C_6 (V2C_992_191),
	.V (V_992)
);

VNU_6 #(quan_width) VNU993 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_993),
	.C2V_2 (C2V_115_993),
	.C2V_3 (C2V_132_993),
	.C2V_4 (C2V_153_993),
	.C2V_5 (C2V_184_993),
	.C2V_6 (C2V_197_993),
	.L (L[14894:14880]),
	.V2C_1 (V2C_993_26),
	.V2C_2 (V2C_993_115),
	.V2C_3 (V2C_993_132),
	.V2C_4 (V2C_993_153),
	.V2C_5 (V2C_993_184),
	.V2C_6 (V2C_993_197),
	.V (V_993)
);

VNU_6 #(quan_width) VNU994 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_994),
	.C2V_2 (C2V_121_994),
	.C2V_3 (C2V_138_994),
	.C2V_4 (C2V_159_994),
	.C2V_5 (C2V_190_994),
	.C2V_6 (C2V_203_994),
	.L (L[14909:14895]),
	.V2C_1 (V2C_994_32),
	.V2C_2 (V2C_994_121),
	.V2C_3 (V2C_994_138),
	.V2C_4 (V2C_994_159),
	.V2C_5 (V2C_994_190),
	.V2C_6 (V2C_994_203),
	.V (V_994)
);

VNU_6 #(quan_width) VNU995 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_995),
	.C2V_2 (C2V_127_995),
	.C2V_3 (C2V_144_995),
	.C2V_4 (C2V_165_995),
	.C2V_5 (C2V_196_995),
	.C2V_6 (C2V_209_995),
	.L (L[14924:14910]),
	.V2C_1 (V2C_995_38),
	.V2C_2 (V2C_995_127),
	.V2C_3 (V2C_995_144),
	.V2C_4 (V2C_995_165),
	.V2C_5 (V2C_995_196),
	.V2C_6 (V2C_995_209),
	.V (V_995)
);

VNU_6 #(quan_width) VNU996 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_996),
	.C2V_2 (C2V_133_996),
	.C2V_3 (C2V_150_996),
	.C2V_4 (C2V_171_996),
	.C2V_5 (C2V_202_996),
	.C2V_6 (C2V_215_996),
	.L (L[14939:14925]),
	.V2C_1 (V2C_996_44),
	.V2C_2 (V2C_996_133),
	.V2C_3 (V2C_996_150),
	.V2C_4 (V2C_996_171),
	.V2C_5 (V2C_996_202),
	.V2C_6 (V2C_996_215),
	.V (V_996)
);

VNU_6 #(quan_width) VNU997 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_997),
	.C2V_2 (C2V_139_997),
	.C2V_3 (C2V_156_997),
	.C2V_4 (C2V_177_997),
	.C2V_5 (C2V_208_997),
	.C2V_6 (C2V_221_997),
	.L (L[14954:14940]),
	.V2C_1 (V2C_997_50),
	.V2C_2 (V2C_997_139),
	.V2C_3 (V2C_997_156),
	.V2C_4 (V2C_997_177),
	.V2C_5 (V2C_997_208),
	.V2C_6 (V2C_997_221),
	.V (V_997)
);

VNU_6 #(quan_width) VNU998 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_998),
	.C2V_2 (C2V_145_998),
	.C2V_3 (C2V_162_998),
	.C2V_4 (C2V_183_998),
	.C2V_5 (C2V_214_998),
	.C2V_6 (C2V_227_998),
	.L (L[14969:14955]),
	.V2C_1 (V2C_998_56),
	.V2C_2 (V2C_998_145),
	.V2C_3 (V2C_998_162),
	.V2C_4 (V2C_998_183),
	.V2C_5 (V2C_998_214),
	.V2C_6 (V2C_998_227),
	.V (V_998)
);

VNU_6 #(quan_width) VNU999 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_999),
	.C2V_2 (C2V_151_999),
	.C2V_3 (C2V_168_999),
	.C2V_4 (C2V_189_999),
	.C2V_5 (C2V_220_999),
	.C2V_6 (C2V_233_999),
	.L (L[14984:14970]),
	.V2C_1 (V2C_999_62),
	.V2C_2 (V2C_999_151),
	.V2C_3 (V2C_999_168),
	.V2C_4 (V2C_999_189),
	.V2C_5 (V2C_999_220),
	.V2C_6 (V2C_999_233),
	.V (V_999)
);

VNU_6 #(quan_width) VNU1000 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_1000),
	.C2V_2 (C2V_157_1000),
	.C2V_3 (C2V_174_1000),
	.C2V_4 (C2V_195_1000),
	.C2V_5 (C2V_226_1000),
	.C2V_6 (C2V_239_1000),
	.L (L[14999:14985]),
	.V2C_1 (V2C_1000_68),
	.V2C_2 (V2C_1000_157),
	.V2C_3 (V2C_1000_174),
	.V2C_4 (V2C_1000_195),
	.V2C_5 (V2C_1000_226),
	.V2C_6 (V2C_1000_239),
	.V (V_1000)
);

VNU_6 #(quan_width) VNU1001 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_1001),
	.C2V_2 (C2V_163_1001),
	.C2V_3 (C2V_180_1001),
	.C2V_4 (C2V_201_1001),
	.C2V_5 (C2V_232_1001),
	.C2V_6 (C2V_245_1001),
	.L (L[15014:15000]),
	.V2C_1 (V2C_1001_74),
	.V2C_2 (V2C_1001_163),
	.V2C_3 (V2C_1001_180),
	.V2C_4 (V2C_1001_201),
	.V2C_5 (V2C_1001_232),
	.V2C_6 (V2C_1001_245),
	.V (V_1001)
);

VNU_6 #(quan_width) VNU1002 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_80_1002),
	.C2V_2 (C2V_169_1002),
	.C2V_3 (C2V_186_1002),
	.C2V_4 (C2V_207_1002),
	.C2V_5 (C2V_238_1002),
	.C2V_6 (C2V_251_1002),
	.L (L[15029:15015]),
	.V2C_1 (V2C_1002_80),
	.V2C_2 (V2C_1002_169),
	.V2C_3 (V2C_1002_186),
	.V2C_4 (V2C_1002_207),
	.V2C_5 (V2C_1002_238),
	.V2C_6 (V2C_1002_251),
	.V (V_1002)
);

VNU_6 #(quan_width) VNU1003 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_86_1003),
	.C2V_2 (C2V_175_1003),
	.C2V_3 (C2V_192_1003),
	.C2V_4 (C2V_213_1003),
	.C2V_5 (C2V_244_1003),
	.C2V_6 (C2V_257_1003),
	.L (L[15044:15030]),
	.V2C_1 (V2C_1003_86),
	.V2C_2 (V2C_1003_175),
	.V2C_3 (V2C_1003_192),
	.V2C_4 (V2C_1003_213),
	.V2C_5 (V2C_1003_244),
	.V2C_6 (V2C_1003_257),
	.V (V_1003)
);

VNU_6 #(quan_width) VNU1004 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_92_1004),
	.C2V_2 (C2V_181_1004),
	.C2V_3 (C2V_198_1004),
	.C2V_4 (C2V_219_1004),
	.C2V_5 (C2V_250_1004),
	.C2V_6 (C2V_263_1004),
	.L (L[15059:15045]),
	.V2C_1 (V2C_1004_92),
	.V2C_2 (V2C_1004_181),
	.V2C_3 (V2C_1004_198),
	.V2C_4 (V2C_1004_219),
	.V2C_5 (V2C_1004_250),
	.V2C_6 (V2C_1004_263),
	.V (V_1004)
);

VNU_6 #(quan_width) VNU1005 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_98_1005),
	.C2V_2 (C2V_187_1005),
	.C2V_3 (C2V_204_1005),
	.C2V_4 (C2V_225_1005),
	.C2V_5 (C2V_256_1005),
	.C2V_6 (C2V_269_1005),
	.L (L[15074:15060]),
	.V2C_1 (V2C_1005_98),
	.V2C_2 (V2C_1005_187),
	.V2C_3 (V2C_1005_204),
	.V2C_4 (V2C_1005_225),
	.V2C_5 (V2C_1005_256),
	.V2C_6 (V2C_1005_269),
	.V (V_1005)
);

VNU_6 #(quan_width) VNU1006 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_104_1006),
	.C2V_2 (C2V_193_1006),
	.C2V_3 (C2V_210_1006),
	.C2V_4 (C2V_231_1006),
	.C2V_5 (C2V_262_1006),
	.C2V_6 (C2V_275_1006),
	.L (L[15089:15075]),
	.V2C_1 (V2C_1006_104),
	.V2C_2 (V2C_1006_193),
	.V2C_3 (V2C_1006_210),
	.V2C_4 (V2C_1006_231),
	.V2C_5 (V2C_1006_262),
	.V2C_6 (V2C_1006_275),
	.V (V_1006)
);

VNU_6 #(quan_width) VNU1007 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_110_1007),
	.C2V_2 (C2V_199_1007),
	.C2V_3 (C2V_216_1007),
	.C2V_4 (C2V_237_1007),
	.C2V_5 (C2V_268_1007),
	.C2V_6 (C2V_281_1007),
	.L (L[15104:15090]),
	.V2C_1 (V2C_1007_110),
	.V2C_2 (V2C_1007_199),
	.V2C_3 (V2C_1007_216),
	.V2C_4 (V2C_1007_237),
	.V2C_5 (V2C_1007_268),
	.V2C_6 (V2C_1007_281),
	.V (V_1007)
);

VNU_6 #(quan_width) VNU1008 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_116_1008),
	.C2V_2 (C2V_205_1008),
	.C2V_3 (C2V_222_1008),
	.C2V_4 (C2V_243_1008),
	.C2V_5 (C2V_274_1008),
	.C2V_6 (C2V_287_1008),
	.L (L[15119:15105]),
	.V2C_1 (V2C_1008_116),
	.V2C_2 (V2C_1008_205),
	.V2C_3 (V2C_1008_222),
	.V2C_4 (V2C_1008_243),
	.V2C_5 (V2C_1008_274),
	.V2C_6 (V2C_1008_287),
	.V (V_1008)
);

VNU_6 #(quan_width) VNU1009 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_1009),
	.C2V_2 (C2V_114_1009),
	.C2V_3 (C2V_177_1009),
	.C2V_4 (C2V_218_1009),
	.C2V_5 (C2V_265_1009),
	.C2V_6 (C2V_269_1009),
	.L (L[15134:15120]),
	.V2C_1 (V2C_1009_100),
	.V2C_2 (V2C_1009_114),
	.V2C_3 (V2C_1009_177),
	.V2C_4 (V2C_1009_218),
	.V2C_5 (V2C_1009_265),
	.V2C_6 (V2C_1009_269),
	.V (V_1009)
);

VNU_6 #(quan_width) VNU1010 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_1010),
	.C2V_2 (C2V_120_1010),
	.C2V_3 (C2V_183_1010),
	.C2V_4 (C2V_224_1010),
	.C2V_5 (C2V_271_1010),
	.C2V_6 (C2V_275_1010),
	.L (L[15149:15135]),
	.V2C_1 (V2C_1010_106),
	.V2C_2 (V2C_1010_120),
	.V2C_3 (V2C_1010_183),
	.V2C_4 (V2C_1010_224),
	.V2C_5 (V2C_1010_271),
	.V2C_6 (V2C_1010_275),
	.V (V_1010)
);

VNU_6 #(quan_width) VNU1011 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_1011),
	.C2V_2 (C2V_126_1011),
	.C2V_3 (C2V_189_1011),
	.C2V_4 (C2V_230_1011),
	.C2V_5 (C2V_277_1011),
	.C2V_6 (C2V_281_1011),
	.L (L[15164:15150]),
	.V2C_1 (V2C_1011_112),
	.V2C_2 (V2C_1011_126),
	.V2C_3 (V2C_1011_189),
	.V2C_4 (V2C_1011_230),
	.V2C_5 (V2C_1011_277),
	.V2C_6 (V2C_1011_281),
	.V (V_1011)
);

VNU_6 #(quan_width) VNU1012 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_118_1012),
	.C2V_2 (C2V_132_1012),
	.C2V_3 (C2V_195_1012),
	.C2V_4 (C2V_236_1012),
	.C2V_5 (C2V_283_1012),
	.C2V_6 (C2V_287_1012),
	.L (L[15179:15165]),
	.V2C_1 (V2C_1012_118),
	.V2C_2 (V2C_1012_132),
	.V2C_3 (V2C_1012_195),
	.V2C_4 (V2C_1012_236),
	.V2C_5 (V2C_1012_283),
	.V2C_6 (V2C_1012_287),
	.V (V_1012)
);

VNU_6 #(quan_width) VNU1013 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_1013),
	.C2V_2 (C2V_5_1013),
	.C2V_3 (C2V_124_1013),
	.C2V_4 (C2V_138_1013),
	.C2V_5 (C2V_201_1013),
	.C2V_6 (C2V_242_1013),
	.L (L[15194:15180]),
	.V2C_1 (V2C_1013_1),
	.V2C_2 (V2C_1013_5),
	.V2C_3 (V2C_1013_124),
	.V2C_4 (V2C_1013_138),
	.V2C_5 (V2C_1013_201),
	.V2C_6 (V2C_1013_242),
	.V (V_1013)
);

VNU_6 #(quan_width) VNU1014 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_1014),
	.C2V_2 (C2V_11_1014),
	.C2V_3 (C2V_130_1014),
	.C2V_4 (C2V_144_1014),
	.C2V_5 (C2V_207_1014),
	.C2V_6 (C2V_248_1014),
	.L (L[15209:15195]),
	.V2C_1 (V2C_1014_7),
	.V2C_2 (V2C_1014_11),
	.V2C_3 (V2C_1014_130),
	.V2C_4 (V2C_1014_144),
	.V2C_5 (V2C_1014_207),
	.V2C_6 (V2C_1014_248),
	.V (V_1014)
);

VNU_6 #(quan_width) VNU1015 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_1015),
	.C2V_2 (C2V_17_1015),
	.C2V_3 (C2V_136_1015),
	.C2V_4 (C2V_150_1015),
	.C2V_5 (C2V_213_1015),
	.C2V_6 (C2V_254_1015),
	.L (L[15224:15210]),
	.V2C_1 (V2C_1015_13),
	.V2C_2 (V2C_1015_17),
	.V2C_3 (V2C_1015_136),
	.V2C_4 (V2C_1015_150),
	.V2C_5 (V2C_1015_213),
	.V2C_6 (V2C_1015_254),
	.V (V_1015)
);

VNU_6 #(quan_width) VNU1016 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_1016),
	.C2V_2 (C2V_23_1016),
	.C2V_3 (C2V_142_1016),
	.C2V_4 (C2V_156_1016),
	.C2V_5 (C2V_219_1016),
	.C2V_6 (C2V_260_1016),
	.L (L[15239:15225]),
	.V2C_1 (V2C_1016_19),
	.V2C_2 (V2C_1016_23),
	.V2C_3 (V2C_1016_142),
	.V2C_4 (V2C_1016_156),
	.V2C_5 (V2C_1016_219),
	.V2C_6 (V2C_1016_260),
	.V (V_1016)
);

VNU_6 #(quan_width) VNU1017 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_1017),
	.C2V_2 (C2V_29_1017),
	.C2V_3 (C2V_148_1017),
	.C2V_4 (C2V_162_1017),
	.C2V_5 (C2V_225_1017),
	.C2V_6 (C2V_266_1017),
	.L (L[15254:15240]),
	.V2C_1 (V2C_1017_25),
	.V2C_2 (V2C_1017_29),
	.V2C_3 (V2C_1017_148),
	.V2C_4 (V2C_1017_162),
	.V2C_5 (V2C_1017_225),
	.V2C_6 (V2C_1017_266),
	.V (V_1017)
);

VNU_6 #(quan_width) VNU1018 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_1018),
	.C2V_2 (C2V_35_1018),
	.C2V_3 (C2V_154_1018),
	.C2V_4 (C2V_168_1018),
	.C2V_5 (C2V_231_1018),
	.C2V_6 (C2V_272_1018),
	.L (L[15269:15255]),
	.V2C_1 (V2C_1018_31),
	.V2C_2 (V2C_1018_35),
	.V2C_3 (V2C_1018_154),
	.V2C_4 (V2C_1018_168),
	.V2C_5 (V2C_1018_231),
	.V2C_6 (V2C_1018_272),
	.V (V_1018)
);

VNU_6 #(quan_width) VNU1019 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_1019),
	.C2V_2 (C2V_41_1019),
	.C2V_3 (C2V_160_1019),
	.C2V_4 (C2V_174_1019),
	.C2V_5 (C2V_237_1019),
	.C2V_6 (C2V_278_1019),
	.L (L[15284:15270]),
	.V2C_1 (V2C_1019_37),
	.V2C_2 (V2C_1019_41),
	.V2C_3 (V2C_1019_160),
	.V2C_4 (V2C_1019_174),
	.V2C_5 (V2C_1019_237),
	.V2C_6 (V2C_1019_278),
	.V (V_1019)
);

VNU_6 #(quan_width) VNU1020 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_1020),
	.C2V_2 (C2V_47_1020),
	.C2V_3 (C2V_166_1020),
	.C2V_4 (C2V_180_1020),
	.C2V_5 (C2V_243_1020),
	.C2V_6 (C2V_284_1020),
	.L (L[15299:15285]),
	.V2C_1 (V2C_1020_43),
	.V2C_2 (V2C_1020_47),
	.V2C_3 (V2C_1020_166),
	.V2C_4 (V2C_1020_180),
	.V2C_5 (V2C_1020_243),
	.V2C_6 (V2C_1020_284),
	.V (V_1020)
);

VNU_6 #(quan_width) VNU1021 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_1021),
	.C2V_2 (C2V_49_1021),
	.C2V_3 (C2V_53_1021),
	.C2V_4 (C2V_172_1021),
	.C2V_5 (C2V_186_1021),
	.C2V_6 (C2V_249_1021),
	.L (L[15314:15300]),
	.V2C_1 (V2C_1021_2),
	.V2C_2 (V2C_1021_49),
	.V2C_3 (V2C_1021_53),
	.V2C_4 (V2C_1021_172),
	.V2C_5 (V2C_1021_186),
	.V2C_6 (V2C_1021_249),
	.V (V_1021)
);

VNU_6 #(quan_width) VNU1022 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_1022),
	.C2V_2 (C2V_55_1022),
	.C2V_3 (C2V_59_1022),
	.C2V_4 (C2V_178_1022),
	.C2V_5 (C2V_192_1022),
	.C2V_6 (C2V_255_1022),
	.L (L[15329:15315]),
	.V2C_1 (V2C_1022_8),
	.V2C_2 (V2C_1022_55),
	.V2C_3 (V2C_1022_59),
	.V2C_4 (V2C_1022_178),
	.V2C_5 (V2C_1022_192),
	.V2C_6 (V2C_1022_255),
	.V (V_1022)
);

VNU_6 #(quan_width) VNU1023 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_1023),
	.C2V_2 (C2V_61_1023),
	.C2V_3 (C2V_65_1023),
	.C2V_4 (C2V_184_1023),
	.C2V_5 (C2V_198_1023),
	.C2V_6 (C2V_261_1023),
	.L (L[15344:15330]),
	.V2C_1 (V2C_1023_14),
	.V2C_2 (V2C_1023_61),
	.V2C_3 (V2C_1023_65),
	.V2C_4 (V2C_1023_184),
	.V2C_5 (V2C_1023_198),
	.V2C_6 (V2C_1023_261),
	.V (V_1023)
);

VNU_6 #(quan_width) VNU1024 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_1024),
	.C2V_2 (C2V_67_1024),
	.C2V_3 (C2V_71_1024),
	.C2V_4 (C2V_190_1024),
	.C2V_5 (C2V_204_1024),
	.C2V_6 (C2V_267_1024),
	.L (L[15359:15345]),
	.V2C_1 (V2C_1024_20),
	.V2C_2 (V2C_1024_67),
	.V2C_3 (V2C_1024_71),
	.V2C_4 (V2C_1024_190),
	.V2C_5 (V2C_1024_204),
	.V2C_6 (V2C_1024_267),
	.V (V_1024)
);

VNU_6 #(quan_width) VNU1025 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_1025),
	.C2V_2 (C2V_73_1025),
	.C2V_3 (C2V_77_1025),
	.C2V_4 (C2V_196_1025),
	.C2V_5 (C2V_210_1025),
	.C2V_6 (C2V_273_1025),
	.L (L[15374:15360]),
	.V2C_1 (V2C_1025_26),
	.V2C_2 (V2C_1025_73),
	.V2C_3 (V2C_1025_77),
	.V2C_4 (V2C_1025_196),
	.V2C_5 (V2C_1025_210),
	.V2C_6 (V2C_1025_273),
	.V (V_1025)
);

VNU_6 #(quan_width) VNU1026 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_1026),
	.C2V_2 (C2V_79_1026),
	.C2V_3 (C2V_83_1026),
	.C2V_4 (C2V_202_1026),
	.C2V_5 (C2V_216_1026),
	.C2V_6 (C2V_279_1026),
	.L (L[15389:15375]),
	.V2C_1 (V2C_1026_32),
	.V2C_2 (V2C_1026_79),
	.V2C_3 (V2C_1026_83),
	.V2C_4 (V2C_1026_202),
	.V2C_5 (V2C_1026_216),
	.V2C_6 (V2C_1026_279),
	.V (V_1026)
);

VNU_6 #(quan_width) VNU1027 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_1027),
	.C2V_2 (C2V_85_1027),
	.C2V_3 (C2V_89_1027),
	.C2V_4 (C2V_208_1027),
	.C2V_5 (C2V_222_1027),
	.C2V_6 (C2V_285_1027),
	.L (L[15404:15390]),
	.V2C_1 (V2C_1027_38),
	.V2C_2 (V2C_1027_85),
	.V2C_3 (V2C_1027_89),
	.V2C_4 (V2C_1027_208),
	.V2C_5 (V2C_1027_222),
	.V2C_6 (V2C_1027_285),
	.V (V_1027)
);

VNU_6 #(quan_width) VNU1028 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_1028),
	.C2V_2 (C2V_44_1028),
	.C2V_3 (C2V_91_1028),
	.C2V_4 (C2V_95_1028),
	.C2V_5 (C2V_214_1028),
	.C2V_6 (C2V_228_1028),
	.L (L[15419:15405]),
	.V2C_1 (V2C_1028_3),
	.V2C_2 (V2C_1028_44),
	.V2C_3 (V2C_1028_91),
	.V2C_4 (V2C_1028_95),
	.V2C_5 (V2C_1028_214),
	.V2C_6 (V2C_1028_228),
	.V (V_1028)
);

VNU_6 #(quan_width) VNU1029 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_1029),
	.C2V_2 (C2V_50_1029),
	.C2V_3 (C2V_97_1029),
	.C2V_4 (C2V_101_1029),
	.C2V_5 (C2V_220_1029),
	.C2V_6 (C2V_234_1029),
	.L (L[15434:15420]),
	.V2C_1 (V2C_1029_9),
	.V2C_2 (V2C_1029_50),
	.V2C_3 (V2C_1029_97),
	.V2C_4 (V2C_1029_101),
	.V2C_5 (V2C_1029_220),
	.V2C_6 (V2C_1029_234),
	.V (V_1029)
);

VNU_6 #(quan_width) VNU1030 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_1030),
	.C2V_2 (C2V_56_1030),
	.C2V_3 (C2V_103_1030),
	.C2V_4 (C2V_107_1030),
	.C2V_5 (C2V_226_1030),
	.C2V_6 (C2V_240_1030),
	.L (L[15449:15435]),
	.V2C_1 (V2C_1030_15),
	.V2C_2 (V2C_1030_56),
	.V2C_3 (V2C_1030_103),
	.V2C_4 (V2C_1030_107),
	.V2C_5 (V2C_1030_226),
	.V2C_6 (V2C_1030_240),
	.V (V_1030)
);

VNU_6 #(quan_width) VNU1031 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_1031),
	.C2V_2 (C2V_62_1031),
	.C2V_3 (C2V_109_1031),
	.C2V_4 (C2V_113_1031),
	.C2V_5 (C2V_232_1031),
	.C2V_6 (C2V_246_1031),
	.L (L[15464:15450]),
	.V2C_1 (V2C_1031_21),
	.V2C_2 (V2C_1031_62),
	.V2C_3 (V2C_1031_109),
	.V2C_4 (V2C_1031_113),
	.V2C_5 (V2C_1031_232),
	.V2C_6 (V2C_1031_246),
	.V (V_1031)
);

VNU_6 #(quan_width) VNU1032 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_1032),
	.C2V_2 (C2V_68_1032),
	.C2V_3 (C2V_115_1032),
	.C2V_4 (C2V_119_1032),
	.C2V_5 (C2V_238_1032),
	.C2V_6 (C2V_252_1032),
	.L (L[15479:15465]),
	.V2C_1 (V2C_1032_27),
	.V2C_2 (V2C_1032_68),
	.V2C_3 (V2C_1032_115),
	.V2C_4 (V2C_1032_119),
	.V2C_5 (V2C_1032_238),
	.V2C_6 (V2C_1032_252),
	.V (V_1032)
);

VNU_6 #(quan_width) VNU1033 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_1033),
	.C2V_2 (C2V_74_1033),
	.C2V_3 (C2V_121_1033),
	.C2V_4 (C2V_125_1033),
	.C2V_5 (C2V_244_1033),
	.C2V_6 (C2V_258_1033),
	.L (L[15494:15480]),
	.V2C_1 (V2C_1033_33),
	.V2C_2 (V2C_1033_74),
	.V2C_3 (V2C_1033_121),
	.V2C_4 (V2C_1033_125),
	.V2C_5 (V2C_1033_244),
	.V2C_6 (V2C_1033_258),
	.V (V_1033)
);

VNU_6 #(quan_width) VNU1034 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_1034),
	.C2V_2 (C2V_80_1034),
	.C2V_3 (C2V_127_1034),
	.C2V_4 (C2V_131_1034),
	.C2V_5 (C2V_250_1034),
	.C2V_6 (C2V_264_1034),
	.L (L[15509:15495]),
	.V2C_1 (V2C_1034_39),
	.V2C_2 (V2C_1034_80),
	.V2C_3 (V2C_1034_127),
	.V2C_4 (V2C_1034_131),
	.V2C_5 (V2C_1034_250),
	.V2C_6 (V2C_1034_264),
	.V (V_1034)
);

VNU_6 #(quan_width) VNU1035 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_1035),
	.C2V_2 (C2V_86_1035),
	.C2V_3 (C2V_133_1035),
	.C2V_4 (C2V_137_1035),
	.C2V_5 (C2V_256_1035),
	.C2V_6 (C2V_270_1035),
	.L (L[15524:15510]),
	.V2C_1 (V2C_1035_45),
	.V2C_2 (V2C_1035_86),
	.V2C_3 (V2C_1035_133),
	.V2C_4 (V2C_1035_137),
	.V2C_5 (V2C_1035_256),
	.V2C_6 (V2C_1035_270),
	.V (V_1035)
);

VNU_6 #(quan_width) VNU1036 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_1036),
	.C2V_2 (C2V_92_1036),
	.C2V_3 (C2V_139_1036),
	.C2V_4 (C2V_143_1036),
	.C2V_5 (C2V_262_1036),
	.C2V_6 (C2V_276_1036),
	.L (L[15539:15525]),
	.V2C_1 (V2C_1036_51),
	.V2C_2 (V2C_1036_92),
	.V2C_3 (V2C_1036_139),
	.V2C_4 (V2C_1036_143),
	.V2C_5 (V2C_1036_262),
	.V2C_6 (V2C_1036_276),
	.V (V_1036)
);

VNU_6 #(quan_width) VNU1037 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_1037),
	.C2V_2 (C2V_98_1037),
	.C2V_3 (C2V_145_1037),
	.C2V_4 (C2V_149_1037),
	.C2V_5 (C2V_268_1037),
	.C2V_6 (C2V_282_1037),
	.L (L[15554:15540]),
	.V2C_1 (V2C_1037_57),
	.V2C_2 (V2C_1037_98),
	.V2C_3 (V2C_1037_145),
	.V2C_4 (V2C_1037_149),
	.V2C_5 (V2C_1037_268),
	.V2C_6 (V2C_1037_282),
	.V (V_1037)
);

VNU_6 #(quan_width) VNU1038 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_1038),
	.C2V_2 (C2V_104_1038),
	.C2V_3 (C2V_151_1038),
	.C2V_4 (C2V_155_1038),
	.C2V_5 (C2V_274_1038),
	.C2V_6 (C2V_288_1038),
	.L (L[15569:15555]),
	.V2C_1 (V2C_1038_63),
	.V2C_2 (V2C_1038_104),
	.V2C_3 (V2C_1038_151),
	.V2C_4 (V2C_1038_155),
	.V2C_5 (V2C_1038_274),
	.V2C_6 (V2C_1038_288),
	.V (V_1038)
);

VNU_6 #(quan_width) VNU1039 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_1039),
	.C2V_2 (C2V_69_1039),
	.C2V_3 (C2V_110_1039),
	.C2V_4 (C2V_157_1039),
	.C2V_5 (C2V_161_1039),
	.C2V_6 (C2V_280_1039),
	.L (L[15584:15570]),
	.V2C_1 (V2C_1039_6),
	.V2C_2 (V2C_1039_69),
	.V2C_3 (V2C_1039_110),
	.V2C_4 (V2C_1039_157),
	.V2C_5 (V2C_1039_161),
	.V2C_6 (V2C_1039_280),
	.V (V_1039)
);

VNU_6 #(quan_width) VNU1040 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_1040),
	.C2V_2 (C2V_75_1040),
	.C2V_3 (C2V_116_1040),
	.C2V_4 (C2V_163_1040),
	.C2V_5 (C2V_167_1040),
	.C2V_6 (C2V_286_1040),
	.L (L[15599:15585]),
	.V2C_1 (V2C_1040_12),
	.V2C_2 (V2C_1040_75),
	.V2C_3 (V2C_1040_116),
	.V2C_4 (V2C_1040_163),
	.V2C_5 (V2C_1040_167),
	.V2C_6 (V2C_1040_286),
	.V (V_1040)
);

VNU_6 #(quan_width) VNU1041 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_1041),
	.C2V_2 (C2V_18_1041),
	.C2V_3 (C2V_81_1041),
	.C2V_4 (C2V_122_1041),
	.C2V_5 (C2V_169_1041),
	.C2V_6 (C2V_173_1041),
	.L (L[15614:15600]),
	.V2C_1 (V2C_1041_4),
	.V2C_2 (V2C_1041_18),
	.V2C_3 (V2C_1041_81),
	.V2C_4 (V2C_1041_122),
	.V2C_5 (V2C_1041_169),
	.V2C_6 (V2C_1041_173),
	.V (V_1041)
);

VNU_6 #(quan_width) VNU1042 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_1042),
	.C2V_2 (C2V_24_1042),
	.C2V_3 (C2V_87_1042),
	.C2V_4 (C2V_128_1042),
	.C2V_5 (C2V_175_1042),
	.C2V_6 (C2V_179_1042),
	.L (L[15629:15615]),
	.V2C_1 (V2C_1042_10),
	.V2C_2 (V2C_1042_24),
	.V2C_3 (V2C_1042_87),
	.V2C_4 (V2C_1042_128),
	.V2C_5 (V2C_1042_175),
	.V2C_6 (V2C_1042_179),
	.V (V_1042)
);

VNU_6 #(quan_width) VNU1043 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_1043),
	.C2V_2 (C2V_30_1043),
	.C2V_3 (C2V_93_1043),
	.C2V_4 (C2V_134_1043),
	.C2V_5 (C2V_181_1043),
	.C2V_6 (C2V_185_1043),
	.L (L[15644:15630]),
	.V2C_1 (V2C_1043_16),
	.V2C_2 (V2C_1043_30),
	.V2C_3 (V2C_1043_93),
	.V2C_4 (V2C_1043_134),
	.V2C_5 (V2C_1043_181),
	.V2C_6 (V2C_1043_185),
	.V (V_1043)
);

VNU_6 #(quan_width) VNU1044 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_1044),
	.C2V_2 (C2V_36_1044),
	.C2V_3 (C2V_99_1044),
	.C2V_4 (C2V_140_1044),
	.C2V_5 (C2V_187_1044),
	.C2V_6 (C2V_191_1044),
	.L (L[15659:15645]),
	.V2C_1 (V2C_1044_22),
	.V2C_2 (V2C_1044_36),
	.V2C_3 (V2C_1044_99),
	.V2C_4 (V2C_1044_140),
	.V2C_5 (V2C_1044_187),
	.V2C_6 (V2C_1044_191),
	.V (V_1044)
);

VNU_6 #(quan_width) VNU1045 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_1045),
	.C2V_2 (C2V_42_1045),
	.C2V_3 (C2V_105_1045),
	.C2V_4 (C2V_146_1045),
	.C2V_5 (C2V_193_1045),
	.C2V_6 (C2V_197_1045),
	.L (L[15674:15660]),
	.V2C_1 (V2C_1045_28),
	.V2C_2 (V2C_1045_42),
	.V2C_3 (V2C_1045_105),
	.V2C_4 (V2C_1045_146),
	.V2C_5 (V2C_1045_193),
	.V2C_6 (V2C_1045_197),
	.V (V_1045)
);

VNU_6 #(quan_width) VNU1046 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_1046),
	.C2V_2 (C2V_48_1046),
	.C2V_3 (C2V_111_1046),
	.C2V_4 (C2V_152_1046),
	.C2V_5 (C2V_199_1046),
	.C2V_6 (C2V_203_1046),
	.L (L[15689:15675]),
	.V2C_1 (V2C_1046_34),
	.V2C_2 (V2C_1046_48),
	.V2C_3 (V2C_1046_111),
	.V2C_4 (V2C_1046_152),
	.V2C_5 (V2C_1046_199),
	.V2C_6 (V2C_1046_203),
	.V (V_1046)
);

VNU_6 #(quan_width) VNU1047 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_1047),
	.C2V_2 (C2V_54_1047),
	.C2V_3 (C2V_117_1047),
	.C2V_4 (C2V_158_1047),
	.C2V_5 (C2V_205_1047),
	.C2V_6 (C2V_209_1047),
	.L (L[15704:15690]),
	.V2C_1 (V2C_1047_40),
	.V2C_2 (V2C_1047_54),
	.V2C_3 (V2C_1047_117),
	.V2C_4 (V2C_1047_158),
	.V2C_5 (V2C_1047_205),
	.V2C_6 (V2C_1047_209),
	.V (V_1047)
);

VNU_6 #(quan_width) VNU1048 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_1048),
	.C2V_2 (C2V_60_1048),
	.C2V_3 (C2V_123_1048),
	.C2V_4 (C2V_164_1048),
	.C2V_5 (C2V_211_1048),
	.C2V_6 (C2V_215_1048),
	.L (L[15719:15705]),
	.V2C_1 (V2C_1048_46),
	.V2C_2 (V2C_1048_60),
	.V2C_3 (V2C_1048_123),
	.V2C_4 (V2C_1048_164),
	.V2C_5 (V2C_1048_211),
	.V2C_6 (V2C_1048_215),
	.V (V_1048)
);

VNU_6 #(quan_width) VNU1049 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_1049),
	.C2V_2 (C2V_66_1049),
	.C2V_3 (C2V_129_1049),
	.C2V_4 (C2V_170_1049),
	.C2V_5 (C2V_217_1049),
	.C2V_6 (C2V_221_1049),
	.L (L[15734:15720]),
	.V2C_1 (V2C_1049_52),
	.V2C_2 (V2C_1049_66),
	.V2C_3 (V2C_1049_129),
	.V2C_4 (V2C_1049_170),
	.V2C_5 (V2C_1049_217),
	.V2C_6 (V2C_1049_221),
	.V (V_1049)
);

VNU_6 #(quan_width) VNU1050 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_1050),
	.C2V_2 (C2V_72_1050),
	.C2V_3 (C2V_135_1050),
	.C2V_4 (C2V_176_1050),
	.C2V_5 (C2V_223_1050),
	.C2V_6 (C2V_227_1050),
	.L (L[15749:15735]),
	.V2C_1 (V2C_1050_58),
	.V2C_2 (V2C_1050_72),
	.V2C_3 (V2C_1050_135),
	.V2C_4 (V2C_1050_176),
	.V2C_5 (V2C_1050_223),
	.V2C_6 (V2C_1050_227),
	.V (V_1050)
);

VNU_6 #(quan_width) VNU1051 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_1051),
	.C2V_2 (C2V_78_1051),
	.C2V_3 (C2V_141_1051),
	.C2V_4 (C2V_182_1051),
	.C2V_5 (C2V_229_1051),
	.C2V_6 (C2V_233_1051),
	.L (L[15764:15750]),
	.V2C_1 (V2C_1051_64),
	.V2C_2 (V2C_1051_78),
	.V2C_3 (V2C_1051_141),
	.V2C_4 (V2C_1051_182),
	.V2C_5 (V2C_1051_229),
	.V2C_6 (V2C_1051_233),
	.V (V_1051)
);

VNU_6 #(quan_width) VNU1052 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_1052),
	.C2V_2 (C2V_84_1052),
	.C2V_3 (C2V_147_1052),
	.C2V_4 (C2V_188_1052),
	.C2V_5 (C2V_235_1052),
	.C2V_6 (C2V_239_1052),
	.L (L[15779:15765]),
	.V2C_1 (V2C_1052_70),
	.V2C_2 (V2C_1052_84),
	.V2C_3 (V2C_1052_147),
	.V2C_4 (V2C_1052_188),
	.V2C_5 (V2C_1052_235),
	.V2C_6 (V2C_1052_239),
	.V (V_1052)
);

VNU_6 #(quan_width) VNU1053 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_1053),
	.C2V_2 (C2V_90_1053),
	.C2V_3 (C2V_153_1053),
	.C2V_4 (C2V_194_1053),
	.C2V_5 (C2V_241_1053),
	.C2V_6 (C2V_245_1053),
	.L (L[15794:15780]),
	.V2C_1 (V2C_1053_76),
	.V2C_2 (V2C_1053_90),
	.V2C_3 (V2C_1053_153),
	.V2C_4 (V2C_1053_194),
	.V2C_5 (V2C_1053_241),
	.V2C_6 (V2C_1053_245),
	.V (V_1053)
);

VNU_6 #(quan_width) VNU1054 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_1054),
	.C2V_2 (C2V_96_1054),
	.C2V_3 (C2V_159_1054),
	.C2V_4 (C2V_200_1054),
	.C2V_5 (C2V_247_1054),
	.C2V_6 (C2V_251_1054),
	.L (L[15809:15795]),
	.V2C_1 (V2C_1054_82),
	.V2C_2 (V2C_1054_96),
	.V2C_3 (V2C_1054_159),
	.V2C_4 (V2C_1054_200),
	.V2C_5 (V2C_1054_247),
	.V2C_6 (V2C_1054_251),
	.V (V_1054)
);

VNU_6 #(quan_width) VNU1055 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_1055),
	.C2V_2 (C2V_102_1055),
	.C2V_3 (C2V_165_1055),
	.C2V_4 (C2V_206_1055),
	.C2V_5 (C2V_253_1055),
	.C2V_6 (C2V_257_1055),
	.L (L[15824:15810]),
	.V2C_1 (V2C_1055_88),
	.V2C_2 (V2C_1055_102),
	.V2C_3 (V2C_1055_165),
	.V2C_4 (V2C_1055_206),
	.V2C_5 (V2C_1055_253),
	.V2C_6 (V2C_1055_257),
	.V (V_1055)
);

VNU_6 #(quan_width) VNU1056 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_1056),
	.C2V_2 (C2V_108_1056),
	.C2V_3 (C2V_171_1056),
	.C2V_4 (C2V_212_1056),
	.C2V_5 (C2V_259_1056),
	.C2V_6 (C2V_263_1056),
	.L (L[15839:15825]),
	.V2C_1 (V2C_1056_94),
	.V2C_2 (V2C_1056_108),
	.V2C_3 (V2C_1056_171),
	.V2C_4 (V2C_1056_212),
	.V2C_5 (V2C_1056_259),
	.V2C_6 (V2C_1056_263),
	.V (V_1056)
);

VNU_6 #(quan_width) VNU1057 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_1057),
	.C2V_2 (C2V_104_1057),
	.C2V_3 (C2V_109_1057),
	.C2V_4 (C2V_226_1057),
	.C2V_5 (C2V_263_1057),
	.C2V_6 (C2V_285_1057),
	.L (L[15854:15840]),
	.V2C_1 (V2C_1057_18),
	.V2C_2 (V2C_1057_104),
	.V2C_3 (V2C_1057_109),
	.V2C_4 (V2C_1057_226),
	.V2C_5 (V2C_1057_263),
	.V2C_6 (V2C_1057_285),
	.V (V_1057)
);

VNU_6 #(quan_width) VNU1058 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_1058),
	.C2V_2 (C2V_24_1058),
	.C2V_3 (C2V_110_1058),
	.C2V_4 (C2V_115_1058),
	.C2V_5 (C2V_232_1058),
	.C2V_6 (C2V_269_1058),
	.L (L[15869:15855]),
	.V2C_1 (V2C_1058_3),
	.V2C_2 (V2C_1058_24),
	.V2C_3 (V2C_1058_110),
	.V2C_4 (V2C_1058_115),
	.V2C_5 (V2C_1058_232),
	.V2C_6 (V2C_1058_269),
	.V (V_1058)
);

VNU_6 #(quan_width) VNU1059 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_1059),
	.C2V_2 (C2V_30_1059),
	.C2V_3 (C2V_116_1059),
	.C2V_4 (C2V_121_1059),
	.C2V_5 (C2V_238_1059),
	.C2V_6 (C2V_275_1059),
	.L (L[15884:15870]),
	.V2C_1 (V2C_1059_9),
	.V2C_2 (V2C_1059_30),
	.V2C_3 (V2C_1059_116),
	.V2C_4 (V2C_1059_121),
	.V2C_5 (V2C_1059_238),
	.V2C_6 (V2C_1059_275),
	.V (V_1059)
);

VNU_6 #(quan_width) VNU1060 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_1060),
	.C2V_2 (C2V_36_1060),
	.C2V_3 (C2V_122_1060),
	.C2V_4 (C2V_127_1060),
	.C2V_5 (C2V_244_1060),
	.C2V_6 (C2V_281_1060),
	.L (L[15899:15885]),
	.V2C_1 (V2C_1060_15),
	.V2C_2 (V2C_1060_36),
	.V2C_3 (V2C_1060_122),
	.V2C_4 (V2C_1060_127),
	.V2C_5 (V2C_1060_244),
	.V2C_6 (V2C_1060_281),
	.V (V_1060)
);

VNU_6 #(quan_width) VNU1061 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_1061),
	.C2V_2 (C2V_42_1061),
	.C2V_3 (C2V_128_1061),
	.C2V_4 (C2V_133_1061),
	.C2V_5 (C2V_250_1061),
	.C2V_6 (C2V_287_1061),
	.L (L[15914:15900]),
	.V2C_1 (V2C_1061_21),
	.V2C_2 (V2C_1061_42),
	.V2C_3 (V2C_1061_128),
	.V2C_4 (V2C_1061_133),
	.V2C_5 (V2C_1061_250),
	.V2C_6 (V2C_1061_287),
	.V (V_1061)
);

VNU_6 #(quan_width) VNU1062 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_1062),
	.C2V_2 (C2V_27_1062),
	.C2V_3 (C2V_48_1062),
	.C2V_4 (C2V_134_1062),
	.C2V_5 (C2V_139_1062),
	.C2V_6 (C2V_256_1062),
	.L (L[15929:15915]),
	.V2C_1 (V2C_1062_5),
	.V2C_2 (V2C_1062_27),
	.V2C_3 (V2C_1062_48),
	.V2C_4 (V2C_1062_134),
	.V2C_5 (V2C_1062_139),
	.V2C_6 (V2C_1062_256),
	.V (V_1062)
);

VNU_6 #(quan_width) VNU1063 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_1063),
	.C2V_2 (C2V_33_1063),
	.C2V_3 (C2V_54_1063),
	.C2V_4 (C2V_140_1063),
	.C2V_5 (C2V_145_1063),
	.C2V_6 (C2V_262_1063),
	.L (L[15944:15930]),
	.V2C_1 (V2C_1063_11),
	.V2C_2 (V2C_1063_33),
	.V2C_3 (V2C_1063_54),
	.V2C_4 (V2C_1063_140),
	.V2C_5 (V2C_1063_145),
	.V2C_6 (V2C_1063_262),
	.V (V_1063)
);

VNU_6 #(quan_width) VNU1064 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_1064),
	.C2V_2 (C2V_39_1064),
	.C2V_3 (C2V_60_1064),
	.C2V_4 (C2V_146_1064),
	.C2V_5 (C2V_151_1064),
	.C2V_6 (C2V_268_1064),
	.L (L[15959:15945]),
	.V2C_1 (V2C_1064_17),
	.V2C_2 (V2C_1064_39),
	.V2C_3 (V2C_1064_60),
	.V2C_4 (V2C_1064_146),
	.V2C_5 (V2C_1064_151),
	.V2C_6 (V2C_1064_268),
	.V (V_1064)
);

VNU_6 #(quan_width) VNU1065 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_1065),
	.C2V_2 (C2V_45_1065),
	.C2V_3 (C2V_66_1065),
	.C2V_4 (C2V_152_1065),
	.C2V_5 (C2V_157_1065),
	.C2V_6 (C2V_274_1065),
	.L (L[15974:15960]),
	.V2C_1 (V2C_1065_23),
	.V2C_2 (V2C_1065_45),
	.V2C_3 (V2C_1065_66),
	.V2C_4 (V2C_1065_152),
	.V2C_5 (V2C_1065_157),
	.V2C_6 (V2C_1065_274),
	.V (V_1065)
);

VNU_6 #(quan_width) VNU1066 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_1066),
	.C2V_2 (C2V_51_1066),
	.C2V_3 (C2V_72_1066),
	.C2V_4 (C2V_158_1066),
	.C2V_5 (C2V_163_1066),
	.C2V_6 (C2V_280_1066),
	.L (L[15989:15975]),
	.V2C_1 (V2C_1066_29),
	.V2C_2 (V2C_1066_51),
	.V2C_3 (V2C_1066_72),
	.V2C_4 (V2C_1066_158),
	.V2C_5 (V2C_1066_163),
	.V2C_6 (V2C_1066_280),
	.V (V_1066)
);

VNU_6 #(quan_width) VNU1067 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_1067),
	.C2V_2 (C2V_57_1067),
	.C2V_3 (C2V_78_1067),
	.C2V_4 (C2V_164_1067),
	.C2V_5 (C2V_169_1067),
	.C2V_6 (C2V_286_1067),
	.L (L[16004:15990]),
	.V2C_1 (V2C_1067_35),
	.V2C_2 (V2C_1067_57),
	.V2C_3 (V2C_1067_78),
	.V2C_4 (V2C_1067_164),
	.V2C_5 (V2C_1067_169),
	.V2C_6 (V2C_1067_286),
	.V (V_1067)
);

VNU_6 #(quan_width) VNU1068 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_1068),
	.C2V_2 (C2V_41_1068),
	.C2V_3 (C2V_63_1068),
	.C2V_4 (C2V_84_1068),
	.C2V_5 (C2V_170_1068),
	.C2V_6 (C2V_175_1068),
	.L (L[16019:16005]),
	.V2C_1 (V2C_1068_4),
	.V2C_2 (V2C_1068_41),
	.V2C_3 (V2C_1068_63),
	.V2C_4 (V2C_1068_84),
	.V2C_5 (V2C_1068_170),
	.V2C_6 (V2C_1068_175),
	.V (V_1068)
);

VNU_6 #(quan_width) VNU1069 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_1069),
	.C2V_2 (C2V_47_1069),
	.C2V_3 (C2V_69_1069),
	.C2V_4 (C2V_90_1069),
	.C2V_5 (C2V_176_1069),
	.C2V_6 (C2V_181_1069),
	.L (L[16034:16020]),
	.V2C_1 (V2C_1069_10),
	.V2C_2 (V2C_1069_47),
	.V2C_3 (V2C_1069_69),
	.V2C_4 (V2C_1069_90),
	.V2C_5 (V2C_1069_176),
	.V2C_6 (V2C_1069_181),
	.V (V_1069)
);

VNU_6 #(quan_width) VNU1070 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_1070),
	.C2V_2 (C2V_53_1070),
	.C2V_3 (C2V_75_1070),
	.C2V_4 (C2V_96_1070),
	.C2V_5 (C2V_182_1070),
	.C2V_6 (C2V_187_1070),
	.L (L[16049:16035]),
	.V2C_1 (V2C_1070_16),
	.V2C_2 (V2C_1070_53),
	.V2C_3 (V2C_1070_75),
	.V2C_4 (V2C_1070_96),
	.V2C_5 (V2C_1070_182),
	.V2C_6 (V2C_1070_187),
	.V (V_1070)
);

VNU_6 #(quan_width) VNU1071 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_1071),
	.C2V_2 (C2V_59_1071),
	.C2V_3 (C2V_81_1071),
	.C2V_4 (C2V_102_1071),
	.C2V_5 (C2V_188_1071),
	.C2V_6 (C2V_193_1071),
	.L (L[16064:16050]),
	.V2C_1 (V2C_1071_22),
	.V2C_2 (V2C_1071_59),
	.V2C_3 (V2C_1071_81),
	.V2C_4 (V2C_1071_102),
	.V2C_5 (V2C_1071_188),
	.V2C_6 (V2C_1071_193),
	.V (V_1071)
);

VNU_6 #(quan_width) VNU1072 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_1072),
	.C2V_2 (C2V_65_1072),
	.C2V_3 (C2V_87_1072),
	.C2V_4 (C2V_108_1072),
	.C2V_5 (C2V_194_1072),
	.C2V_6 (C2V_199_1072),
	.L (L[16079:16065]),
	.V2C_1 (V2C_1072_28),
	.V2C_2 (V2C_1072_65),
	.V2C_3 (V2C_1072_87),
	.V2C_4 (V2C_1072_108),
	.V2C_5 (V2C_1072_194),
	.V2C_6 (V2C_1072_199),
	.V (V_1072)
);

VNU_6 #(quan_width) VNU1073 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_1073),
	.C2V_2 (C2V_71_1073),
	.C2V_3 (C2V_93_1073),
	.C2V_4 (C2V_114_1073),
	.C2V_5 (C2V_200_1073),
	.C2V_6 (C2V_205_1073),
	.L (L[16094:16080]),
	.V2C_1 (V2C_1073_34),
	.V2C_2 (V2C_1073_71),
	.V2C_3 (V2C_1073_93),
	.V2C_4 (V2C_1073_114),
	.V2C_5 (V2C_1073_200),
	.V2C_6 (V2C_1073_205),
	.V (V_1073)
);

VNU_6 #(quan_width) VNU1074 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_1074),
	.C2V_2 (C2V_77_1074),
	.C2V_3 (C2V_99_1074),
	.C2V_4 (C2V_120_1074),
	.C2V_5 (C2V_206_1074),
	.C2V_6 (C2V_211_1074),
	.L (L[16109:16095]),
	.V2C_1 (V2C_1074_40),
	.V2C_2 (V2C_1074_77),
	.V2C_3 (V2C_1074_99),
	.V2C_4 (V2C_1074_120),
	.V2C_5 (V2C_1074_206),
	.V2C_6 (V2C_1074_211),
	.V (V_1074)
);

VNU_6 #(quan_width) VNU1075 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_1075),
	.C2V_2 (C2V_83_1075),
	.C2V_3 (C2V_105_1075),
	.C2V_4 (C2V_126_1075),
	.C2V_5 (C2V_212_1075),
	.C2V_6 (C2V_217_1075),
	.L (L[16124:16110]),
	.V2C_1 (V2C_1075_46),
	.V2C_2 (V2C_1075_83),
	.V2C_3 (V2C_1075_105),
	.V2C_4 (V2C_1075_126),
	.V2C_5 (V2C_1075_212),
	.V2C_6 (V2C_1075_217),
	.V (V_1075)
);

VNU_6 #(quan_width) VNU1076 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_1076),
	.C2V_2 (C2V_89_1076),
	.C2V_3 (C2V_111_1076),
	.C2V_4 (C2V_132_1076),
	.C2V_5 (C2V_218_1076),
	.C2V_6 (C2V_223_1076),
	.L (L[16139:16125]),
	.V2C_1 (V2C_1076_52),
	.V2C_2 (V2C_1076_89),
	.V2C_3 (V2C_1076_111),
	.V2C_4 (V2C_1076_132),
	.V2C_5 (V2C_1076_218),
	.V2C_6 (V2C_1076_223),
	.V (V_1076)
);

VNU_6 #(quan_width) VNU1077 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_1077),
	.C2V_2 (C2V_95_1077),
	.C2V_3 (C2V_117_1077),
	.C2V_4 (C2V_138_1077),
	.C2V_5 (C2V_224_1077),
	.C2V_6 (C2V_229_1077),
	.L (L[16154:16140]),
	.V2C_1 (V2C_1077_58),
	.V2C_2 (V2C_1077_95),
	.V2C_3 (V2C_1077_117),
	.V2C_4 (V2C_1077_138),
	.V2C_5 (V2C_1077_224),
	.V2C_6 (V2C_1077_229),
	.V (V_1077)
);

VNU_6 #(quan_width) VNU1078 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_1078),
	.C2V_2 (C2V_101_1078),
	.C2V_3 (C2V_123_1078),
	.C2V_4 (C2V_144_1078),
	.C2V_5 (C2V_230_1078),
	.C2V_6 (C2V_235_1078),
	.L (L[16169:16155]),
	.V2C_1 (V2C_1078_64),
	.V2C_2 (V2C_1078_101),
	.V2C_3 (V2C_1078_123),
	.V2C_4 (V2C_1078_144),
	.V2C_5 (V2C_1078_230),
	.V2C_6 (V2C_1078_235),
	.V (V_1078)
);

VNU_6 #(quan_width) VNU1079 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_1079),
	.C2V_2 (C2V_107_1079),
	.C2V_3 (C2V_129_1079),
	.C2V_4 (C2V_150_1079),
	.C2V_5 (C2V_236_1079),
	.C2V_6 (C2V_241_1079),
	.L (L[16184:16170]),
	.V2C_1 (V2C_1079_70),
	.V2C_2 (V2C_1079_107),
	.V2C_3 (V2C_1079_129),
	.V2C_4 (V2C_1079_150),
	.V2C_5 (V2C_1079_236),
	.V2C_6 (V2C_1079_241),
	.V (V_1079)
);

VNU_6 #(quan_width) VNU1080 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_1080),
	.C2V_2 (C2V_113_1080),
	.C2V_3 (C2V_135_1080),
	.C2V_4 (C2V_156_1080),
	.C2V_5 (C2V_242_1080),
	.C2V_6 (C2V_247_1080),
	.L (L[16199:16185]),
	.V2C_1 (V2C_1080_76),
	.V2C_2 (V2C_1080_113),
	.V2C_3 (V2C_1080_135),
	.V2C_4 (V2C_1080_156),
	.V2C_5 (V2C_1080_242),
	.V2C_6 (V2C_1080_247),
	.V (V_1080)
);

VNU_6 #(quan_width) VNU1081 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_1081),
	.C2V_2 (C2V_119_1081),
	.C2V_3 (C2V_141_1081),
	.C2V_4 (C2V_162_1081),
	.C2V_5 (C2V_248_1081),
	.C2V_6 (C2V_253_1081),
	.L (L[16214:16200]),
	.V2C_1 (V2C_1081_82),
	.V2C_2 (V2C_1081_119),
	.V2C_3 (V2C_1081_141),
	.V2C_4 (V2C_1081_162),
	.V2C_5 (V2C_1081_248),
	.V2C_6 (V2C_1081_253),
	.V (V_1081)
);

VNU_6 #(quan_width) VNU1082 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_1082),
	.C2V_2 (C2V_125_1082),
	.C2V_3 (C2V_147_1082),
	.C2V_4 (C2V_168_1082),
	.C2V_5 (C2V_254_1082),
	.C2V_6 (C2V_259_1082),
	.L (L[16229:16215]),
	.V2C_1 (V2C_1082_88),
	.V2C_2 (V2C_1082_125),
	.V2C_3 (V2C_1082_147),
	.V2C_4 (V2C_1082_168),
	.V2C_5 (V2C_1082_254),
	.V2C_6 (V2C_1082_259),
	.V (V_1082)
);

VNU_6 #(quan_width) VNU1083 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_1083),
	.C2V_2 (C2V_131_1083),
	.C2V_3 (C2V_153_1083),
	.C2V_4 (C2V_174_1083),
	.C2V_5 (C2V_260_1083),
	.C2V_6 (C2V_265_1083),
	.L (L[16244:16230]),
	.V2C_1 (V2C_1083_94),
	.V2C_2 (V2C_1083_131),
	.V2C_3 (V2C_1083_153),
	.V2C_4 (V2C_1083_174),
	.V2C_5 (V2C_1083_260),
	.V2C_6 (V2C_1083_265),
	.V (V_1083)
);

VNU_6 #(quan_width) VNU1084 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_1084),
	.C2V_2 (C2V_137_1084),
	.C2V_3 (C2V_159_1084),
	.C2V_4 (C2V_180_1084),
	.C2V_5 (C2V_266_1084),
	.C2V_6 (C2V_271_1084),
	.L (L[16259:16245]),
	.V2C_1 (V2C_1084_100),
	.V2C_2 (V2C_1084_137),
	.V2C_3 (V2C_1084_159),
	.V2C_4 (V2C_1084_180),
	.V2C_5 (V2C_1084_266),
	.V2C_6 (V2C_1084_271),
	.V (V_1084)
);

VNU_6 #(quan_width) VNU1085 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_1085),
	.C2V_2 (C2V_143_1085),
	.C2V_3 (C2V_165_1085),
	.C2V_4 (C2V_186_1085),
	.C2V_5 (C2V_272_1085),
	.C2V_6 (C2V_277_1085),
	.L (L[16274:16260]),
	.V2C_1 (V2C_1085_106),
	.V2C_2 (V2C_1085_143),
	.V2C_3 (V2C_1085_165),
	.V2C_4 (V2C_1085_186),
	.V2C_5 (V2C_1085_272),
	.V2C_6 (V2C_1085_277),
	.V (V_1085)
);

VNU_6 #(quan_width) VNU1086 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_1086),
	.C2V_2 (C2V_149_1086),
	.C2V_3 (C2V_171_1086),
	.C2V_4 (C2V_192_1086),
	.C2V_5 (C2V_278_1086),
	.C2V_6 (C2V_283_1086),
	.L (L[16289:16275]),
	.V2C_1 (V2C_1086_112),
	.V2C_2 (V2C_1086_149),
	.V2C_3 (V2C_1086_171),
	.V2C_4 (V2C_1086_192),
	.V2C_5 (V2C_1086_278),
	.V2C_6 (V2C_1086_283),
	.V (V_1086)
);

VNU_6 #(quan_width) VNU1087 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_1087),
	.C2V_2 (C2V_118_1087),
	.C2V_3 (C2V_155_1087),
	.C2V_4 (C2V_177_1087),
	.C2V_5 (C2V_198_1087),
	.C2V_6 (C2V_284_1087),
	.L (L[16304:16290]),
	.V2C_1 (V2C_1087_1),
	.V2C_2 (V2C_1087_118),
	.V2C_3 (V2C_1087_155),
	.V2C_4 (V2C_1087_177),
	.V2C_5 (V2C_1087_198),
	.V2C_6 (V2C_1087_284),
	.V (V_1087)
);

VNU_6 #(quan_width) VNU1088 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_1088),
	.C2V_2 (C2V_7_1088),
	.C2V_3 (C2V_124_1088),
	.C2V_4 (C2V_161_1088),
	.C2V_5 (C2V_183_1088),
	.C2V_6 (C2V_204_1088),
	.L (L[16319:16305]),
	.V2C_1 (V2C_1088_2),
	.V2C_2 (V2C_1088_7),
	.V2C_3 (V2C_1088_124),
	.V2C_4 (V2C_1088_161),
	.V2C_5 (V2C_1088_183),
	.V2C_6 (V2C_1088_204),
	.V (V_1088)
);

VNU_6 #(quan_width) VNU1089 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_1089),
	.C2V_2 (C2V_13_1089),
	.C2V_3 (C2V_130_1089),
	.C2V_4 (C2V_167_1089),
	.C2V_5 (C2V_189_1089),
	.C2V_6 (C2V_210_1089),
	.L (L[16334:16320]),
	.V2C_1 (V2C_1089_8),
	.V2C_2 (V2C_1089_13),
	.V2C_3 (V2C_1089_130),
	.V2C_4 (V2C_1089_167),
	.V2C_5 (V2C_1089_189),
	.V2C_6 (V2C_1089_210),
	.V (V_1089)
);

VNU_6 #(quan_width) VNU1090 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_1090),
	.C2V_2 (C2V_19_1090),
	.C2V_3 (C2V_136_1090),
	.C2V_4 (C2V_173_1090),
	.C2V_5 (C2V_195_1090),
	.C2V_6 (C2V_216_1090),
	.L (L[16349:16335]),
	.V2C_1 (V2C_1090_14),
	.V2C_2 (V2C_1090_19),
	.V2C_3 (V2C_1090_136),
	.V2C_4 (V2C_1090_173),
	.V2C_5 (V2C_1090_195),
	.V2C_6 (V2C_1090_216),
	.V (V_1090)
);

VNU_6 #(quan_width) VNU1091 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_1091),
	.C2V_2 (C2V_25_1091),
	.C2V_3 (C2V_142_1091),
	.C2V_4 (C2V_179_1091),
	.C2V_5 (C2V_201_1091),
	.C2V_6 (C2V_222_1091),
	.L (L[16364:16350]),
	.V2C_1 (V2C_1091_20),
	.V2C_2 (V2C_1091_25),
	.V2C_3 (V2C_1091_142),
	.V2C_4 (V2C_1091_179),
	.V2C_5 (V2C_1091_201),
	.V2C_6 (V2C_1091_222),
	.V (V_1091)
);

VNU_6 #(quan_width) VNU1092 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_1092),
	.C2V_2 (C2V_31_1092),
	.C2V_3 (C2V_148_1092),
	.C2V_4 (C2V_185_1092),
	.C2V_5 (C2V_207_1092),
	.C2V_6 (C2V_228_1092),
	.L (L[16379:16365]),
	.V2C_1 (V2C_1092_26),
	.V2C_2 (V2C_1092_31),
	.V2C_3 (V2C_1092_148),
	.V2C_4 (V2C_1092_185),
	.V2C_5 (V2C_1092_207),
	.V2C_6 (V2C_1092_228),
	.V (V_1092)
);

VNU_6 #(quan_width) VNU1093 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_1093),
	.C2V_2 (C2V_37_1093),
	.C2V_3 (C2V_154_1093),
	.C2V_4 (C2V_191_1093),
	.C2V_5 (C2V_213_1093),
	.C2V_6 (C2V_234_1093),
	.L (L[16394:16380]),
	.V2C_1 (V2C_1093_32),
	.V2C_2 (V2C_1093_37),
	.V2C_3 (V2C_1093_154),
	.V2C_4 (V2C_1093_191),
	.V2C_5 (V2C_1093_213),
	.V2C_6 (V2C_1093_234),
	.V (V_1093)
);

VNU_6 #(quan_width) VNU1094 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_1094),
	.C2V_2 (C2V_43_1094),
	.C2V_3 (C2V_160_1094),
	.C2V_4 (C2V_197_1094),
	.C2V_5 (C2V_219_1094),
	.C2V_6 (C2V_240_1094),
	.L (L[16409:16395]),
	.V2C_1 (V2C_1094_38),
	.V2C_2 (V2C_1094_43),
	.V2C_3 (V2C_1094_160),
	.V2C_4 (V2C_1094_197),
	.V2C_5 (V2C_1094_219),
	.V2C_6 (V2C_1094_240),
	.V (V_1094)
);

VNU_6 #(quan_width) VNU1095 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_1095),
	.C2V_2 (C2V_49_1095),
	.C2V_3 (C2V_166_1095),
	.C2V_4 (C2V_203_1095),
	.C2V_5 (C2V_225_1095),
	.C2V_6 (C2V_246_1095),
	.L (L[16424:16410]),
	.V2C_1 (V2C_1095_44),
	.V2C_2 (V2C_1095_49),
	.V2C_3 (V2C_1095_166),
	.V2C_4 (V2C_1095_203),
	.V2C_5 (V2C_1095_225),
	.V2C_6 (V2C_1095_246),
	.V (V_1095)
);

VNU_6 #(quan_width) VNU1096 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_1096),
	.C2V_2 (C2V_55_1096),
	.C2V_3 (C2V_172_1096),
	.C2V_4 (C2V_209_1096),
	.C2V_5 (C2V_231_1096),
	.C2V_6 (C2V_252_1096),
	.L (L[16439:16425]),
	.V2C_1 (V2C_1096_50),
	.V2C_2 (V2C_1096_55),
	.V2C_3 (V2C_1096_172),
	.V2C_4 (V2C_1096_209),
	.V2C_5 (V2C_1096_231),
	.V2C_6 (V2C_1096_252),
	.V (V_1096)
);

VNU_6 #(quan_width) VNU1097 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_1097),
	.C2V_2 (C2V_61_1097),
	.C2V_3 (C2V_178_1097),
	.C2V_4 (C2V_215_1097),
	.C2V_5 (C2V_237_1097),
	.C2V_6 (C2V_258_1097),
	.L (L[16454:16440]),
	.V2C_1 (V2C_1097_56),
	.V2C_2 (V2C_1097_61),
	.V2C_3 (V2C_1097_178),
	.V2C_4 (V2C_1097_215),
	.V2C_5 (V2C_1097_237),
	.V2C_6 (V2C_1097_258),
	.V (V_1097)
);

VNU_6 #(quan_width) VNU1098 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_1098),
	.C2V_2 (C2V_67_1098),
	.C2V_3 (C2V_184_1098),
	.C2V_4 (C2V_221_1098),
	.C2V_5 (C2V_243_1098),
	.C2V_6 (C2V_264_1098),
	.L (L[16469:16455]),
	.V2C_1 (V2C_1098_62),
	.V2C_2 (V2C_1098_67),
	.V2C_3 (V2C_1098_184),
	.V2C_4 (V2C_1098_221),
	.V2C_5 (V2C_1098_243),
	.V2C_6 (V2C_1098_264),
	.V (V_1098)
);

VNU_6 #(quan_width) VNU1099 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_1099),
	.C2V_2 (C2V_73_1099),
	.C2V_3 (C2V_190_1099),
	.C2V_4 (C2V_227_1099),
	.C2V_5 (C2V_249_1099),
	.C2V_6 (C2V_270_1099),
	.L (L[16484:16470]),
	.V2C_1 (V2C_1099_68),
	.V2C_2 (V2C_1099_73),
	.V2C_3 (V2C_1099_190),
	.V2C_4 (V2C_1099_227),
	.V2C_5 (V2C_1099_249),
	.V2C_6 (V2C_1099_270),
	.V (V_1099)
);

VNU_6 #(quan_width) VNU1100 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_1100),
	.C2V_2 (C2V_79_1100),
	.C2V_3 (C2V_196_1100),
	.C2V_4 (C2V_233_1100),
	.C2V_5 (C2V_255_1100),
	.C2V_6 (C2V_276_1100),
	.L (L[16499:16485]),
	.V2C_1 (V2C_1100_74),
	.V2C_2 (V2C_1100_79),
	.V2C_3 (V2C_1100_196),
	.V2C_4 (V2C_1100_233),
	.V2C_5 (V2C_1100_255),
	.V2C_6 (V2C_1100_276),
	.V (V_1100)
);

VNU_6 #(quan_width) VNU1101 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_80_1101),
	.C2V_2 (C2V_85_1101),
	.C2V_3 (C2V_202_1101),
	.C2V_4 (C2V_239_1101),
	.C2V_5 (C2V_261_1101),
	.C2V_6 (C2V_282_1101),
	.L (L[16514:16500]),
	.V2C_1 (V2C_1101_80),
	.V2C_2 (V2C_1101_85),
	.V2C_3 (V2C_1101_202),
	.V2C_4 (V2C_1101_239),
	.V2C_5 (V2C_1101_261),
	.V2C_6 (V2C_1101_282),
	.V (V_1101)
);

VNU_6 #(quan_width) VNU1102 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_86_1102),
	.C2V_2 (C2V_91_1102),
	.C2V_3 (C2V_208_1102),
	.C2V_4 (C2V_245_1102),
	.C2V_5 (C2V_267_1102),
	.C2V_6 (C2V_288_1102),
	.L (L[16529:16515]),
	.V2C_1 (V2C_1102_86),
	.V2C_2 (V2C_1102_91),
	.V2C_3 (V2C_1102_208),
	.V2C_4 (V2C_1102_245),
	.V2C_5 (V2C_1102_267),
	.V2C_6 (V2C_1102_288),
	.V (V_1102)
);

VNU_6 #(quan_width) VNU1103 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_1103),
	.C2V_2 (C2V_92_1103),
	.C2V_3 (C2V_97_1103),
	.C2V_4 (C2V_214_1103),
	.C2V_5 (C2V_251_1103),
	.C2V_6 (C2V_273_1103),
	.L (L[16544:16530]),
	.V2C_1 (V2C_1103_6),
	.V2C_2 (V2C_1103_92),
	.V2C_3 (V2C_1103_97),
	.V2C_4 (V2C_1103_214),
	.V2C_5 (V2C_1103_251),
	.V2C_6 (V2C_1103_273),
	.V (V_1103)
);

VNU_6 #(quan_width) VNU1104 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_1104),
	.C2V_2 (C2V_98_1104),
	.C2V_3 (C2V_103_1104),
	.C2V_4 (C2V_220_1104),
	.C2V_5 (C2V_257_1104),
	.C2V_6 (C2V_279_1104),
	.L (L[16559:16545]),
	.V2C_1 (V2C_1104_12),
	.V2C_2 (V2C_1104_98),
	.V2C_3 (V2C_1104_103),
	.V2C_4 (V2C_1104_220),
	.V2C_5 (V2C_1104_257),
	.V2C_6 (V2C_1104_279),
	.V (V_1104)
);

VNU_6 #(quan_width) VNU1105 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_1105),
	.C2V_2 (C2V_15_1105),
	.C2V_3 (C2V_43_1105),
	.C2V_4 (C2V_130_1105),
	.C2V_5 (C2V_206_1105),
	.C2V_6 (C2V_263_1105),
	.L (L[16574:16560]),
	.V2C_1 (V2C_1105_6),
	.V2C_2 (V2C_1105_15),
	.V2C_3 (V2C_1105_43),
	.V2C_4 (V2C_1105_130),
	.V2C_5 (V2C_1105_206),
	.V2C_6 (V2C_1105_263),
	.V (V_1105)
);

VNU_6 #(quan_width) VNU1106 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_1106),
	.C2V_2 (C2V_21_1106),
	.C2V_3 (C2V_49_1106),
	.C2V_4 (C2V_136_1106),
	.C2V_5 (C2V_212_1106),
	.C2V_6 (C2V_269_1106),
	.L (L[16589:16575]),
	.V2C_1 (V2C_1106_12),
	.V2C_2 (V2C_1106_21),
	.V2C_3 (V2C_1106_49),
	.V2C_4 (V2C_1106_136),
	.V2C_5 (V2C_1106_212),
	.V2C_6 (V2C_1106_269),
	.V (V_1106)
);

VNU_6 #(quan_width) VNU1107 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_1107),
	.C2V_2 (C2V_27_1107),
	.C2V_3 (C2V_55_1107),
	.C2V_4 (C2V_142_1107),
	.C2V_5 (C2V_218_1107),
	.C2V_6 (C2V_275_1107),
	.L (L[16604:16590]),
	.V2C_1 (V2C_1107_18),
	.V2C_2 (V2C_1107_27),
	.V2C_3 (V2C_1107_55),
	.V2C_4 (V2C_1107_142),
	.V2C_5 (V2C_1107_218),
	.V2C_6 (V2C_1107_275),
	.V (V_1107)
);

VNU_6 #(quan_width) VNU1108 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_1108),
	.C2V_2 (C2V_33_1108),
	.C2V_3 (C2V_61_1108),
	.C2V_4 (C2V_148_1108),
	.C2V_5 (C2V_224_1108),
	.C2V_6 (C2V_281_1108),
	.L (L[16619:16605]),
	.V2C_1 (V2C_1108_24),
	.V2C_2 (V2C_1108_33),
	.V2C_3 (V2C_1108_61),
	.V2C_4 (V2C_1108_148),
	.V2C_5 (V2C_1108_224),
	.V2C_6 (V2C_1108_281),
	.V (V_1108)
);

VNU_6 #(quan_width) VNU1109 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_1109),
	.C2V_2 (C2V_39_1109),
	.C2V_3 (C2V_67_1109),
	.C2V_4 (C2V_154_1109),
	.C2V_5 (C2V_230_1109),
	.C2V_6 (C2V_287_1109),
	.L (L[16634:16620]),
	.V2C_1 (V2C_1109_30),
	.V2C_2 (V2C_1109_39),
	.V2C_3 (V2C_1109_67),
	.V2C_4 (V2C_1109_154),
	.V2C_5 (V2C_1109_230),
	.V2C_6 (V2C_1109_287),
	.V (V_1109)
);

VNU_6 #(quan_width) VNU1110 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_1110),
	.C2V_2 (C2V_36_1110),
	.C2V_3 (C2V_45_1110),
	.C2V_4 (C2V_73_1110),
	.C2V_5 (C2V_160_1110),
	.C2V_6 (C2V_236_1110),
	.L (L[16649:16635]),
	.V2C_1 (V2C_1110_5),
	.V2C_2 (V2C_1110_36),
	.V2C_3 (V2C_1110_45),
	.V2C_4 (V2C_1110_73),
	.V2C_5 (V2C_1110_160),
	.V2C_6 (V2C_1110_236),
	.V (V_1110)
);

VNU_6 #(quan_width) VNU1111 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_1111),
	.C2V_2 (C2V_42_1111),
	.C2V_3 (C2V_51_1111),
	.C2V_4 (C2V_79_1111),
	.C2V_5 (C2V_166_1111),
	.C2V_6 (C2V_242_1111),
	.L (L[16664:16650]),
	.V2C_1 (V2C_1111_11),
	.V2C_2 (V2C_1111_42),
	.V2C_3 (V2C_1111_51),
	.V2C_4 (V2C_1111_79),
	.V2C_5 (V2C_1111_166),
	.V2C_6 (V2C_1111_242),
	.V (V_1111)
);

VNU_6 #(quan_width) VNU1112 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_1112),
	.C2V_2 (C2V_48_1112),
	.C2V_3 (C2V_57_1112),
	.C2V_4 (C2V_85_1112),
	.C2V_5 (C2V_172_1112),
	.C2V_6 (C2V_248_1112),
	.L (L[16679:16665]),
	.V2C_1 (V2C_1112_17),
	.V2C_2 (V2C_1112_48),
	.V2C_3 (V2C_1112_57),
	.V2C_4 (V2C_1112_85),
	.V2C_5 (V2C_1112_172),
	.V2C_6 (V2C_1112_248),
	.V (V_1112)
);

VNU_6 #(quan_width) VNU1113 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_1113),
	.C2V_2 (C2V_54_1113),
	.C2V_3 (C2V_63_1113),
	.C2V_4 (C2V_91_1113),
	.C2V_5 (C2V_178_1113),
	.C2V_6 (C2V_254_1113),
	.L (L[16694:16680]),
	.V2C_1 (V2C_1113_23),
	.V2C_2 (V2C_1113_54),
	.V2C_3 (V2C_1113_63),
	.V2C_4 (V2C_1113_91),
	.V2C_5 (V2C_1113_178),
	.V2C_6 (V2C_1113_254),
	.V (V_1113)
);

VNU_6 #(quan_width) VNU1114 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_1114),
	.C2V_2 (C2V_60_1114),
	.C2V_3 (C2V_69_1114),
	.C2V_4 (C2V_97_1114),
	.C2V_5 (C2V_184_1114),
	.C2V_6 (C2V_260_1114),
	.L (L[16709:16695]),
	.V2C_1 (V2C_1114_29),
	.V2C_2 (V2C_1114_60),
	.V2C_3 (V2C_1114_69),
	.V2C_4 (V2C_1114_97),
	.V2C_5 (V2C_1114_184),
	.V2C_6 (V2C_1114_260),
	.V (V_1114)
);

VNU_6 #(quan_width) VNU1115 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_1115),
	.C2V_2 (C2V_66_1115),
	.C2V_3 (C2V_75_1115),
	.C2V_4 (C2V_103_1115),
	.C2V_5 (C2V_190_1115),
	.C2V_6 (C2V_266_1115),
	.L (L[16724:16710]),
	.V2C_1 (V2C_1115_35),
	.V2C_2 (V2C_1115_66),
	.V2C_3 (V2C_1115_75),
	.V2C_4 (V2C_1115_103),
	.V2C_5 (V2C_1115_190),
	.V2C_6 (V2C_1115_266),
	.V (V_1115)
);

VNU_6 #(quan_width) VNU1116 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_1116),
	.C2V_2 (C2V_72_1116),
	.C2V_3 (C2V_81_1116),
	.C2V_4 (C2V_109_1116),
	.C2V_5 (C2V_196_1116),
	.C2V_6 (C2V_272_1116),
	.L (L[16739:16725]),
	.V2C_1 (V2C_1116_41),
	.V2C_2 (V2C_1116_72),
	.V2C_3 (V2C_1116_81),
	.V2C_4 (V2C_1116_109),
	.V2C_5 (V2C_1116_196),
	.V2C_6 (V2C_1116_272),
	.V (V_1116)
);

VNU_6 #(quan_width) VNU1117 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_1117),
	.C2V_2 (C2V_78_1117),
	.C2V_3 (C2V_87_1117),
	.C2V_4 (C2V_115_1117),
	.C2V_5 (C2V_202_1117),
	.C2V_6 (C2V_278_1117),
	.L (L[16754:16740]),
	.V2C_1 (V2C_1117_47),
	.V2C_2 (V2C_1117_78),
	.V2C_3 (V2C_1117_87),
	.V2C_4 (V2C_1117_115),
	.V2C_5 (V2C_1117_202),
	.V2C_6 (V2C_1117_278),
	.V (V_1117)
);

VNU_6 #(quan_width) VNU1118 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_1118),
	.C2V_2 (C2V_84_1118),
	.C2V_3 (C2V_93_1118),
	.C2V_4 (C2V_121_1118),
	.C2V_5 (C2V_208_1118),
	.C2V_6 (C2V_284_1118),
	.L (L[16769:16755]),
	.V2C_1 (V2C_1118_53),
	.V2C_2 (V2C_1118_84),
	.V2C_3 (V2C_1118_93),
	.V2C_4 (V2C_1118_121),
	.V2C_5 (V2C_1118_208),
	.V2C_6 (V2C_1118_284),
	.V (V_1118)
);

VNU_6 #(quan_width) VNU1119 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_1119),
	.C2V_2 (C2V_59_1119),
	.C2V_3 (C2V_90_1119),
	.C2V_4 (C2V_99_1119),
	.C2V_5 (C2V_127_1119),
	.C2V_6 (C2V_214_1119),
	.L (L[16784:16770]),
	.V2C_1 (V2C_1119_2),
	.V2C_2 (V2C_1119_59),
	.V2C_3 (V2C_1119_90),
	.V2C_4 (V2C_1119_99),
	.V2C_5 (V2C_1119_127),
	.V2C_6 (V2C_1119_214),
	.V (V_1119)
);

VNU_6 #(quan_width) VNU1120 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_1120),
	.C2V_2 (C2V_65_1120),
	.C2V_3 (C2V_96_1120),
	.C2V_4 (C2V_105_1120),
	.C2V_5 (C2V_133_1120),
	.C2V_6 (C2V_220_1120),
	.L (L[16799:16785]),
	.V2C_1 (V2C_1120_8),
	.V2C_2 (V2C_1120_65),
	.V2C_3 (V2C_1120_96),
	.V2C_4 (V2C_1120_105),
	.V2C_5 (V2C_1120_133),
	.V2C_6 (V2C_1120_220),
	.V (V_1120)
);

VNU_6 #(quan_width) VNU1121 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_1121),
	.C2V_2 (C2V_71_1121),
	.C2V_3 (C2V_102_1121),
	.C2V_4 (C2V_111_1121),
	.C2V_5 (C2V_139_1121),
	.C2V_6 (C2V_226_1121),
	.L (L[16814:16800]),
	.V2C_1 (V2C_1121_14),
	.V2C_2 (V2C_1121_71),
	.V2C_3 (V2C_1121_102),
	.V2C_4 (V2C_1121_111),
	.V2C_5 (V2C_1121_139),
	.V2C_6 (V2C_1121_226),
	.V (V_1121)
);

VNU_6 #(quan_width) VNU1122 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_1122),
	.C2V_2 (C2V_77_1122),
	.C2V_3 (C2V_108_1122),
	.C2V_4 (C2V_117_1122),
	.C2V_5 (C2V_145_1122),
	.C2V_6 (C2V_232_1122),
	.L (L[16829:16815]),
	.V2C_1 (V2C_1122_20),
	.V2C_2 (V2C_1122_77),
	.V2C_3 (V2C_1122_108),
	.V2C_4 (V2C_1122_117),
	.V2C_5 (V2C_1122_145),
	.V2C_6 (V2C_1122_232),
	.V (V_1122)
);

VNU_6 #(quan_width) VNU1123 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_1123),
	.C2V_2 (C2V_83_1123),
	.C2V_3 (C2V_114_1123),
	.C2V_4 (C2V_123_1123),
	.C2V_5 (C2V_151_1123),
	.C2V_6 (C2V_238_1123),
	.L (L[16844:16830]),
	.V2C_1 (V2C_1123_26),
	.V2C_2 (V2C_1123_83),
	.V2C_3 (V2C_1123_114),
	.V2C_4 (V2C_1123_123),
	.V2C_5 (V2C_1123_151),
	.V2C_6 (V2C_1123_238),
	.V (V_1123)
);

VNU_6 #(quan_width) VNU1124 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_1124),
	.C2V_2 (C2V_89_1124),
	.C2V_3 (C2V_120_1124),
	.C2V_4 (C2V_129_1124),
	.C2V_5 (C2V_157_1124),
	.C2V_6 (C2V_244_1124),
	.L (L[16859:16845]),
	.V2C_1 (V2C_1124_32),
	.V2C_2 (V2C_1124_89),
	.V2C_3 (V2C_1124_120),
	.V2C_4 (V2C_1124_129),
	.V2C_5 (V2C_1124_157),
	.V2C_6 (V2C_1124_244),
	.V (V_1124)
);

VNU_6 #(quan_width) VNU1125 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_1125),
	.C2V_2 (C2V_95_1125),
	.C2V_3 (C2V_126_1125),
	.C2V_4 (C2V_135_1125),
	.C2V_5 (C2V_163_1125),
	.C2V_6 (C2V_250_1125),
	.L (L[16874:16860]),
	.V2C_1 (V2C_1125_38),
	.V2C_2 (V2C_1125_95),
	.V2C_3 (V2C_1125_126),
	.V2C_4 (V2C_1125_135),
	.V2C_5 (V2C_1125_163),
	.V2C_6 (V2C_1125_250),
	.V (V_1125)
);

VNU_6 #(quan_width) VNU1126 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_1126),
	.C2V_2 (C2V_101_1126),
	.C2V_3 (C2V_132_1126),
	.C2V_4 (C2V_141_1126),
	.C2V_5 (C2V_169_1126),
	.C2V_6 (C2V_256_1126),
	.L (L[16889:16875]),
	.V2C_1 (V2C_1126_44),
	.V2C_2 (V2C_1126_101),
	.V2C_3 (V2C_1126_132),
	.V2C_4 (V2C_1126_141),
	.V2C_5 (V2C_1126_169),
	.V2C_6 (V2C_1126_256),
	.V (V_1126)
);

VNU_6 #(quan_width) VNU1127 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_1127),
	.C2V_2 (C2V_107_1127),
	.C2V_3 (C2V_138_1127),
	.C2V_4 (C2V_147_1127),
	.C2V_5 (C2V_175_1127),
	.C2V_6 (C2V_262_1127),
	.L (L[16904:16890]),
	.V2C_1 (V2C_1127_50),
	.V2C_2 (V2C_1127_107),
	.V2C_3 (V2C_1127_138),
	.V2C_4 (V2C_1127_147),
	.V2C_5 (V2C_1127_175),
	.V2C_6 (V2C_1127_262),
	.V (V_1127)
);

VNU_6 #(quan_width) VNU1128 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_1128),
	.C2V_2 (C2V_113_1128),
	.C2V_3 (C2V_144_1128),
	.C2V_4 (C2V_153_1128),
	.C2V_5 (C2V_181_1128),
	.C2V_6 (C2V_268_1128),
	.L (L[16919:16905]),
	.V2C_1 (V2C_1128_56),
	.V2C_2 (V2C_1128_113),
	.V2C_3 (V2C_1128_144),
	.V2C_4 (V2C_1128_153),
	.V2C_5 (V2C_1128_181),
	.V2C_6 (V2C_1128_268),
	.V (V_1128)
);

VNU_6 #(quan_width) VNU1129 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_1129),
	.C2V_2 (C2V_119_1129),
	.C2V_3 (C2V_150_1129),
	.C2V_4 (C2V_159_1129),
	.C2V_5 (C2V_187_1129),
	.C2V_6 (C2V_274_1129),
	.L (L[16934:16920]),
	.V2C_1 (V2C_1129_62),
	.V2C_2 (V2C_1129_119),
	.V2C_3 (V2C_1129_150),
	.V2C_4 (V2C_1129_159),
	.V2C_5 (V2C_1129_187),
	.V2C_6 (V2C_1129_274),
	.V (V_1129)
);

VNU_6 #(quan_width) VNU1130 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_1130),
	.C2V_2 (C2V_125_1130),
	.C2V_3 (C2V_156_1130),
	.C2V_4 (C2V_165_1130),
	.C2V_5 (C2V_193_1130),
	.C2V_6 (C2V_280_1130),
	.L (L[16949:16935]),
	.V2C_1 (V2C_1130_68),
	.V2C_2 (V2C_1130_125),
	.V2C_3 (V2C_1130_156),
	.V2C_4 (V2C_1130_165),
	.V2C_5 (V2C_1130_193),
	.V2C_6 (V2C_1130_280),
	.V (V_1130)
);

VNU_6 #(quan_width) VNU1131 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_1131),
	.C2V_2 (C2V_131_1131),
	.C2V_3 (C2V_162_1131),
	.C2V_4 (C2V_171_1131),
	.C2V_5 (C2V_199_1131),
	.C2V_6 (C2V_286_1131),
	.L (L[16964:16950]),
	.V2C_1 (V2C_1131_74),
	.V2C_2 (V2C_1131_131),
	.V2C_3 (V2C_1131_162),
	.V2C_4 (V2C_1131_171),
	.V2C_5 (V2C_1131_199),
	.V2C_6 (V2C_1131_286),
	.V (V_1131)
);

VNU_6 #(quan_width) VNU1132 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_1132),
	.C2V_2 (C2V_80_1132),
	.C2V_3 (C2V_137_1132),
	.C2V_4 (C2V_168_1132),
	.C2V_5 (C2V_177_1132),
	.C2V_6 (C2V_205_1132),
	.L (L[16979:16965]),
	.V2C_1 (V2C_1132_4),
	.V2C_2 (V2C_1132_80),
	.V2C_3 (V2C_1132_137),
	.V2C_4 (V2C_1132_168),
	.V2C_5 (V2C_1132_177),
	.V2C_6 (V2C_1132_205),
	.V (V_1132)
);

VNU_6 #(quan_width) VNU1133 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_1133),
	.C2V_2 (C2V_86_1133),
	.C2V_3 (C2V_143_1133),
	.C2V_4 (C2V_174_1133),
	.C2V_5 (C2V_183_1133),
	.C2V_6 (C2V_211_1133),
	.L (L[16994:16980]),
	.V2C_1 (V2C_1133_10),
	.V2C_2 (V2C_1133_86),
	.V2C_3 (V2C_1133_143),
	.V2C_4 (V2C_1133_174),
	.V2C_5 (V2C_1133_183),
	.V2C_6 (V2C_1133_211),
	.V (V_1133)
);

VNU_6 #(quan_width) VNU1134 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_1134),
	.C2V_2 (C2V_92_1134),
	.C2V_3 (C2V_149_1134),
	.C2V_4 (C2V_180_1134),
	.C2V_5 (C2V_189_1134),
	.C2V_6 (C2V_217_1134),
	.L (L[17009:16995]),
	.V2C_1 (V2C_1134_16),
	.V2C_2 (V2C_1134_92),
	.V2C_3 (V2C_1134_149),
	.V2C_4 (V2C_1134_180),
	.V2C_5 (V2C_1134_189),
	.V2C_6 (V2C_1134_217),
	.V (V_1134)
);

VNU_6 #(quan_width) VNU1135 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_1135),
	.C2V_2 (C2V_98_1135),
	.C2V_3 (C2V_155_1135),
	.C2V_4 (C2V_186_1135),
	.C2V_5 (C2V_195_1135),
	.C2V_6 (C2V_223_1135),
	.L (L[17024:17010]),
	.V2C_1 (V2C_1135_22),
	.V2C_2 (V2C_1135_98),
	.V2C_3 (V2C_1135_155),
	.V2C_4 (V2C_1135_186),
	.V2C_5 (V2C_1135_195),
	.V2C_6 (V2C_1135_223),
	.V (V_1135)
);

VNU_6 #(quan_width) VNU1136 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_1136),
	.C2V_2 (C2V_104_1136),
	.C2V_3 (C2V_161_1136),
	.C2V_4 (C2V_192_1136),
	.C2V_5 (C2V_201_1136),
	.C2V_6 (C2V_229_1136),
	.L (L[17039:17025]),
	.V2C_1 (V2C_1136_28),
	.V2C_2 (V2C_1136_104),
	.V2C_3 (V2C_1136_161),
	.V2C_4 (V2C_1136_192),
	.V2C_5 (V2C_1136_201),
	.V2C_6 (V2C_1136_229),
	.V (V_1136)
);

VNU_6 #(quan_width) VNU1137 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_1137),
	.C2V_2 (C2V_110_1137),
	.C2V_3 (C2V_167_1137),
	.C2V_4 (C2V_198_1137),
	.C2V_5 (C2V_207_1137),
	.C2V_6 (C2V_235_1137),
	.L (L[17054:17040]),
	.V2C_1 (V2C_1137_34),
	.V2C_2 (V2C_1137_110),
	.V2C_3 (V2C_1137_167),
	.V2C_4 (V2C_1137_198),
	.V2C_5 (V2C_1137_207),
	.V2C_6 (V2C_1137_235),
	.V (V_1137)
);

VNU_6 #(quan_width) VNU1138 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_1138),
	.C2V_2 (C2V_116_1138),
	.C2V_3 (C2V_173_1138),
	.C2V_4 (C2V_204_1138),
	.C2V_5 (C2V_213_1138),
	.C2V_6 (C2V_241_1138),
	.L (L[17069:17055]),
	.V2C_1 (V2C_1138_40),
	.V2C_2 (V2C_1138_116),
	.V2C_3 (V2C_1138_173),
	.V2C_4 (V2C_1138_204),
	.V2C_5 (V2C_1138_213),
	.V2C_6 (V2C_1138_241),
	.V (V_1138)
);

VNU_6 #(quan_width) VNU1139 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_1139),
	.C2V_2 (C2V_122_1139),
	.C2V_3 (C2V_179_1139),
	.C2V_4 (C2V_210_1139),
	.C2V_5 (C2V_219_1139),
	.C2V_6 (C2V_247_1139),
	.L (L[17084:17070]),
	.V2C_1 (V2C_1139_46),
	.V2C_2 (V2C_1139_122),
	.V2C_3 (V2C_1139_179),
	.V2C_4 (V2C_1139_210),
	.V2C_5 (V2C_1139_219),
	.V2C_6 (V2C_1139_247),
	.V (V_1139)
);

VNU_6 #(quan_width) VNU1140 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_1140),
	.C2V_2 (C2V_128_1140),
	.C2V_3 (C2V_185_1140),
	.C2V_4 (C2V_216_1140),
	.C2V_5 (C2V_225_1140),
	.C2V_6 (C2V_253_1140),
	.L (L[17099:17085]),
	.V2C_1 (V2C_1140_52),
	.V2C_2 (V2C_1140_128),
	.V2C_3 (V2C_1140_185),
	.V2C_4 (V2C_1140_216),
	.V2C_5 (V2C_1140_225),
	.V2C_6 (V2C_1140_253),
	.V (V_1140)
);

VNU_6 #(quan_width) VNU1141 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_1141),
	.C2V_2 (C2V_134_1141),
	.C2V_3 (C2V_191_1141),
	.C2V_4 (C2V_222_1141),
	.C2V_5 (C2V_231_1141),
	.C2V_6 (C2V_259_1141),
	.L (L[17114:17100]),
	.V2C_1 (V2C_1141_58),
	.V2C_2 (V2C_1141_134),
	.V2C_3 (V2C_1141_191),
	.V2C_4 (V2C_1141_222),
	.V2C_5 (V2C_1141_231),
	.V2C_6 (V2C_1141_259),
	.V (V_1141)
);

VNU_6 #(quan_width) VNU1142 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_1142),
	.C2V_2 (C2V_140_1142),
	.C2V_3 (C2V_197_1142),
	.C2V_4 (C2V_228_1142),
	.C2V_5 (C2V_237_1142),
	.C2V_6 (C2V_265_1142),
	.L (L[17129:17115]),
	.V2C_1 (V2C_1142_64),
	.V2C_2 (V2C_1142_140),
	.V2C_3 (V2C_1142_197),
	.V2C_4 (V2C_1142_228),
	.V2C_5 (V2C_1142_237),
	.V2C_6 (V2C_1142_265),
	.V (V_1142)
);

VNU_6 #(quan_width) VNU1143 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_1143),
	.C2V_2 (C2V_146_1143),
	.C2V_3 (C2V_203_1143),
	.C2V_4 (C2V_234_1143),
	.C2V_5 (C2V_243_1143),
	.C2V_6 (C2V_271_1143),
	.L (L[17144:17130]),
	.V2C_1 (V2C_1143_70),
	.V2C_2 (V2C_1143_146),
	.V2C_3 (V2C_1143_203),
	.V2C_4 (V2C_1143_234),
	.V2C_5 (V2C_1143_243),
	.V2C_6 (V2C_1143_271),
	.V (V_1143)
);

VNU_6 #(quan_width) VNU1144 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_1144),
	.C2V_2 (C2V_152_1144),
	.C2V_3 (C2V_209_1144),
	.C2V_4 (C2V_240_1144),
	.C2V_5 (C2V_249_1144),
	.C2V_6 (C2V_277_1144),
	.L (L[17159:17145]),
	.V2C_1 (V2C_1144_76),
	.V2C_2 (V2C_1144_152),
	.V2C_3 (V2C_1144_209),
	.V2C_4 (V2C_1144_240),
	.V2C_5 (V2C_1144_249),
	.V2C_6 (V2C_1144_277),
	.V (V_1144)
);

VNU_6 #(quan_width) VNU1145 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_1145),
	.C2V_2 (C2V_158_1145),
	.C2V_3 (C2V_215_1145),
	.C2V_4 (C2V_246_1145),
	.C2V_5 (C2V_255_1145),
	.C2V_6 (C2V_283_1145),
	.L (L[17174:17160]),
	.V2C_1 (V2C_1145_82),
	.V2C_2 (V2C_1145_158),
	.V2C_3 (V2C_1145_215),
	.V2C_4 (V2C_1145_246),
	.V2C_5 (V2C_1145_255),
	.V2C_6 (V2C_1145_283),
	.V (V_1145)
);

VNU_6 #(quan_width) VNU1146 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_1146),
	.C2V_2 (C2V_88_1146),
	.C2V_3 (C2V_164_1146),
	.C2V_4 (C2V_221_1146),
	.C2V_5 (C2V_252_1146),
	.C2V_6 (C2V_261_1146),
	.L (L[17189:17175]),
	.V2C_1 (V2C_1146_1),
	.V2C_2 (V2C_1146_88),
	.V2C_3 (V2C_1146_164),
	.V2C_4 (V2C_1146_221),
	.V2C_5 (V2C_1146_252),
	.V2C_6 (V2C_1146_261),
	.V (V_1146)
);

VNU_6 #(quan_width) VNU1147 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_1147),
	.C2V_2 (C2V_94_1147),
	.C2V_3 (C2V_170_1147),
	.C2V_4 (C2V_227_1147),
	.C2V_5 (C2V_258_1147),
	.C2V_6 (C2V_267_1147),
	.L (L[17204:17190]),
	.V2C_1 (V2C_1147_7),
	.V2C_2 (V2C_1147_94),
	.V2C_3 (V2C_1147_170),
	.V2C_4 (V2C_1147_227),
	.V2C_5 (V2C_1147_258),
	.V2C_6 (V2C_1147_267),
	.V (V_1147)
);

VNU_6 #(quan_width) VNU1148 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_1148),
	.C2V_2 (C2V_100_1148),
	.C2V_3 (C2V_176_1148),
	.C2V_4 (C2V_233_1148),
	.C2V_5 (C2V_264_1148),
	.C2V_6 (C2V_273_1148),
	.L (L[17219:17205]),
	.V2C_1 (V2C_1148_13),
	.V2C_2 (V2C_1148_100),
	.V2C_3 (V2C_1148_176),
	.V2C_4 (V2C_1148_233),
	.V2C_5 (V2C_1148_264),
	.V2C_6 (V2C_1148_273),
	.V (V_1148)
);

VNU_6 #(quan_width) VNU1149 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_1149),
	.C2V_2 (C2V_106_1149),
	.C2V_3 (C2V_182_1149),
	.C2V_4 (C2V_239_1149),
	.C2V_5 (C2V_270_1149),
	.C2V_6 (C2V_279_1149),
	.L (L[17234:17220]),
	.V2C_1 (V2C_1149_19),
	.V2C_2 (V2C_1149_106),
	.V2C_3 (V2C_1149_182),
	.V2C_4 (V2C_1149_239),
	.V2C_5 (V2C_1149_270),
	.V2C_6 (V2C_1149_279),
	.V (V_1149)
);

VNU_6 #(quan_width) VNU1150 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_1150),
	.C2V_2 (C2V_112_1150),
	.C2V_3 (C2V_188_1150),
	.C2V_4 (C2V_245_1150),
	.C2V_5 (C2V_276_1150),
	.C2V_6 (C2V_285_1150),
	.L (L[17249:17235]),
	.V2C_1 (V2C_1150_25),
	.V2C_2 (V2C_1150_112),
	.V2C_3 (V2C_1150_188),
	.V2C_4 (V2C_1150_245),
	.V2C_5 (V2C_1150_276),
	.V2C_6 (V2C_1150_285),
	.V (V_1150)
);

VNU_6 #(quan_width) VNU1151 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_1151),
	.C2V_2 (C2V_31_1151),
	.C2V_3 (C2V_118_1151),
	.C2V_4 (C2V_194_1151),
	.C2V_5 (C2V_251_1151),
	.C2V_6 (C2V_282_1151),
	.L (L[17264:17250]),
	.V2C_1 (V2C_1151_3),
	.V2C_2 (V2C_1151_31),
	.V2C_3 (V2C_1151_118),
	.V2C_4 (V2C_1151_194),
	.V2C_5 (V2C_1151_251),
	.V2C_6 (V2C_1151_282),
	.V (V_1151)
);

VNU_6 #(quan_width) VNU1152 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_1152),
	.C2V_2 (C2V_37_1152),
	.C2V_3 (C2V_124_1152),
	.C2V_4 (C2V_200_1152),
	.C2V_5 (C2V_257_1152),
	.C2V_6 (C2V_288_1152),
	.L (L[17279:17265]),
	.V2C_1 (V2C_1152_9),
	.V2C_2 (V2C_1152_37),
	.V2C_3 (V2C_1152_124),
	.V2C_4 (V2C_1152_200),
	.V2C_5 (V2C_1152_257),
	.V2C_6 (V2C_1152_288),
	.V (V_1152)
);

VNU_2 #(quan_width) VNU1153 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_1153),
	.C2V_2 (C2V_2_1153),
	.L (L[17294:17280]),
	.V2C_1 (V2C_1153_1),
	.V2C_2 (V2C_1153_2),
	.V (V_1153)
);

VNU_2 #(quan_width) VNU1154 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_1154),
	.C2V_2 (C2V_3_1154),
	.L (L[17309:17295]),
	.V2C_1 (V2C_1154_2),
	.V2C_2 (V2C_1154_3),
	.V (V_1154)
);

VNU_2 #(quan_width) VNU1155 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_1155),
	.C2V_2 (C2V_4_1155),
	.L (L[17324:17310]),
	.V2C_1 (V2C_1155_3),
	.V2C_2 (V2C_1155_4),
	.V (V_1155)
);

VNU_2 #(quan_width) VNU1156 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_1156),
	.C2V_2 (C2V_5_1156),
	.L (L[17339:17325]),
	.V2C_1 (V2C_1156_4),
	.V2C_2 (V2C_1156_5),
	.V (V_1156)
);

VNU_2 #(quan_width) VNU1157 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_1157),
	.C2V_2 (C2V_6_1157),
	.L (L[17354:17340]),
	.V2C_1 (V2C_1157_5),
	.V2C_2 (V2C_1157_6),
	.V (V_1157)
);

VNU_2 #(quan_width) VNU1158 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_1158),
	.C2V_2 (C2V_7_1158),
	.L (L[17369:17355]),
	.V2C_1 (V2C_1158_6),
	.V2C_2 (V2C_1158_7),
	.V (V_1158)
);

VNU_2 #(quan_width) VNU1159 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_1159),
	.C2V_2 (C2V_8_1159),
	.L (L[17384:17370]),
	.V2C_1 (V2C_1159_7),
	.V2C_2 (V2C_1159_8),
	.V (V_1159)
);

VNU_2 #(quan_width) VNU1160 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_1160),
	.C2V_2 (C2V_9_1160),
	.L (L[17399:17385]),
	.V2C_1 (V2C_1160_8),
	.V2C_2 (V2C_1160_9),
	.V (V_1160)
);

VNU_2 #(quan_width) VNU1161 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_1161),
	.C2V_2 (C2V_10_1161),
	.L (L[17414:17400]),
	.V2C_1 (V2C_1161_9),
	.V2C_2 (V2C_1161_10),
	.V (V_1161)
);

VNU_2 #(quan_width) VNU1162 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_1162),
	.C2V_2 (C2V_11_1162),
	.L (L[17429:17415]),
	.V2C_1 (V2C_1162_10),
	.V2C_2 (V2C_1162_11),
	.V (V_1162)
);

VNU_2 #(quan_width) VNU1163 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_1163),
	.C2V_2 (C2V_12_1163),
	.L (L[17444:17430]),
	.V2C_1 (V2C_1163_11),
	.V2C_2 (V2C_1163_12),
	.V (V_1163)
);

VNU_2 #(quan_width) VNU1164 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_1164),
	.C2V_2 (C2V_13_1164),
	.L (L[17459:17445]),
	.V2C_1 (V2C_1164_12),
	.V2C_2 (V2C_1164_13),
	.V (V_1164)
);

VNU_2 #(quan_width) VNU1165 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_1165),
	.C2V_2 (C2V_14_1165),
	.L (L[17474:17460]),
	.V2C_1 (V2C_1165_13),
	.V2C_2 (V2C_1165_14),
	.V (V_1165)
);

VNU_2 #(quan_width) VNU1166 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_1166),
	.C2V_2 (C2V_15_1166),
	.L (L[17489:17475]),
	.V2C_1 (V2C_1166_14),
	.V2C_2 (V2C_1166_15),
	.V (V_1166)
);

VNU_2 #(quan_width) VNU1167 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_1167),
	.C2V_2 (C2V_16_1167),
	.L (L[17504:17490]),
	.V2C_1 (V2C_1167_15),
	.V2C_2 (V2C_1167_16),
	.V (V_1167)
);

VNU_2 #(quan_width) VNU1168 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_1168),
	.C2V_2 (C2V_17_1168),
	.L (L[17519:17505]),
	.V2C_1 (V2C_1168_16),
	.V2C_2 (V2C_1168_17),
	.V (V_1168)
);

VNU_2 #(quan_width) VNU1169 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_1169),
	.C2V_2 (C2V_18_1169),
	.L (L[17534:17520]),
	.V2C_1 (V2C_1169_17),
	.V2C_2 (V2C_1169_18),
	.V (V_1169)
);

VNU_2 #(quan_width) VNU1170 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_1170),
	.C2V_2 (C2V_19_1170),
	.L (L[17549:17535]),
	.V2C_1 (V2C_1170_18),
	.V2C_2 (V2C_1170_19),
	.V (V_1170)
);

VNU_2 #(quan_width) VNU1171 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_1171),
	.C2V_2 (C2V_20_1171),
	.L (L[17564:17550]),
	.V2C_1 (V2C_1171_19),
	.V2C_2 (V2C_1171_20),
	.V (V_1171)
);

VNU_2 #(quan_width) VNU1172 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_1172),
	.C2V_2 (C2V_21_1172),
	.L (L[17579:17565]),
	.V2C_1 (V2C_1172_20),
	.V2C_2 (V2C_1172_21),
	.V (V_1172)
);

VNU_2 #(quan_width) VNU1173 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_1173),
	.C2V_2 (C2V_22_1173),
	.L (L[17594:17580]),
	.V2C_1 (V2C_1173_21),
	.V2C_2 (V2C_1173_22),
	.V (V_1173)
);

VNU_2 #(quan_width) VNU1174 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_1174),
	.C2V_2 (C2V_23_1174),
	.L (L[17609:17595]),
	.V2C_1 (V2C_1174_22),
	.V2C_2 (V2C_1174_23),
	.V (V_1174)
);

VNU_2 #(quan_width) VNU1175 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_1175),
	.C2V_2 (C2V_24_1175),
	.L (L[17624:17610]),
	.V2C_1 (V2C_1175_23),
	.V2C_2 (V2C_1175_24),
	.V (V_1175)
);

VNU_2 #(quan_width) VNU1176 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_1176),
	.C2V_2 (C2V_25_1176),
	.L (L[17639:17625]),
	.V2C_1 (V2C_1176_24),
	.V2C_2 (V2C_1176_25),
	.V (V_1176)
);

VNU_2 #(quan_width) VNU1177 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_1177),
	.C2V_2 (C2V_26_1177),
	.L (L[17654:17640]),
	.V2C_1 (V2C_1177_25),
	.V2C_2 (V2C_1177_26),
	.V (V_1177)
);

VNU_2 #(quan_width) VNU1178 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_1178),
	.C2V_2 (C2V_27_1178),
	.L (L[17669:17655]),
	.V2C_1 (V2C_1178_26),
	.V2C_2 (V2C_1178_27),
	.V (V_1178)
);

VNU_2 #(quan_width) VNU1179 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_1179),
	.C2V_2 (C2V_28_1179),
	.L (L[17684:17670]),
	.V2C_1 (V2C_1179_27),
	.V2C_2 (V2C_1179_28),
	.V (V_1179)
);

VNU_2 #(quan_width) VNU1180 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_1180),
	.C2V_2 (C2V_29_1180),
	.L (L[17699:17685]),
	.V2C_1 (V2C_1180_28),
	.V2C_2 (V2C_1180_29),
	.V (V_1180)
);

VNU_2 #(quan_width) VNU1181 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_1181),
	.C2V_2 (C2V_30_1181),
	.L (L[17714:17700]),
	.V2C_1 (V2C_1181_29),
	.V2C_2 (V2C_1181_30),
	.V (V_1181)
);

VNU_2 #(quan_width) VNU1182 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_1182),
	.C2V_2 (C2V_31_1182),
	.L (L[17729:17715]),
	.V2C_1 (V2C_1182_30),
	.V2C_2 (V2C_1182_31),
	.V (V_1182)
);

VNU_2 #(quan_width) VNU1183 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_1183),
	.C2V_2 (C2V_32_1183),
	.L (L[17744:17730]),
	.V2C_1 (V2C_1183_31),
	.V2C_2 (V2C_1183_32),
	.V (V_1183)
);

VNU_2 #(quan_width) VNU1184 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_1184),
	.C2V_2 (C2V_33_1184),
	.L (L[17759:17745]),
	.V2C_1 (V2C_1184_32),
	.V2C_2 (V2C_1184_33),
	.V (V_1184)
);

VNU_2 #(quan_width) VNU1185 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_1185),
	.C2V_2 (C2V_34_1185),
	.L (L[17774:17760]),
	.V2C_1 (V2C_1185_33),
	.V2C_2 (V2C_1185_34),
	.V (V_1185)
);

VNU_2 #(quan_width) VNU1186 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_1186),
	.C2V_2 (C2V_35_1186),
	.L (L[17789:17775]),
	.V2C_1 (V2C_1186_34),
	.V2C_2 (V2C_1186_35),
	.V (V_1186)
);

VNU_2 #(quan_width) VNU1187 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_1187),
	.C2V_2 (C2V_36_1187),
	.L (L[17804:17790]),
	.V2C_1 (V2C_1187_35),
	.V2C_2 (V2C_1187_36),
	.V (V_1187)
);

VNU_2 #(quan_width) VNU1188 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_1188),
	.C2V_2 (C2V_37_1188),
	.L (L[17819:17805]),
	.V2C_1 (V2C_1188_36),
	.V2C_2 (V2C_1188_37),
	.V (V_1188)
);

VNU_2 #(quan_width) VNU1189 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_1189),
	.C2V_2 (C2V_38_1189),
	.L (L[17834:17820]),
	.V2C_1 (V2C_1189_37),
	.V2C_2 (V2C_1189_38),
	.V (V_1189)
);

VNU_2 #(quan_width) VNU1190 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_1190),
	.C2V_2 (C2V_39_1190),
	.L (L[17849:17835]),
	.V2C_1 (V2C_1190_38),
	.V2C_2 (V2C_1190_39),
	.V (V_1190)
);

VNU_2 #(quan_width) VNU1191 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_1191),
	.C2V_2 (C2V_40_1191),
	.L (L[17864:17850]),
	.V2C_1 (V2C_1191_39),
	.V2C_2 (V2C_1191_40),
	.V (V_1191)
);

VNU_2 #(quan_width) VNU1192 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_1192),
	.C2V_2 (C2V_41_1192),
	.L (L[17879:17865]),
	.V2C_1 (V2C_1192_40),
	.V2C_2 (V2C_1192_41),
	.V (V_1192)
);

VNU_2 #(quan_width) VNU1193 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_1193),
	.C2V_2 (C2V_42_1193),
	.L (L[17894:17880]),
	.V2C_1 (V2C_1193_41),
	.V2C_2 (V2C_1193_42),
	.V (V_1193)
);

VNU_2 #(quan_width) VNU1194 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_1194),
	.C2V_2 (C2V_43_1194),
	.L (L[17909:17895]),
	.V2C_1 (V2C_1194_42),
	.V2C_2 (V2C_1194_43),
	.V (V_1194)
);

VNU_2 #(quan_width) VNU1195 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_1195),
	.C2V_2 (C2V_44_1195),
	.L (L[17924:17910]),
	.V2C_1 (V2C_1195_43),
	.V2C_2 (V2C_1195_44),
	.V (V_1195)
);

VNU_2 #(quan_width) VNU1196 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_1196),
	.C2V_2 (C2V_45_1196),
	.L (L[17939:17925]),
	.V2C_1 (V2C_1196_44),
	.V2C_2 (V2C_1196_45),
	.V (V_1196)
);

VNU_2 #(quan_width) VNU1197 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_1197),
	.C2V_2 (C2V_46_1197),
	.L (L[17954:17940]),
	.V2C_1 (V2C_1197_45),
	.V2C_2 (V2C_1197_46),
	.V (V_1197)
);

VNU_2 #(quan_width) VNU1198 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_1198),
	.C2V_2 (C2V_47_1198),
	.L (L[17969:17955]),
	.V2C_1 (V2C_1198_46),
	.V2C_2 (V2C_1198_47),
	.V (V_1198)
);

VNU_2 #(quan_width) VNU1199 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_1199),
	.C2V_2 (C2V_48_1199),
	.L (L[17984:17970]),
	.V2C_1 (V2C_1199_47),
	.V2C_2 (V2C_1199_48),
	.V (V_1199)
);

VNU_2 #(quan_width) VNU1200 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_1200),
	.C2V_2 (C2V_49_1200),
	.L (L[17999:17985]),
	.V2C_1 (V2C_1200_48),
	.V2C_2 (V2C_1200_49),
	.V (V_1200)
);

VNU_2 #(quan_width) VNU1201 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_1201),
	.C2V_2 (C2V_50_1201),
	.L (L[18014:18000]),
	.V2C_1 (V2C_1201_49),
	.V2C_2 (V2C_1201_50),
	.V (V_1201)
);

VNU_2 #(quan_width) VNU1202 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_1202),
	.C2V_2 (C2V_51_1202),
	.L (L[18029:18015]),
	.V2C_1 (V2C_1202_50),
	.V2C_2 (V2C_1202_51),
	.V (V_1202)
);

VNU_2 #(quan_width) VNU1203 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_1203),
	.C2V_2 (C2V_52_1203),
	.L (L[18044:18030]),
	.V2C_1 (V2C_1203_51),
	.V2C_2 (V2C_1203_52),
	.V (V_1203)
);

VNU_2 #(quan_width) VNU1204 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_1204),
	.C2V_2 (C2V_53_1204),
	.L (L[18059:18045]),
	.V2C_1 (V2C_1204_52),
	.V2C_2 (V2C_1204_53),
	.V (V_1204)
);

VNU_2 #(quan_width) VNU1205 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_1205),
	.C2V_2 (C2V_54_1205),
	.L (L[18074:18060]),
	.V2C_1 (V2C_1205_53),
	.V2C_2 (V2C_1205_54),
	.V (V_1205)
);

VNU_2 #(quan_width) VNU1206 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_54_1206),
	.C2V_2 (C2V_55_1206),
	.L (L[18089:18075]),
	.V2C_1 (V2C_1206_54),
	.V2C_2 (V2C_1206_55),
	.V (V_1206)
);

VNU_2 #(quan_width) VNU1207 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_1207),
	.C2V_2 (C2V_56_1207),
	.L (L[18104:18090]),
	.V2C_1 (V2C_1207_55),
	.V2C_2 (V2C_1207_56),
	.V (V_1207)
);

VNU_2 #(quan_width) VNU1208 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_1208),
	.C2V_2 (C2V_57_1208),
	.L (L[18119:18105]),
	.V2C_1 (V2C_1208_56),
	.V2C_2 (V2C_1208_57),
	.V (V_1208)
);

VNU_2 #(quan_width) VNU1209 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_1209),
	.C2V_2 (C2V_58_1209),
	.L (L[18134:18120]),
	.V2C_1 (V2C_1209_57),
	.V2C_2 (V2C_1209_58),
	.V (V_1209)
);

VNU_2 #(quan_width) VNU1210 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_1210),
	.C2V_2 (C2V_59_1210),
	.L (L[18149:18135]),
	.V2C_1 (V2C_1210_58),
	.V2C_2 (V2C_1210_59),
	.V (V_1210)
);

VNU_2 #(quan_width) VNU1211 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_59_1211),
	.C2V_2 (C2V_60_1211),
	.L (L[18164:18150]),
	.V2C_1 (V2C_1211_59),
	.V2C_2 (V2C_1211_60),
	.V (V_1211)
);

VNU_2 #(quan_width) VNU1212 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_60_1212),
	.C2V_2 (C2V_61_1212),
	.L (L[18179:18165]),
	.V2C_1 (V2C_1212_60),
	.V2C_2 (V2C_1212_61),
	.V (V_1212)
);

VNU_2 #(quan_width) VNU1213 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_1213),
	.C2V_2 (C2V_62_1213),
	.L (L[18194:18180]),
	.V2C_1 (V2C_1213_61),
	.V2C_2 (V2C_1213_62),
	.V (V_1213)
);

VNU_2 #(quan_width) VNU1214 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_1214),
	.C2V_2 (C2V_63_1214),
	.L (L[18209:18195]),
	.V2C_1 (V2C_1214_62),
	.V2C_2 (V2C_1214_63),
	.V (V_1214)
);

VNU_2 #(quan_width) VNU1215 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_1215),
	.C2V_2 (C2V_64_1215),
	.L (L[18224:18210]),
	.V2C_1 (V2C_1215_63),
	.V2C_2 (V2C_1215_64),
	.V (V_1215)
);

VNU_2 #(quan_width) VNU1216 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_1216),
	.C2V_2 (C2V_65_1216),
	.L (L[18239:18225]),
	.V2C_1 (V2C_1216_64),
	.V2C_2 (V2C_1216_65),
	.V (V_1216)
);

VNU_2 #(quan_width) VNU1217 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_65_1217),
	.C2V_2 (C2V_66_1217),
	.L (L[18254:18240]),
	.V2C_1 (V2C_1217_65),
	.V2C_2 (V2C_1217_66),
	.V (V_1217)
);

VNU_2 #(quan_width) VNU1218 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_66_1218),
	.C2V_2 (C2V_67_1218),
	.L (L[18269:18255]),
	.V2C_1 (V2C_1218_66),
	.V2C_2 (V2C_1218_67),
	.V (V_1218)
);

VNU_2 #(quan_width) VNU1219 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_1219),
	.C2V_2 (C2V_68_1219),
	.L (L[18284:18270]),
	.V2C_1 (V2C_1219_67),
	.V2C_2 (V2C_1219_68),
	.V (V_1219)
);

VNU_2 #(quan_width) VNU1220 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_1220),
	.C2V_2 (C2V_69_1220),
	.L (L[18299:18285]),
	.V2C_1 (V2C_1220_68),
	.V2C_2 (V2C_1220_69),
	.V (V_1220)
);

VNU_2 #(quan_width) VNU1221 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_1221),
	.C2V_2 (C2V_70_1221),
	.L (L[18314:18300]),
	.V2C_1 (V2C_1221_69),
	.V2C_2 (V2C_1221_70),
	.V (V_1221)
);

VNU_2 #(quan_width) VNU1222 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_1222),
	.C2V_2 (C2V_71_1222),
	.L (L[18329:18315]),
	.V2C_1 (V2C_1222_70),
	.V2C_2 (V2C_1222_71),
	.V (V_1222)
);

VNU_2 #(quan_width) VNU1223 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_71_1223),
	.C2V_2 (C2V_72_1223),
	.L (L[18344:18330]),
	.V2C_1 (V2C_1223_71),
	.V2C_2 (V2C_1223_72),
	.V (V_1223)
);

VNU_2 #(quan_width) VNU1224 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_72_1224),
	.C2V_2 (C2V_73_1224),
	.L (L[18359:18345]),
	.V2C_1 (V2C_1224_72),
	.V2C_2 (V2C_1224_73),
	.V (V_1224)
);

VNU_2 #(quan_width) VNU1225 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_1225),
	.C2V_2 (C2V_74_1225),
	.L (L[18374:18360]),
	.V2C_1 (V2C_1225_73),
	.V2C_2 (V2C_1225_74),
	.V (V_1225)
);

VNU_2 #(quan_width) VNU1226 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_1226),
	.C2V_2 (C2V_75_1226),
	.L (L[18389:18375]),
	.V2C_1 (V2C_1226_74),
	.V2C_2 (V2C_1226_75),
	.V (V_1226)
);

VNU_2 #(quan_width) VNU1227 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_1227),
	.C2V_2 (C2V_76_1227),
	.L (L[18404:18390]),
	.V2C_1 (V2C_1227_75),
	.V2C_2 (V2C_1227_76),
	.V (V_1227)
);

VNU_2 #(quan_width) VNU1228 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_1228),
	.C2V_2 (C2V_77_1228),
	.L (L[18419:18405]),
	.V2C_1 (V2C_1228_76),
	.V2C_2 (V2C_1228_77),
	.V (V_1228)
);

VNU_2 #(quan_width) VNU1229 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_77_1229),
	.C2V_2 (C2V_78_1229),
	.L (L[18434:18420]),
	.V2C_1 (V2C_1229_77),
	.V2C_2 (V2C_1229_78),
	.V (V_1229)
);

VNU_2 #(quan_width) VNU1230 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_78_1230),
	.C2V_2 (C2V_79_1230),
	.L (L[18449:18435]),
	.V2C_1 (V2C_1230_78),
	.V2C_2 (V2C_1230_79),
	.V (V_1230)
);

VNU_2 #(quan_width) VNU1231 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_1231),
	.C2V_2 (C2V_80_1231),
	.L (L[18464:18450]),
	.V2C_1 (V2C_1231_79),
	.V2C_2 (V2C_1231_80),
	.V (V_1231)
);

VNU_2 #(quan_width) VNU1232 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_80_1232),
	.C2V_2 (C2V_81_1232),
	.L (L[18479:18465]),
	.V2C_1 (V2C_1232_80),
	.V2C_2 (V2C_1232_81),
	.V (V_1232)
);

VNU_2 #(quan_width) VNU1233 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_1233),
	.C2V_2 (C2V_82_1233),
	.L (L[18494:18480]),
	.V2C_1 (V2C_1233_81),
	.V2C_2 (V2C_1233_82),
	.V (V_1233)
);

VNU_2 #(quan_width) VNU1234 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_1234),
	.C2V_2 (C2V_83_1234),
	.L (L[18509:18495]),
	.V2C_1 (V2C_1234_82),
	.V2C_2 (V2C_1234_83),
	.V (V_1234)
);

VNU_2 #(quan_width) VNU1235 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_83_1235),
	.C2V_2 (C2V_84_1235),
	.L (L[18524:18510]),
	.V2C_1 (V2C_1235_83),
	.V2C_2 (V2C_1235_84),
	.V (V_1235)
);

VNU_2 #(quan_width) VNU1236 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_84_1236),
	.C2V_2 (C2V_85_1236),
	.L (L[18539:18525]),
	.V2C_1 (V2C_1236_84),
	.V2C_2 (V2C_1236_85),
	.V (V_1236)
);

VNU_2 #(quan_width) VNU1237 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_1237),
	.C2V_2 (C2V_86_1237),
	.L (L[18554:18540]),
	.V2C_1 (V2C_1237_85),
	.V2C_2 (V2C_1237_86),
	.V (V_1237)
);

VNU_2 #(quan_width) VNU1238 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_86_1238),
	.C2V_2 (C2V_87_1238),
	.L (L[18569:18555]),
	.V2C_1 (V2C_1238_86),
	.V2C_2 (V2C_1238_87),
	.V (V_1238)
);

VNU_2 #(quan_width) VNU1239 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_1239),
	.C2V_2 (C2V_88_1239),
	.L (L[18584:18570]),
	.V2C_1 (V2C_1239_87),
	.V2C_2 (V2C_1239_88),
	.V (V_1239)
);

VNU_2 #(quan_width) VNU1240 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_1240),
	.C2V_2 (C2V_89_1240),
	.L (L[18599:18585]),
	.V2C_1 (V2C_1240_88),
	.V2C_2 (V2C_1240_89),
	.V (V_1240)
);

VNU_2 #(quan_width) VNU1241 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_89_1241),
	.C2V_2 (C2V_90_1241),
	.L (L[18614:18600]),
	.V2C_1 (V2C_1241_89),
	.V2C_2 (V2C_1241_90),
	.V (V_1241)
);

VNU_2 #(quan_width) VNU1242 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_90_1242),
	.C2V_2 (C2V_91_1242),
	.L (L[18629:18615]),
	.V2C_1 (V2C_1242_90),
	.V2C_2 (V2C_1242_91),
	.V (V_1242)
);

VNU_2 #(quan_width) VNU1243 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_91_1243),
	.C2V_2 (C2V_92_1243),
	.L (L[18644:18630]),
	.V2C_1 (V2C_1243_91),
	.V2C_2 (V2C_1243_92),
	.V (V_1243)
);

VNU_2 #(quan_width) VNU1244 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_92_1244),
	.C2V_2 (C2V_93_1244),
	.L (L[18659:18645]),
	.V2C_1 (V2C_1244_92),
	.V2C_2 (V2C_1244_93),
	.V (V_1244)
);

VNU_2 #(quan_width) VNU1245 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_93_1245),
	.C2V_2 (C2V_94_1245),
	.L (L[18674:18660]),
	.V2C_1 (V2C_1245_93),
	.V2C_2 (V2C_1245_94),
	.V (V_1245)
);

VNU_2 #(quan_width) VNU1246 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_1246),
	.C2V_2 (C2V_95_1246),
	.L (L[18689:18675]),
	.V2C_1 (V2C_1246_94),
	.V2C_2 (V2C_1246_95),
	.V (V_1246)
);

VNU_2 #(quan_width) VNU1247 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_95_1247),
	.C2V_2 (C2V_96_1247),
	.L (L[18704:18690]),
	.V2C_1 (V2C_1247_95),
	.V2C_2 (V2C_1247_96),
	.V (V_1247)
);

VNU_2 #(quan_width) VNU1248 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_96_1248),
	.C2V_2 (C2V_97_1248),
	.L (L[18719:18705]),
	.V2C_1 (V2C_1248_96),
	.V2C_2 (V2C_1248_97),
	.V (V_1248)
);

VNU_2 #(quan_width) VNU1249 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_97_1249),
	.C2V_2 (C2V_98_1249),
	.L (L[18734:18720]),
	.V2C_1 (V2C_1249_97),
	.V2C_2 (V2C_1249_98),
	.V (V_1249)
);

VNU_2 #(quan_width) VNU1250 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_98_1250),
	.C2V_2 (C2V_99_1250),
	.L (L[18749:18735]),
	.V2C_1 (V2C_1250_98),
	.V2C_2 (V2C_1250_99),
	.V (V_1250)
);

VNU_2 #(quan_width) VNU1251 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_99_1251),
	.C2V_2 (C2V_100_1251),
	.L (L[18764:18750]),
	.V2C_1 (V2C_1251_99),
	.V2C_2 (V2C_1251_100),
	.V (V_1251)
);

VNU_2 #(quan_width) VNU1252 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_1252),
	.C2V_2 (C2V_101_1252),
	.L (L[18779:18765]),
	.V2C_1 (V2C_1252_100),
	.V2C_2 (V2C_1252_101),
	.V (V_1252)
);

VNU_2 #(quan_width) VNU1253 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_101_1253),
	.C2V_2 (C2V_102_1253),
	.L (L[18794:18780]),
	.V2C_1 (V2C_1253_101),
	.V2C_2 (V2C_1253_102),
	.V (V_1253)
);

VNU_2 #(quan_width) VNU1254 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_102_1254),
	.C2V_2 (C2V_103_1254),
	.L (L[18809:18795]),
	.V2C_1 (V2C_1254_102),
	.V2C_2 (V2C_1254_103),
	.V (V_1254)
);

VNU_2 #(quan_width) VNU1255 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_103_1255),
	.C2V_2 (C2V_104_1255),
	.L (L[18824:18810]),
	.V2C_1 (V2C_1255_103),
	.V2C_2 (V2C_1255_104),
	.V (V_1255)
);

VNU_2 #(quan_width) VNU1256 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_104_1256),
	.C2V_2 (C2V_105_1256),
	.L (L[18839:18825]),
	.V2C_1 (V2C_1256_104),
	.V2C_2 (V2C_1256_105),
	.V (V_1256)
);

VNU_2 #(quan_width) VNU1257 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_105_1257),
	.C2V_2 (C2V_106_1257),
	.L (L[18854:18840]),
	.V2C_1 (V2C_1257_105),
	.V2C_2 (V2C_1257_106),
	.V (V_1257)
);

VNU_2 #(quan_width) VNU1258 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_1258),
	.C2V_2 (C2V_107_1258),
	.L (L[18869:18855]),
	.V2C_1 (V2C_1258_106),
	.V2C_2 (V2C_1258_107),
	.V (V_1258)
);

VNU_2 #(quan_width) VNU1259 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_107_1259),
	.C2V_2 (C2V_108_1259),
	.L (L[18884:18870]),
	.V2C_1 (V2C_1259_107),
	.V2C_2 (V2C_1259_108),
	.V (V_1259)
);

VNU_2 #(quan_width) VNU1260 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_108_1260),
	.C2V_2 (C2V_109_1260),
	.L (L[18899:18885]),
	.V2C_1 (V2C_1260_108),
	.V2C_2 (V2C_1260_109),
	.V (V_1260)
);

VNU_2 #(quan_width) VNU1261 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_109_1261),
	.C2V_2 (C2V_110_1261),
	.L (L[18914:18900]),
	.V2C_1 (V2C_1261_109),
	.V2C_2 (V2C_1261_110),
	.V (V_1261)
);

VNU_2 #(quan_width) VNU1262 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_110_1262),
	.C2V_2 (C2V_111_1262),
	.L (L[18929:18915]),
	.V2C_1 (V2C_1262_110),
	.V2C_2 (V2C_1262_111),
	.V (V_1262)
);

VNU_2 #(quan_width) VNU1263 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_111_1263),
	.C2V_2 (C2V_112_1263),
	.L (L[18944:18930]),
	.V2C_1 (V2C_1263_111),
	.V2C_2 (V2C_1263_112),
	.V (V_1263)
);

VNU_2 #(quan_width) VNU1264 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_1264),
	.C2V_2 (C2V_113_1264),
	.L (L[18959:18945]),
	.V2C_1 (V2C_1264_112),
	.V2C_2 (V2C_1264_113),
	.V (V_1264)
);

VNU_2 #(quan_width) VNU1265 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_113_1265),
	.C2V_2 (C2V_114_1265),
	.L (L[18974:18960]),
	.V2C_1 (V2C_1265_113),
	.V2C_2 (V2C_1265_114),
	.V (V_1265)
);

VNU_2 #(quan_width) VNU1266 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_114_1266),
	.C2V_2 (C2V_115_1266),
	.L (L[18989:18975]),
	.V2C_1 (V2C_1266_114),
	.V2C_2 (V2C_1266_115),
	.V (V_1266)
);

VNU_2 #(quan_width) VNU1267 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_115_1267),
	.C2V_2 (C2V_116_1267),
	.L (L[19004:18990]),
	.V2C_1 (V2C_1267_115),
	.V2C_2 (V2C_1267_116),
	.V (V_1267)
);

VNU_2 #(quan_width) VNU1268 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_116_1268),
	.C2V_2 (C2V_117_1268),
	.L (L[19019:19005]),
	.V2C_1 (V2C_1268_116),
	.V2C_2 (V2C_1268_117),
	.V (V_1268)
);

VNU_2 #(quan_width) VNU1269 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_117_1269),
	.C2V_2 (C2V_118_1269),
	.L (L[19034:19020]),
	.V2C_1 (V2C_1269_117),
	.V2C_2 (V2C_1269_118),
	.V (V_1269)
);

VNU_2 #(quan_width) VNU1270 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_118_1270),
	.C2V_2 (C2V_119_1270),
	.L (L[19049:19035]),
	.V2C_1 (V2C_1270_118),
	.V2C_2 (V2C_1270_119),
	.V (V_1270)
);

VNU_2 #(quan_width) VNU1271 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_119_1271),
	.C2V_2 (C2V_120_1271),
	.L (L[19064:19050]),
	.V2C_1 (V2C_1271_119),
	.V2C_2 (V2C_1271_120),
	.V (V_1271)
);

VNU_2 #(quan_width) VNU1272 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_120_1272),
	.C2V_2 (C2V_121_1272),
	.L (L[19079:19065]),
	.V2C_1 (V2C_1272_120),
	.V2C_2 (V2C_1272_121),
	.V (V_1272)
);

VNU_2 #(quan_width) VNU1273 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_121_1273),
	.C2V_2 (C2V_122_1273),
	.L (L[19094:19080]),
	.V2C_1 (V2C_1273_121),
	.V2C_2 (V2C_1273_122),
	.V (V_1273)
);

VNU_2 #(quan_width) VNU1274 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_122_1274),
	.C2V_2 (C2V_123_1274),
	.L (L[19109:19095]),
	.V2C_1 (V2C_1274_122),
	.V2C_2 (V2C_1274_123),
	.V (V_1274)
);

VNU_2 #(quan_width) VNU1275 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_123_1275),
	.C2V_2 (C2V_124_1275),
	.L (L[19124:19110]),
	.V2C_1 (V2C_1275_123),
	.V2C_2 (V2C_1275_124),
	.V (V_1275)
);

VNU_2 #(quan_width) VNU1276 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_124_1276),
	.C2V_2 (C2V_125_1276),
	.L (L[19139:19125]),
	.V2C_1 (V2C_1276_124),
	.V2C_2 (V2C_1276_125),
	.V (V_1276)
);

VNU_2 #(quan_width) VNU1277 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_125_1277),
	.C2V_2 (C2V_126_1277),
	.L (L[19154:19140]),
	.V2C_1 (V2C_1277_125),
	.V2C_2 (V2C_1277_126),
	.V (V_1277)
);

VNU_2 #(quan_width) VNU1278 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_126_1278),
	.C2V_2 (C2V_127_1278),
	.L (L[19169:19155]),
	.V2C_1 (V2C_1278_126),
	.V2C_2 (V2C_1278_127),
	.V (V_1278)
);

VNU_2 #(quan_width) VNU1279 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_127_1279),
	.C2V_2 (C2V_128_1279),
	.L (L[19184:19170]),
	.V2C_1 (V2C_1279_127),
	.V2C_2 (V2C_1279_128),
	.V (V_1279)
);

VNU_2 #(quan_width) VNU1280 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_128_1280),
	.C2V_2 (C2V_129_1280),
	.L (L[19199:19185]),
	.V2C_1 (V2C_1280_128),
	.V2C_2 (V2C_1280_129),
	.V (V_1280)
);

VNU_2 #(quan_width) VNU1281 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_129_1281),
	.C2V_2 (C2V_130_1281),
	.L (L[19214:19200]),
	.V2C_1 (V2C_1281_129),
	.V2C_2 (V2C_1281_130),
	.V (V_1281)
);

VNU_2 #(quan_width) VNU1282 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_130_1282),
	.C2V_2 (C2V_131_1282),
	.L (L[19229:19215]),
	.V2C_1 (V2C_1282_130),
	.V2C_2 (V2C_1282_131),
	.V (V_1282)
);

VNU_2 #(quan_width) VNU1283 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_131_1283),
	.C2V_2 (C2V_132_1283),
	.L (L[19244:19230]),
	.V2C_1 (V2C_1283_131),
	.V2C_2 (V2C_1283_132),
	.V (V_1283)
);

VNU_2 #(quan_width) VNU1284 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_132_1284),
	.C2V_2 (C2V_133_1284),
	.L (L[19259:19245]),
	.V2C_1 (V2C_1284_132),
	.V2C_2 (V2C_1284_133),
	.V (V_1284)
);

VNU_2 #(quan_width) VNU1285 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_133_1285),
	.C2V_2 (C2V_134_1285),
	.L (L[19274:19260]),
	.V2C_1 (V2C_1285_133),
	.V2C_2 (V2C_1285_134),
	.V (V_1285)
);

VNU_2 #(quan_width) VNU1286 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_134_1286),
	.C2V_2 (C2V_135_1286),
	.L (L[19289:19275]),
	.V2C_1 (V2C_1286_134),
	.V2C_2 (V2C_1286_135),
	.V (V_1286)
);

VNU_2 #(quan_width) VNU1287 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_135_1287),
	.C2V_2 (C2V_136_1287),
	.L (L[19304:19290]),
	.V2C_1 (V2C_1287_135),
	.V2C_2 (V2C_1287_136),
	.V (V_1287)
);

VNU_2 #(quan_width) VNU1288 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_136_1288),
	.C2V_2 (C2V_137_1288),
	.L (L[19319:19305]),
	.V2C_1 (V2C_1288_136),
	.V2C_2 (V2C_1288_137),
	.V (V_1288)
);

VNU_2 #(quan_width) VNU1289 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_137_1289),
	.C2V_2 (C2V_138_1289),
	.L (L[19334:19320]),
	.V2C_1 (V2C_1289_137),
	.V2C_2 (V2C_1289_138),
	.V (V_1289)
);

VNU_2 #(quan_width) VNU1290 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_138_1290),
	.C2V_2 (C2V_139_1290),
	.L (L[19349:19335]),
	.V2C_1 (V2C_1290_138),
	.V2C_2 (V2C_1290_139),
	.V (V_1290)
);

VNU_2 #(quan_width) VNU1291 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_139_1291),
	.C2V_2 (C2V_140_1291),
	.L (L[19364:19350]),
	.V2C_1 (V2C_1291_139),
	.V2C_2 (V2C_1291_140),
	.V (V_1291)
);

VNU_2 #(quan_width) VNU1292 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_140_1292),
	.C2V_2 (C2V_141_1292),
	.L (L[19379:19365]),
	.V2C_1 (V2C_1292_140),
	.V2C_2 (V2C_1292_141),
	.V (V_1292)
);

VNU_2 #(quan_width) VNU1293 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_141_1293),
	.C2V_2 (C2V_142_1293),
	.L (L[19394:19380]),
	.V2C_1 (V2C_1293_141),
	.V2C_2 (V2C_1293_142),
	.V (V_1293)
);

VNU_2 #(quan_width) VNU1294 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_142_1294),
	.C2V_2 (C2V_143_1294),
	.L (L[19409:19395]),
	.V2C_1 (V2C_1294_142),
	.V2C_2 (V2C_1294_143),
	.V (V_1294)
);

VNU_2 #(quan_width) VNU1295 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_143_1295),
	.C2V_2 (C2V_144_1295),
	.L (L[19424:19410]),
	.V2C_1 (V2C_1295_143),
	.V2C_2 (V2C_1295_144),
	.V (V_1295)
);

VNU_2 #(quan_width) VNU1296 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_144_1296),
	.C2V_2 (C2V_145_1296),
	.L (L[19439:19425]),
	.V2C_1 (V2C_1296_144),
	.V2C_2 (V2C_1296_145),
	.V (V_1296)
);

VNU_2 #(quan_width) VNU1297 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_145_1297),
	.C2V_2 (C2V_146_1297),
	.L (L[19454:19440]),
	.V2C_1 (V2C_1297_145),
	.V2C_2 (V2C_1297_146),
	.V (V_1297)
);

VNU_2 #(quan_width) VNU1298 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_146_1298),
	.C2V_2 (C2V_147_1298),
	.L (L[19469:19455]),
	.V2C_1 (V2C_1298_146),
	.V2C_2 (V2C_1298_147),
	.V (V_1298)
);

VNU_2 #(quan_width) VNU1299 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_147_1299),
	.C2V_2 (C2V_148_1299),
	.L (L[19484:19470]),
	.V2C_1 (V2C_1299_147),
	.V2C_2 (V2C_1299_148),
	.V (V_1299)
);

VNU_2 #(quan_width) VNU1300 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_148_1300),
	.C2V_2 (C2V_149_1300),
	.L (L[19499:19485]),
	.V2C_1 (V2C_1300_148),
	.V2C_2 (V2C_1300_149),
	.V (V_1300)
);

VNU_2 #(quan_width) VNU1301 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_149_1301),
	.C2V_2 (C2V_150_1301),
	.L (L[19514:19500]),
	.V2C_1 (V2C_1301_149),
	.V2C_2 (V2C_1301_150),
	.V (V_1301)
);

VNU_2 #(quan_width) VNU1302 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_150_1302),
	.C2V_2 (C2V_151_1302),
	.L (L[19529:19515]),
	.V2C_1 (V2C_1302_150),
	.V2C_2 (V2C_1302_151),
	.V (V_1302)
);

VNU_2 #(quan_width) VNU1303 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_151_1303),
	.C2V_2 (C2V_152_1303),
	.L (L[19544:19530]),
	.V2C_1 (V2C_1303_151),
	.V2C_2 (V2C_1303_152),
	.V (V_1303)
);

VNU_2 #(quan_width) VNU1304 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_152_1304),
	.C2V_2 (C2V_153_1304),
	.L (L[19559:19545]),
	.V2C_1 (V2C_1304_152),
	.V2C_2 (V2C_1304_153),
	.V (V_1304)
);

VNU_2 #(quan_width) VNU1305 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_153_1305),
	.C2V_2 (C2V_154_1305),
	.L (L[19574:19560]),
	.V2C_1 (V2C_1305_153),
	.V2C_2 (V2C_1305_154),
	.V (V_1305)
);

VNU_2 #(quan_width) VNU1306 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_154_1306),
	.C2V_2 (C2V_155_1306),
	.L (L[19589:19575]),
	.V2C_1 (V2C_1306_154),
	.V2C_2 (V2C_1306_155),
	.V (V_1306)
);

VNU_2 #(quan_width) VNU1307 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_155_1307),
	.C2V_2 (C2V_156_1307),
	.L (L[19604:19590]),
	.V2C_1 (V2C_1307_155),
	.V2C_2 (V2C_1307_156),
	.V (V_1307)
);

VNU_2 #(quan_width) VNU1308 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_156_1308),
	.C2V_2 (C2V_157_1308),
	.L (L[19619:19605]),
	.V2C_1 (V2C_1308_156),
	.V2C_2 (V2C_1308_157),
	.V (V_1308)
);

VNU_2 #(quan_width) VNU1309 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_157_1309),
	.C2V_2 (C2V_158_1309),
	.L (L[19634:19620]),
	.V2C_1 (V2C_1309_157),
	.V2C_2 (V2C_1309_158),
	.V (V_1309)
);

VNU_2 #(quan_width) VNU1310 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_158_1310),
	.C2V_2 (C2V_159_1310),
	.L (L[19649:19635]),
	.V2C_1 (V2C_1310_158),
	.V2C_2 (V2C_1310_159),
	.V (V_1310)
);

VNU_2 #(quan_width) VNU1311 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_159_1311),
	.C2V_2 (C2V_160_1311),
	.L (L[19664:19650]),
	.V2C_1 (V2C_1311_159),
	.V2C_2 (V2C_1311_160),
	.V (V_1311)
);

VNU_2 #(quan_width) VNU1312 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_160_1312),
	.C2V_2 (C2V_161_1312),
	.L (L[19679:19665]),
	.V2C_1 (V2C_1312_160),
	.V2C_2 (V2C_1312_161),
	.V (V_1312)
);

VNU_2 #(quan_width) VNU1313 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_161_1313),
	.C2V_2 (C2V_162_1313),
	.L (L[19694:19680]),
	.V2C_1 (V2C_1313_161),
	.V2C_2 (V2C_1313_162),
	.V (V_1313)
);

VNU_2 #(quan_width) VNU1314 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_162_1314),
	.C2V_2 (C2V_163_1314),
	.L (L[19709:19695]),
	.V2C_1 (V2C_1314_162),
	.V2C_2 (V2C_1314_163),
	.V (V_1314)
);

VNU_2 #(quan_width) VNU1315 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_163_1315),
	.C2V_2 (C2V_164_1315),
	.L (L[19724:19710]),
	.V2C_1 (V2C_1315_163),
	.V2C_2 (V2C_1315_164),
	.V (V_1315)
);

VNU_2 #(quan_width) VNU1316 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_164_1316),
	.C2V_2 (C2V_165_1316),
	.L (L[19739:19725]),
	.V2C_1 (V2C_1316_164),
	.V2C_2 (V2C_1316_165),
	.V (V_1316)
);

VNU_2 #(quan_width) VNU1317 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_165_1317),
	.C2V_2 (C2V_166_1317),
	.L (L[19754:19740]),
	.V2C_1 (V2C_1317_165),
	.V2C_2 (V2C_1317_166),
	.V (V_1317)
);

VNU_2 #(quan_width) VNU1318 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_166_1318),
	.C2V_2 (C2V_167_1318),
	.L (L[19769:19755]),
	.V2C_1 (V2C_1318_166),
	.V2C_2 (V2C_1318_167),
	.V (V_1318)
);

VNU_2 #(quan_width) VNU1319 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_167_1319),
	.C2V_2 (C2V_168_1319),
	.L (L[19784:19770]),
	.V2C_1 (V2C_1319_167),
	.V2C_2 (V2C_1319_168),
	.V (V_1319)
);

VNU_2 #(quan_width) VNU1320 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_168_1320),
	.C2V_2 (C2V_169_1320),
	.L (L[19799:19785]),
	.V2C_1 (V2C_1320_168),
	.V2C_2 (V2C_1320_169),
	.V (V_1320)
);

VNU_2 #(quan_width) VNU1321 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_169_1321),
	.C2V_2 (C2V_170_1321),
	.L (L[19814:19800]),
	.V2C_1 (V2C_1321_169),
	.V2C_2 (V2C_1321_170),
	.V (V_1321)
);

VNU_2 #(quan_width) VNU1322 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_170_1322),
	.C2V_2 (C2V_171_1322),
	.L (L[19829:19815]),
	.V2C_1 (V2C_1322_170),
	.V2C_2 (V2C_1322_171),
	.V (V_1322)
);

VNU_2 #(quan_width) VNU1323 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_171_1323),
	.C2V_2 (C2V_172_1323),
	.L (L[19844:19830]),
	.V2C_1 (V2C_1323_171),
	.V2C_2 (V2C_1323_172),
	.V (V_1323)
);

VNU_2 #(quan_width) VNU1324 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_172_1324),
	.C2V_2 (C2V_173_1324),
	.L (L[19859:19845]),
	.V2C_1 (V2C_1324_172),
	.V2C_2 (V2C_1324_173),
	.V (V_1324)
);

VNU_2 #(quan_width) VNU1325 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_173_1325),
	.C2V_2 (C2V_174_1325),
	.L (L[19874:19860]),
	.V2C_1 (V2C_1325_173),
	.V2C_2 (V2C_1325_174),
	.V (V_1325)
);

VNU_2 #(quan_width) VNU1326 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_174_1326),
	.C2V_2 (C2V_175_1326),
	.L (L[19889:19875]),
	.V2C_1 (V2C_1326_174),
	.V2C_2 (V2C_1326_175),
	.V (V_1326)
);

VNU_2 #(quan_width) VNU1327 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_175_1327),
	.C2V_2 (C2V_176_1327),
	.L (L[19904:19890]),
	.V2C_1 (V2C_1327_175),
	.V2C_2 (V2C_1327_176),
	.V (V_1327)
);

VNU_2 #(quan_width) VNU1328 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_176_1328),
	.C2V_2 (C2V_177_1328),
	.L (L[19919:19905]),
	.V2C_1 (V2C_1328_176),
	.V2C_2 (V2C_1328_177),
	.V (V_1328)
);

VNU_2 #(quan_width) VNU1329 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_177_1329),
	.C2V_2 (C2V_178_1329),
	.L (L[19934:19920]),
	.V2C_1 (V2C_1329_177),
	.V2C_2 (V2C_1329_178),
	.V (V_1329)
);

VNU_2 #(quan_width) VNU1330 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_178_1330),
	.C2V_2 (C2V_179_1330),
	.L (L[19949:19935]),
	.V2C_1 (V2C_1330_178),
	.V2C_2 (V2C_1330_179),
	.V (V_1330)
);

VNU_2 #(quan_width) VNU1331 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_179_1331),
	.C2V_2 (C2V_180_1331),
	.L (L[19964:19950]),
	.V2C_1 (V2C_1331_179),
	.V2C_2 (V2C_1331_180),
	.V (V_1331)
);

VNU_2 #(quan_width) VNU1332 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_180_1332),
	.C2V_2 (C2V_181_1332),
	.L (L[19979:19965]),
	.V2C_1 (V2C_1332_180),
	.V2C_2 (V2C_1332_181),
	.V (V_1332)
);

VNU_2 #(quan_width) VNU1333 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_181_1333),
	.C2V_2 (C2V_182_1333),
	.L (L[19994:19980]),
	.V2C_1 (V2C_1333_181),
	.V2C_2 (V2C_1333_182),
	.V (V_1333)
);

VNU_2 #(quan_width) VNU1334 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_182_1334),
	.C2V_2 (C2V_183_1334),
	.L (L[20009:19995]),
	.V2C_1 (V2C_1334_182),
	.V2C_2 (V2C_1334_183),
	.V (V_1334)
);

VNU_2 #(quan_width) VNU1335 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_183_1335),
	.C2V_2 (C2V_184_1335),
	.L (L[20024:20010]),
	.V2C_1 (V2C_1335_183),
	.V2C_2 (V2C_1335_184),
	.V (V_1335)
);

VNU_2 #(quan_width) VNU1336 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_184_1336),
	.C2V_2 (C2V_185_1336),
	.L (L[20039:20025]),
	.V2C_1 (V2C_1336_184),
	.V2C_2 (V2C_1336_185),
	.V (V_1336)
);

VNU_2 #(quan_width) VNU1337 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_185_1337),
	.C2V_2 (C2V_186_1337),
	.L (L[20054:20040]),
	.V2C_1 (V2C_1337_185),
	.V2C_2 (V2C_1337_186),
	.V (V_1337)
);

VNU_2 #(quan_width) VNU1338 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_186_1338),
	.C2V_2 (C2V_187_1338),
	.L (L[20069:20055]),
	.V2C_1 (V2C_1338_186),
	.V2C_2 (V2C_1338_187),
	.V (V_1338)
);

VNU_2 #(quan_width) VNU1339 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_187_1339),
	.C2V_2 (C2V_188_1339),
	.L (L[20084:20070]),
	.V2C_1 (V2C_1339_187),
	.V2C_2 (V2C_1339_188),
	.V (V_1339)
);

VNU_2 #(quan_width) VNU1340 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_188_1340),
	.C2V_2 (C2V_189_1340),
	.L (L[20099:20085]),
	.V2C_1 (V2C_1340_188),
	.V2C_2 (V2C_1340_189),
	.V (V_1340)
);

VNU_2 #(quan_width) VNU1341 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_189_1341),
	.C2V_2 (C2V_190_1341),
	.L (L[20114:20100]),
	.V2C_1 (V2C_1341_189),
	.V2C_2 (V2C_1341_190),
	.V (V_1341)
);

VNU_2 #(quan_width) VNU1342 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_190_1342),
	.C2V_2 (C2V_191_1342),
	.L (L[20129:20115]),
	.V2C_1 (V2C_1342_190),
	.V2C_2 (V2C_1342_191),
	.V (V_1342)
);

VNU_2 #(quan_width) VNU1343 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_191_1343),
	.C2V_2 (C2V_192_1343),
	.L (L[20144:20130]),
	.V2C_1 (V2C_1343_191),
	.V2C_2 (V2C_1343_192),
	.V (V_1343)
);

VNU_2 #(quan_width) VNU1344 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_192_1344),
	.C2V_2 (C2V_193_1344),
	.L (L[20159:20145]),
	.V2C_1 (V2C_1344_192),
	.V2C_2 (V2C_1344_193),
	.V (V_1344)
);

VNU_2 #(quan_width) VNU1345 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_193_1345),
	.C2V_2 (C2V_194_1345),
	.L (L[20174:20160]),
	.V2C_1 (V2C_1345_193),
	.V2C_2 (V2C_1345_194),
	.V (V_1345)
);

VNU_2 #(quan_width) VNU1346 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_194_1346),
	.C2V_2 (C2V_195_1346),
	.L (L[20189:20175]),
	.V2C_1 (V2C_1346_194),
	.V2C_2 (V2C_1346_195),
	.V (V_1346)
);

VNU_2 #(quan_width) VNU1347 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_195_1347),
	.C2V_2 (C2V_196_1347),
	.L (L[20204:20190]),
	.V2C_1 (V2C_1347_195),
	.V2C_2 (V2C_1347_196),
	.V (V_1347)
);

VNU_2 #(quan_width) VNU1348 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_196_1348),
	.C2V_2 (C2V_197_1348),
	.L (L[20219:20205]),
	.V2C_1 (V2C_1348_196),
	.V2C_2 (V2C_1348_197),
	.V (V_1348)
);

VNU_2 #(quan_width) VNU1349 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_197_1349),
	.C2V_2 (C2V_198_1349),
	.L (L[20234:20220]),
	.V2C_1 (V2C_1349_197),
	.V2C_2 (V2C_1349_198),
	.V (V_1349)
);

VNU_2 #(quan_width) VNU1350 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_198_1350),
	.C2V_2 (C2V_199_1350),
	.L (L[20249:20235]),
	.V2C_1 (V2C_1350_198),
	.V2C_2 (V2C_1350_199),
	.V (V_1350)
);

VNU_2 #(quan_width) VNU1351 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_199_1351),
	.C2V_2 (C2V_200_1351),
	.L (L[20264:20250]),
	.V2C_1 (V2C_1351_199),
	.V2C_2 (V2C_1351_200),
	.V (V_1351)
);

VNU_2 #(quan_width) VNU1352 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_200_1352),
	.C2V_2 (C2V_201_1352),
	.L (L[20279:20265]),
	.V2C_1 (V2C_1352_200),
	.V2C_2 (V2C_1352_201),
	.V (V_1352)
);

VNU_2 #(quan_width) VNU1353 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_201_1353),
	.C2V_2 (C2V_202_1353),
	.L (L[20294:20280]),
	.V2C_1 (V2C_1353_201),
	.V2C_2 (V2C_1353_202),
	.V (V_1353)
);

VNU_2 #(quan_width) VNU1354 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_202_1354),
	.C2V_2 (C2V_203_1354),
	.L (L[20309:20295]),
	.V2C_1 (V2C_1354_202),
	.V2C_2 (V2C_1354_203),
	.V (V_1354)
);

VNU_2 #(quan_width) VNU1355 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_203_1355),
	.C2V_2 (C2V_204_1355),
	.L (L[20324:20310]),
	.V2C_1 (V2C_1355_203),
	.V2C_2 (V2C_1355_204),
	.V (V_1355)
);

VNU_2 #(quan_width) VNU1356 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_204_1356),
	.C2V_2 (C2V_205_1356),
	.L (L[20339:20325]),
	.V2C_1 (V2C_1356_204),
	.V2C_2 (V2C_1356_205),
	.V (V_1356)
);

VNU_2 #(quan_width) VNU1357 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_205_1357),
	.C2V_2 (C2V_206_1357),
	.L (L[20354:20340]),
	.V2C_1 (V2C_1357_205),
	.V2C_2 (V2C_1357_206),
	.V (V_1357)
);

VNU_2 #(quan_width) VNU1358 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_206_1358),
	.C2V_2 (C2V_207_1358),
	.L (L[20369:20355]),
	.V2C_1 (V2C_1358_206),
	.V2C_2 (V2C_1358_207),
	.V (V_1358)
);

VNU_2 #(quan_width) VNU1359 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_207_1359),
	.C2V_2 (C2V_208_1359),
	.L (L[20384:20370]),
	.V2C_1 (V2C_1359_207),
	.V2C_2 (V2C_1359_208),
	.V (V_1359)
);

VNU_2 #(quan_width) VNU1360 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_208_1360),
	.C2V_2 (C2V_209_1360),
	.L (L[20399:20385]),
	.V2C_1 (V2C_1360_208),
	.V2C_2 (V2C_1360_209),
	.V (V_1360)
);

VNU_2 #(quan_width) VNU1361 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_209_1361),
	.C2V_2 (C2V_210_1361),
	.L (L[20414:20400]),
	.V2C_1 (V2C_1361_209),
	.V2C_2 (V2C_1361_210),
	.V (V_1361)
);

VNU_2 #(quan_width) VNU1362 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_210_1362),
	.C2V_2 (C2V_211_1362),
	.L (L[20429:20415]),
	.V2C_1 (V2C_1362_210),
	.V2C_2 (V2C_1362_211),
	.V (V_1362)
);

VNU_2 #(quan_width) VNU1363 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_211_1363),
	.C2V_2 (C2V_212_1363),
	.L (L[20444:20430]),
	.V2C_1 (V2C_1363_211),
	.V2C_2 (V2C_1363_212),
	.V (V_1363)
);

VNU_2 #(quan_width) VNU1364 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_212_1364),
	.C2V_2 (C2V_213_1364),
	.L (L[20459:20445]),
	.V2C_1 (V2C_1364_212),
	.V2C_2 (V2C_1364_213),
	.V (V_1364)
);

VNU_2 #(quan_width) VNU1365 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_213_1365),
	.C2V_2 (C2V_214_1365),
	.L (L[20474:20460]),
	.V2C_1 (V2C_1365_213),
	.V2C_2 (V2C_1365_214),
	.V (V_1365)
);

VNU_2 #(quan_width) VNU1366 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_214_1366),
	.C2V_2 (C2V_215_1366),
	.L (L[20489:20475]),
	.V2C_1 (V2C_1366_214),
	.V2C_2 (V2C_1366_215),
	.V (V_1366)
);

VNU_2 #(quan_width) VNU1367 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_215_1367),
	.C2V_2 (C2V_216_1367),
	.L (L[20504:20490]),
	.V2C_1 (V2C_1367_215),
	.V2C_2 (V2C_1367_216),
	.V (V_1367)
);

VNU_2 #(quan_width) VNU1368 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_216_1368),
	.C2V_2 (C2V_217_1368),
	.L (L[20519:20505]),
	.V2C_1 (V2C_1368_216),
	.V2C_2 (V2C_1368_217),
	.V (V_1368)
);

VNU_2 #(quan_width) VNU1369 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_217_1369),
	.C2V_2 (C2V_218_1369),
	.L (L[20534:20520]),
	.V2C_1 (V2C_1369_217),
	.V2C_2 (V2C_1369_218),
	.V (V_1369)
);

VNU_2 #(quan_width) VNU1370 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_218_1370),
	.C2V_2 (C2V_219_1370),
	.L (L[20549:20535]),
	.V2C_1 (V2C_1370_218),
	.V2C_2 (V2C_1370_219),
	.V (V_1370)
);

VNU_2 #(quan_width) VNU1371 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_219_1371),
	.C2V_2 (C2V_220_1371),
	.L (L[20564:20550]),
	.V2C_1 (V2C_1371_219),
	.V2C_2 (V2C_1371_220),
	.V (V_1371)
);

VNU_2 #(quan_width) VNU1372 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_220_1372),
	.C2V_2 (C2V_221_1372),
	.L (L[20579:20565]),
	.V2C_1 (V2C_1372_220),
	.V2C_2 (V2C_1372_221),
	.V (V_1372)
);

VNU_2 #(quan_width) VNU1373 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_221_1373),
	.C2V_2 (C2V_222_1373),
	.L (L[20594:20580]),
	.V2C_1 (V2C_1373_221),
	.V2C_2 (V2C_1373_222),
	.V (V_1373)
);

VNU_2 #(quan_width) VNU1374 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_222_1374),
	.C2V_2 (C2V_223_1374),
	.L (L[20609:20595]),
	.V2C_1 (V2C_1374_222),
	.V2C_2 (V2C_1374_223),
	.V (V_1374)
);

VNU_2 #(quan_width) VNU1375 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_223_1375),
	.C2V_2 (C2V_224_1375),
	.L (L[20624:20610]),
	.V2C_1 (V2C_1375_223),
	.V2C_2 (V2C_1375_224),
	.V (V_1375)
);

VNU_2 #(quan_width) VNU1376 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_224_1376),
	.C2V_2 (C2V_225_1376),
	.L (L[20639:20625]),
	.V2C_1 (V2C_1376_224),
	.V2C_2 (V2C_1376_225),
	.V (V_1376)
);

VNU_2 #(quan_width) VNU1377 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_225_1377),
	.C2V_2 (C2V_226_1377),
	.L (L[20654:20640]),
	.V2C_1 (V2C_1377_225),
	.V2C_2 (V2C_1377_226),
	.V (V_1377)
);

VNU_2 #(quan_width) VNU1378 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_226_1378),
	.C2V_2 (C2V_227_1378),
	.L (L[20669:20655]),
	.V2C_1 (V2C_1378_226),
	.V2C_2 (V2C_1378_227),
	.V (V_1378)
);

VNU_2 #(quan_width) VNU1379 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_227_1379),
	.C2V_2 (C2V_228_1379),
	.L (L[20684:20670]),
	.V2C_1 (V2C_1379_227),
	.V2C_2 (V2C_1379_228),
	.V (V_1379)
);

VNU_2 #(quan_width) VNU1380 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_228_1380),
	.C2V_2 (C2V_229_1380),
	.L (L[20699:20685]),
	.V2C_1 (V2C_1380_228),
	.V2C_2 (V2C_1380_229),
	.V (V_1380)
);

VNU_2 #(quan_width) VNU1381 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_229_1381),
	.C2V_2 (C2V_230_1381),
	.L (L[20714:20700]),
	.V2C_1 (V2C_1381_229),
	.V2C_2 (V2C_1381_230),
	.V (V_1381)
);

VNU_2 #(quan_width) VNU1382 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_230_1382),
	.C2V_2 (C2V_231_1382),
	.L (L[20729:20715]),
	.V2C_1 (V2C_1382_230),
	.V2C_2 (V2C_1382_231),
	.V (V_1382)
);

VNU_2 #(quan_width) VNU1383 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_231_1383),
	.C2V_2 (C2V_232_1383),
	.L (L[20744:20730]),
	.V2C_1 (V2C_1383_231),
	.V2C_2 (V2C_1383_232),
	.V (V_1383)
);

VNU_2 #(quan_width) VNU1384 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_232_1384),
	.C2V_2 (C2V_233_1384),
	.L (L[20759:20745]),
	.V2C_1 (V2C_1384_232),
	.V2C_2 (V2C_1384_233),
	.V (V_1384)
);

VNU_2 #(quan_width) VNU1385 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_233_1385),
	.C2V_2 (C2V_234_1385),
	.L (L[20774:20760]),
	.V2C_1 (V2C_1385_233),
	.V2C_2 (V2C_1385_234),
	.V (V_1385)
);

VNU_2 #(quan_width) VNU1386 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_234_1386),
	.C2V_2 (C2V_235_1386),
	.L (L[20789:20775]),
	.V2C_1 (V2C_1386_234),
	.V2C_2 (V2C_1386_235),
	.V (V_1386)
);

VNU_2 #(quan_width) VNU1387 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_235_1387),
	.C2V_2 (C2V_236_1387),
	.L (L[20804:20790]),
	.V2C_1 (V2C_1387_235),
	.V2C_2 (V2C_1387_236),
	.V (V_1387)
);

VNU_2 #(quan_width) VNU1388 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_236_1388),
	.C2V_2 (C2V_237_1388),
	.L (L[20819:20805]),
	.V2C_1 (V2C_1388_236),
	.V2C_2 (V2C_1388_237),
	.V (V_1388)
);

VNU_2 #(quan_width) VNU1389 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_237_1389),
	.C2V_2 (C2V_238_1389),
	.L (L[20834:20820]),
	.V2C_1 (V2C_1389_237),
	.V2C_2 (V2C_1389_238),
	.V (V_1389)
);

VNU_2 #(quan_width) VNU1390 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_238_1390),
	.C2V_2 (C2V_239_1390),
	.L (L[20849:20835]),
	.V2C_1 (V2C_1390_238),
	.V2C_2 (V2C_1390_239),
	.V (V_1390)
);

VNU_2 #(quan_width) VNU1391 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_239_1391),
	.C2V_2 (C2V_240_1391),
	.L (L[20864:20850]),
	.V2C_1 (V2C_1391_239),
	.V2C_2 (V2C_1391_240),
	.V (V_1391)
);

VNU_2 #(quan_width) VNU1392 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_240_1392),
	.C2V_2 (C2V_241_1392),
	.L (L[20879:20865]),
	.V2C_1 (V2C_1392_240),
	.V2C_2 (V2C_1392_241),
	.V (V_1392)
);

VNU_2 #(quan_width) VNU1393 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_241_1393),
	.C2V_2 (C2V_242_1393),
	.L (L[20894:20880]),
	.V2C_1 (V2C_1393_241),
	.V2C_2 (V2C_1393_242),
	.V (V_1393)
);

VNU_2 #(quan_width) VNU1394 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_242_1394),
	.C2V_2 (C2V_243_1394),
	.L (L[20909:20895]),
	.V2C_1 (V2C_1394_242),
	.V2C_2 (V2C_1394_243),
	.V (V_1394)
);

VNU_2 #(quan_width) VNU1395 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_243_1395),
	.C2V_2 (C2V_244_1395),
	.L (L[20924:20910]),
	.V2C_1 (V2C_1395_243),
	.V2C_2 (V2C_1395_244),
	.V (V_1395)
);

VNU_2 #(quan_width) VNU1396 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_244_1396),
	.C2V_2 (C2V_245_1396),
	.L (L[20939:20925]),
	.V2C_1 (V2C_1396_244),
	.V2C_2 (V2C_1396_245),
	.V (V_1396)
);

VNU_2 #(quan_width) VNU1397 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_245_1397),
	.C2V_2 (C2V_246_1397),
	.L (L[20954:20940]),
	.V2C_1 (V2C_1397_245),
	.V2C_2 (V2C_1397_246),
	.V (V_1397)
);

VNU_2 #(quan_width) VNU1398 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_246_1398),
	.C2V_2 (C2V_247_1398),
	.L (L[20969:20955]),
	.V2C_1 (V2C_1398_246),
	.V2C_2 (V2C_1398_247),
	.V (V_1398)
);

VNU_2 #(quan_width) VNU1399 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_247_1399),
	.C2V_2 (C2V_248_1399),
	.L (L[20984:20970]),
	.V2C_1 (V2C_1399_247),
	.V2C_2 (V2C_1399_248),
	.V (V_1399)
);

VNU_2 #(quan_width) VNU1400 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_248_1400),
	.C2V_2 (C2V_249_1400),
	.L (L[20999:20985]),
	.V2C_1 (V2C_1400_248),
	.V2C_2 (V2C_1400_249),
	.V (V_1400)
);

VNU_2 #(quan_width) VNU1401 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_249_1401),
	.C2V_2 (C2V_250_1401),
	.L (L[21014:21000]),
	.V2C_1 (V2C_1401_249),
	.V2C_2 (V2C_1401_250),
	.V (V_1401)
);

VNU_2 #(quan_width) VNU1402 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_250_1402),
	.C2V_2 (C2V_251_1402),
	.L (L[21029:21015]),
	.V2C_1 (V2C_1402_250),
	.V2C_2 (V2C_1402_251),
	.V (V_1402)
);

VNU_2 #(quan_width) VNU1403 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_251_1403),
	.C2V_2 (C2V_252_1403),
	.L (L[21044:21030]),
	.V2C_1 (V2C_1403_251),
	.V2C_2 (V2C_1403_252),
	.V (V_1403)
);

VNU_2 #(quan_width) VNU1404 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_252_1404),
	.C2V_2 (C2V_253_1404),
	.L (L[21059:21045]),
	.V2C_1 (V2C_1404_252),
	.V2C_2 (V2C_1404_253),
	.V (V_1404)
);

VNU_2 #(quan_width) VNU1405 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_253_1405),
	.C2V_2 (C2V_254_1405),
	.L (L[21074:21060]),
	.V2C_1 (V2C_1405_253),
	.V2C_2 (V2C_1405_254),
	.V (V_1405)
);

VNU_2 #(quan_width) VNU1406 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_254_1406),
	.C2V_2 (C2V_255_1406),
	.L (L[21089:21075]),
	.V2C_1 (V2C_1406_254),
	.V2C_2 (V2C_1406_255),
	.V (V_1406)
);

VNU_2 #(quan_width) VNU1407 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_255_1407),
	.C2V_2 (C2V_256_1407),
	.L (L[21104:21090]),
	.V2C_1 (V2C_1407_255),
	.V2C_2 (V2C_1407_256),
	.V (V_1407)
);

VNU_2 #(quan_width) VNU1408 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_256_1408),
	.C2V_2 (C2V_257_1408),
	.L (L[21119:21105]),
	.V2C_1 (V2C_1408_256),
	.V2C_2 (V2C_1408_257),
	.V (V_1408)
);

VNU_2 #(quan_width) VNU1409 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_257_1409),
	.C2V_2 (C2V_258_1409),
	.L (L[21134:21120]),
	.V2C_1 (V2C_1409_257),
	.V2C_2 (V2C_1409_258),
	.V (V_1409)
);

VNU_2 #(quan_width) VNU1410 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_258_1410),
	.C2V_2 (C2V_259_1410),
	.L (L[21149:21135]),
	.V2C_1 (V2C_1410_258),
	.V2C_2 (V2C_1410_259),
	.V (V_1410)
);

VNU_2 #(quan_width) VNU1411 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_259_1411),
	.C2V_2 (C2V_260_1411),
	.L (L[21164:21150]),
	.V2C_1 (V2C_1411_259),
	.V2C_2 (V2C_1411_260),
	.V (V_1411)
);

VNU_2 #(quan_width) VNU1412 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_260_1412),
	.C2V_2 (C2V_261_1412),
	.L (L[21179:21165]),
	.V2C_1 (V2C_1412_260),
	.V2C_2 (V2C_1412_261),
	.V (V_1412)
);

VNU_2 #(quan_width) VNU1413 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_261_1413),
	.C2V_2 (C2V_262_1413),
	.L (L[21194:21180]),
	.V2C_1 (V2C_1413_261),
	.V2C_2 (V2C_1413_262),
	.V (V_1413)
);

VNU_2 #(quan_width) VNU1414 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_262_1414),
	.C2V_2 (C2V_263_1414),
	.L (L[21209:21195]),
	.V2C_1 (V2C_1414_262),
	.V2C_2 (V2C_1414_263),
	.V (V_1414)
);

VNU_2 #(quan_width) VNU1415 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_263_1415),
	.C2V_2 (C2V_264_1415),
	.L (L[21224:21210]),
	.V2C_1 (V2C_1415_263),
	.V2C_2 (V2C_1415_264),
	.V (V_1415)
);

VNU_2 #(quan_width) VNU1416 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_264_1416),
	.C2V_2 (C2V_265_1416),
	.L (L[21239:21225]),
	.V2C_1 (V2C_1416_264),
	.V2C_2 (V2C_1416_265),
	.V (V_1416)
);

VNU_2 #(quan_width) VNU1417 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_265_1417),
	.C2V_2 (C2V_266_1417),
	.L (L[21254:21240]),
	.V2C_1 (V2C_1417_265),
	.V2C_2 (V2C_1417_266),
	.V (V_1417)
);

VNU_2 #(quan_width) VNU1418 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_266_1418),
	.C2V_2 (C2V_267_1418),
	.L (L[21269:21255]),
	.V2C_1 (V2C_1418_266),
	.V2C_2 (V2C_1418_267),
	.V (V_1418)
);

VNU_2 #(quan_width) VNU1419 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_267_1419),
	.C2V_2 (C2V_268_1419),
	.L (L[21284:21270]),
	.V2C_1 (V2C_1419_267),
	.V2C_2 (V2C_1419_268),
	.V (V_1419)
);

VNU_2 #(quan_width) VNU1420 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_268_1420),
	.C2V_2 (C2V_269_1420),
	.L (L[21299:21285]),
	.V2C_1 (V2C_1420_268),
	.V2C_2 (V2C_1420_269),
	.V (V_1420)
);

VNU_2 #(quan_width) VNU1421 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_269_1421),
	.C2V_2 (C2V_270_1421),
	.L (L[21314:21300]),
	.V2C_1 (V2C_1421_269),
	.V2C_2 (V2C_1421_270),
	.V (V_1421)
);

VNU_2 #(quan_width) VNU1422 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_270_1422),
	.C2V_2 (C2V_271_1422),
	.L (L[21329:21315]),
	.V2C_1 (V2C_1422_270),
	.V2C_2 (V2C_1422_271),
	.V (V_1422)
);

VNU_2 #(quan_width) VNU1423 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_271_1423),
	.C2V_2 (C2V_272_1423),
	.L (L[21344:21330]),
	.V2C_1 (V2C_1423_271),
	.V2C_2 (V2C_1423_272),
	.V (V_1423)
);

VNU_2 #(quan_width) VNU1424 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_272_1424),
	.C2V_2 (C2V_273_1424),
	.L (L[21359:21345]),
	.V2C_1 (V2C_1424_272),
	.V2C_2 (V2C_1424_273),
	.V (V_1424)
);

VNU_2 #(quan_width) VNU1425 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_273_1425),
	.C2V_2 (C2V_274_1425),
	.L (L[21374:21360]),
	.V2C_1 (V2C_1425_273),
	.V2C_2 (V2C_1425_274),
	.V (V_1425)
);

VNU_2 #(quan_width) VNU1426 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_274_1426),
	.C2V_2 (C2V_275_1426),
	.L (L[21389:21375]),
	.V2C_1 (V2C_1426_274),
	.V2C_2 (V2C_1426_275),
	.V (V_1426)
);

VNU_2 #(quan_width) VNU1427 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_275_1427),
	.C2V_2 (C2V_276_1427),
	.L (L[21404:21390]),
	.V2C_1 (V2C_1427_275),
	.V2C_2 (V2C_1427_276),
	.V (V_1427)
);

VNU_2 #(quan_width) VNU1428 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_276_1428),
	.C2V_2 (C2V_277_1428),
	.L (L[21419:21405]),
	.V2C_1 (V2C_1428_276),
	.V2C_2 (V2C_1428_277),
	.V (V_1428)
);

VNU_2 #(quan_width) VNU1429 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_277_1429),
	.C2V_2 (C2V_278_1429),
	.L (L[21434:21420]),
	.V2C_1 (V2C_1429_277),
	.V2C_2 (V2C_1429_278),
	.V (V_1429)
);

VNU_2 #(quan_width) VNU1430 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_278_1430),
	.C2V_2 (C2V_279_1430),
	.L (L[21449:21435]),
	.V2C_1 (V2C_1430_278),
	.V2C_2 (V2C_1430_279),
	.V (V_1430)
);

VNU_2 #(quan_width) VNU1431 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_279_1431),
	.C2V_2 (C2V_280_1431),
	.L (L[21464:21450]),
	.V2C_1 (V2C_1431_279),
	.V2C_2 (V2C_1431_280),
	.V (V_1431)
);

VNU_2 #(quan_width) VNU1432 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_280_1432),
	.C2V_2 (C2V_281_1432),
	.L (L[21479:21465]),
	.V2C_1 (V2C_1432_280),
	.V2C_2 (V2C_1432_281),
	.V (V_1432)
);

VNU_2 #(quan_width) VNU1433 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_281_1433),
	.C2V_2 (C2V_282_1433),
	.L (L[21494:21480]),
	.V2C_1 (V2C_1433_281),
	.V2C_2 (V2C_1433_282),
	.V (V_1433)
);

VNU_2 #(quan_width) VNU1434 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_282_1434),
	.C2V_2 (C2V_283_1434),
	.L (L[21509:21495]),
	.V2C_1 (V2C_1434_282),
	.V2C_2 (V2C_1434_283),
	.V (V_1434)
);

VNU_2 #(quan_width) VNU1435 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_283_1435),
	.C2V_2 (C2V_284_1435),
	.L (L[21524:21510]),
	.V2C_1 (V2C_1435_283),
	.V2C_2 (V2C_1435_284),
	.V (V_1435)
);

VNU_2 #(quan_width) VNU1436 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_284_1436),
	.C2V_2 (C2V_285_1436),
	.L (L[21539:21525]),
	.V2C_1 (V2C_1436_284),
	.V2C_2 (V2C_1436_285),
	.V (V_1436)
);

VNU_2 #(quan_width) VNU1437 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_285_1437),
	.C2V_2 (C2V_286_1437),
	.L (L[21554:21540]),
	.V2C_1 (V2C_1437_285),
	.V2C_2 (V2C_1437_286),
	.V (V_1437)
);

VNU_2 #(quan_width) VNU1438 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_286_1438),
	.C2V_2 (C2V_287_1438),
	.L (L[21569:21555]),
	.V2C_1 (V2C_1438_286),
	.V2C_2 (V2C_1438_287),
	.V (V_1438)
);

VNU_2 #(quan_width) VNU1439 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_287_1439),
	.C2V_2 (C2V_288_1439),
	.L (L[21584:21570]),
	.V2C_1 (V2C_1439_287),
	.V2C_2 (V2C_1439_288),
	.V (V_1439)
);

VNU_1 #(quan_width) VNU1440 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_288_1440),
	.L (L[21599:21585]),
	.V2C_1 (V2C_1440_288),
	.V (V_1440)
);

endmodule