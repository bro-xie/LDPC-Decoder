module Decoder #(
	parameter code_length = 1440,
	parameter quan_width = 10
)
(
	input wire clk,
	input wire rst,
	input wire in_valid,
	input wire [15:0] in_index,
	input wire [4 * quan_width - 1: 0] data_in,
	output reg out_valid,
	output reg [15:0] out_index,
	output reg [4 - 1: 0] data_out
);

//wire [code_length - 1:0] Bit;
wire Bit_1, Bit_2, Bit_3, Bit_4, Bit_5, Bit_6, Bit_7, Bit_8, Bit_9, Bit_10, Bit_11, Bit_12, Bit_13, Bit_14, Bit_15, Bit_16, Bit_17, Bit_18, Bit_19, Bit_20, Bit_21, Bit_22, Bit_23, Bit_24, Bit_25, Bit_26, Bit_27, Bit_28, Bit_29, Bit_30, Bit_31, Bit_32, Bit_33, Bit_34, Bit_35, Bit_36, Bit_37, Bit_38, Bit_39, Bit_40, Bit_41, Bit_42, Bit_43, Bit_44, Bit_45, Bit_46, Bit_47, Bit_48, Bit_49, Bit_50, Bit_51, Bit_52, Bit_53, Bit_54, Bit_55, Bit_56, Bit_57, Bit_58, Bit_59, Bit_60, Bit_61, Bit_62, Bit_63, Bit_64, Bit_65, Bit_66, Bit_67, Bit_68, Bit_69, Bit_70, Bit_71, Bit_72, Bit_73, Bit_74, Bit_75, Bit_76, Bit_77, Bit_78, Bit_79, Bit_80, Bit_81, Bit_82, Bit_83, Bit_84, Bit_85, Bit_86, Bit_87, Bit_88, Bit_89, Bit_90, Bit_91, Bit_92, Bit_93, Bit_94, Bit_95, Bit_96, Bit_97, Bit_98, Bit_99, Bit_100, Bit_101, Bit_102, Bit_103, Bit_104, Bit_105, Bit_106, Bit_107, Bit_108, Bit_109, Bit_110, Bit_111, Bit_112, Bit_113, Bit_114, Bit_115, Bit_116, Bit_117, Bit_118, Bit_119, Bit_120, Bit_121, Bit_122, Bit_123, Bit_124, Bit_125, Bit_126, Bit_127, Bit_128, Bit_129, Bit_130, Bit_131, Bit_132, Bit_133, Bit_134, Bit_135, Bit_136, Bit_137, Bit_138, Bit_139, Bit_140, Bit_141, Bit_142, Bit_143, Bit_144, Bit_145, Bit_146, Bit_147, Bit_148, Bit_149, Bit_150, Bit_151, Bit_152, Bit_153, Bit_154, Bit_155, Bit_156, Bit_157, Bit_158, Bit_159, Bit_160, Bit_161, Bit_162, Bit_163, Bit_164, Bit_165, Bit_166, Bit_167, Bit_168, Bit_169, Bit_170, Bit_171, Bit_172, Bit_173, Bit_174, Bit_175, Bit_176, Bit_177, Bit_178, Bit_179, Bit_180, Bit_181, Bit_182, Bit_183, Bit_184, Bit_185, Bit_186, Bit_187, Bit_188, Bit_189, Bit_190, Bit_191, Bit_192, Bit_193, Bit_194, Bit_195, Bit_196, Bit_197, Bit_198, Bit_199, Bit_200, Bit_201, Bit_202, Bit_203, Bit_204, Bit_205, Bit_206, Bit_207, Bit_208, Bit_209, Bit_210, Bit_211, Bit_212, Bit_213, Bit_214, Bit_215, Bit_216, Bit_217, Bit_218, Bit_219, Bit_220, Bit_221, Bit_222, Bit_223, Bit_224, Bit_225, Bit_226, Bit_227, Bit_228, Bit_229, Bit_230, Bit_231, Bit_232, Bit_233, Bit_234, Bit_235, Bit_236, Bit_237, Bit_238, Bit_239, Bit_240, Bit_241, Bit_242, Bit_243, Bit_244, Bit_245, Bit_246, Bit_247, Bit_248, Bit_249, Bit_250, Bit_251, Bit_252, Bit_253, Bit_254, Bit_255, Bit_256, Bit_257, Bit_258, Bit_259, Bit_260, Bit_261, Bit_262, Bit_263, Bit_264, Bit_265, Bit_266, Bit_267, Bit_268, Bit_269, Bit_270, Bit_271, Bit_272, Bit_273, Bit_274, Bit_275, Bit_276, Bit_277, Bit_278, Bit_279, Bit_280, Bit_281, Bit_282, Bit_283, Bit_284, Bit_285, Bit_286, Bit_287, Bit_288, Bit_289, Bit_290, Bit_291, Bit_292, Bit_293, Bit_294, Bit_295, Bit_296, Bit_297, Bit_298, Bit_299, Bit_300, Bit_301, Bit_302, Bit_303, Bit_304, Bit_305, Bit_306, Bit_307, Bit_308, Bit_309, Bit_310, Bit_311, Bit_312, Bit_313, Bit_314, Bit_315, Bit_316, Bit_317, Bit_318, Bit_319, Bit_320, Bit_321, Bit_322, Bit_323, Bit_324, Bit_325, Bit_326, Bit_327, Bit_328, Bit_329, Bit_330, Bit_331, Bit_332, Bit_333, Bit_334, Bit_335, Bit_336, Bit_337, Bit_338, Bit_339, Bit_340, Bit_341, Bit_342, Bit_343, Bit_344, Bit_345, Bit_346, Bit_347, Bit_348, Bit_349, Bit_350, Bit_351, Bit_352, Bit_353, Bit_354, Bit_355, Bit_356, Bit_357, Bit_358, Bit_359, Bit_360, Bit_361, Bit_362, Bit_363, Bit_364, Bit_365, Bit_366, Bit_367, Bit_368, Bit_369, Bit_370, Bit_371, Bit_372, Bit_373, Bit_374, Bit_375, Bit_376, Bit_377, Bit_378, Bit_379, Bit_380, Bit_381, Bit_382, Bit_383, Bit_384, Bit_385, Bit_386, Bit_387, Bit_388, Bit_389, Bit_390, Bit_391, Bit_392, Bit_393, Bit_394, Bit_395, Bit_396, Bit_397, Bit_398, Bit_399, Bit_400, Bit_401, Bit_402, Bit_403, Bit_404, Bit_405, Bit_406, Bit_407, Bit_408, Bit_409, Bit_410, Bit_411, Bit_412, Bit_413, Bit_414, Bit_415, Bit_416, Bit_417, Bit_418, Bit_419, Bit_420, Bit_421, Bit_422, Bit_423, Bit_424, Bit_425, Bit_426, Bit_427, Bit_428, Bit_429, Bit_430, Bit_431, Bit_432, Bit_433, Bit_434, Bit_435, Bit_436, Bit_437, Bit_438, Bit_439, Bit_440, Bit_441, Bit_442, Bit_443, Bit_444, Bit_445, Bit_446, Bit_447, Bit_448, Bit_449, Bit_450, Bit_451, Bit_452, Bit_453, Bit_454, Bit_455, Bit_456, Bit_457, Bit_458, Bit_459, Bit_460, Bit_461, Bit_462, Bit_463, Bit_464, Bit_465, Bit_466, Bit_467, Bit_468, Bit_469, Bit_470, Bit_471, Bit_472, Bit_473, Bit_474, Bit_475, Bit_476, Bit_477, Bit_478, Bit_479, Bit_480, Bit_481, Bit_482, Bit_483, Bit_484, Bit_485, Bit_486, Bit_487, Bit_488, Bit_489, Bit_490, Bit_491, Bit_492, Bit_493, Bit_494, Bit_495, Bit_496, Bit_497, Bit_498, Bit_499, Bit_500, Bit_501, Bit_502, Bit_503, Bit_504, Bit_505, Bit_506, Bit_507, Bit_508, Bit_509, Bit_510, Bit_511, Bit_512, Bit_513, Bit_514, Bit_515, Bit_516, Bit_517, Bit_518, Bit_519, Bit_520, Bit_521, Bit_522, Bit_523, Bit_524, Bit_525, Bit_526, Bit_527, Bit_528, Bit_529, Bit_530, Bit_531, Bit_532, Bit_533, Bit_534, Bit_535, Bit_536, Bit_537, Bit_538, Bit_539, Bit_540, Bit_541, Bit_542, Bit_543, Bit_544, Bit_545, Bit_546, Bit_547, Bit_548, Bit_549, Bit_550, Bit_551, Bit_552, Bit_553, Bit_554, Bit_555, Bit_556, Bit_557, Bit_558, Bit_559, Bit_560, Bit_561, Bit_562, Bit_563, Bit_564, Bit_565, Bit_566, Bit_567, Bit_568, Bit_569, Bit_570, Bit_571, Bit_572, Bit_573, Bit_574, Bit_575, Bit_576, Bit_577, Bit_578, Bit_579, Bit_580, Bit_581, Bit_582, Bit_583, Bit_584, Bit_585, Bit_586, Bit_587, Bit_588, Bit_589, Bit_590, Bit_591, Bit_592, Bit_593, Bit_594, Bit_595, Bit_596, Bit_597, Bit_598, Bit_599, Bit_600, Bit_601, Bit_602, Bit_603, Bit_604, Bit_605, Bit_606, Bit_607, Bit_608, Bit_609, Bit_610, Bit_611, Bit_612, Bit_613, Bit_614, Bit_615, Bit_616, Bit_617, Bit_618, Bit_619, Bit_620, Bit_621, Bit_622, Bit_623, Bit_624, Bit_625, Bit_626, Bit_627, Bit_628, Bit_629, Bit_630, Bit_631, Bit_632, Bit_633, Bit_634, Bit_635, Bit_636, Bit_637, Bit_638, Bit_639, Bit_640, Bit_641, Bit_642, Bit_643, Bit_644, Bit_645, Bit_646, Bit_647, Bit_648, Bit_649, Bit_650, Bit_651, Bit_652, Bit_653, Bit_654, Bit_655, Bit_656, Bit_657, Bit_658, Bit_659, Bit_660, Bit_661, Bit_662, Bit_663, Bit_664, Bit_665, Bit_666, Bit_667, Bit_668, Bit_669, Bit_670, Bit_671, Bit_672, Bit_673, Bit_674, Bit_675, Bit_676, Bit_677, Bit_678, Bit_679, Bit_680, Bit_681, Bit_682, Bit_683, Bit_684, Bit_685, Bit_686, Bit_687, Bit_688, Bit_689, Bit_690, Bit_691, Bit_692, Bit_693, Bit_694, Bit_695, Bit_696, Bit_697, Bit_698, Bit_699, Bit_700, Bit_701, Bit_702, Bit_703, Bit_704, Bit_705, Bit_706, Bit_707, Bit_708, Bit_709, Bit_710, Bit_711, Bit_712, Bit_713, Bit_714, Bit_715, Bit_716, Bit_717, Bit_718, Bit_719, Bit_720, Bit_721, Bit_722, Bit_723, Bit_724, Bit_725, Bit_726, Bit_727, Bit_728, Bit_729, Bit_730, Bit_731, Bit_732, Bit_733, Bit_734, Bit_735, Bit_736, Bit_737, Bit_738, Bit_739, Bit_740, Bit_741, Bit_742, Bit_743, Bit_744, Bit_745, Bit_746, Bit_747, Bit_748, Bit_749, Bit_750, Bit_751, Bit_752, Bit_753, Bit_754, Bit_755, Bit_756, Bit_757, Bit_758, Bit_759, Bit_760, Bit_761, Bit_762, Bit_763, Bit_764, Bit_765, Bit_766, Bit_767, Bit_768, Bit_769, Bit_770, Bit_771, Bit_772, Bit_773, Bit_774, Bit_775, Bit_776, Bit_777, Bit_778, Bit_779, Bit_780, Bit_781, Bit_782, Bit_783, Bit_784, Bit_785, Bit_786, Bit_787, Bit_788, Bit_789, Bit_790, Bit_791, Bit_792, Bit_793, Bit_794, Bit_795, Bit_796, Bit_797, Bit_798, Bit_799, Bit_800, Bit_801, Bit_802, Bit_803, Bit_804, Bit_805, Bit_806, Bit_807, Bit_808, Bit_809, Bit_810, Bit_811, Bit_812, Bit_813, Bit_814, Bit_815, Bit_816, Bit_817, Bit_818, Bit_819, Bit_820, Bit_821, Bit_822, Bit_823, Bit_824, Bit_825, Bit_826, Bit_827, Bit_828, Bit_829, Bit_830, Bit_831, Bit_832, Bit_833, Bit_834, Bit_835, Bit_836, Bit_837, Bit_838, Bit_839, Bit_840, Bit_841, Bit_842, Bit_843, Bit_844, Bit_845, Bit_846, Bit_847, Bit_848, Bit_849, Bit_850, Bit_851, Bit_852, Bit_853, Bit_854, Bit_855, Bit_856, Bit_857, Bit_858, Bit_859, Bit_860, Bit_861, Bit_862, Bit_863, Bit_864, Bit_865, Bit_866, Bit_867, Bit_868, Bit_869, Bit_870, Bit_871, Bit_872, Bit_873, Bit_874, Bit_875, Bit_876, Bit_877, Bit_878, Bit_879, Bit_880, Bit_881, Bit_882, Bit_883, Bit_884, Bit_885, Bit_886, Bit_887, Bit_888, Bit_889, Bit_890, Bit_891, Bit_892, Bit_893, Bit_894, Bit_895, Bit_896, Bit_897, Bit_898, Bit_899, Bit_900, Bit_901, Bit_902, Bit_903, Bit_904, Bit_905, Bit_906, Bit_907, Bit_908, Bit_909, Bit_910, Bit_911, Bit_912, Bit_913, Bit_914, Bit_915, Bit_916, Bit_917, Bit_918, Bit_919, Bit_920, Bit_921, Bit_922, Bit_923, Bit_924, Bit_925, Bit_926, Bit_927, Bit_928, Bit_929, Bit_930, Bit_931, Bit_932, Bit_933, Bit_934, Bit_935, Bit_936, Bit_937, Bit_938, Bit_939, Bit_940, Bit_941, Bit_942, Bit_943, Bit_944, Bit_945, Bit_946, Bit_947, Bit_948, Bit_949, Bit_950, Bit_951, Bit_952, Bit_953, Bit_954, Bit_955, Bit_956, Bit_957, Bit_958, Bit_959, Bit_960, Bit_961, Bit_962, Bit_963, Bit_964, Bit_965, Bit_966, Bit_967, Bit_968, Bit_969, Bit_970, Bit_971, Bit_972, Bit_973, Bit_974, Bit_975, Bit_976, Bit_977, Bit_978, Bit_979, Bit_980, Bit_981, Bit_982, Bit_983, Bit_984, Bit_985, Bit_986, Bit_987, Bit_988, Bit_989, Bit_990, Bit_991, Bit_992, Bit_993, Bit_994, Bit_995, Bit_996, Bit_997, Bit_998, Bit_999, Bit_1000, Bit_1001, Bit_1002, Bit_1003, Bit_1004, Bit_1005, Bit_1006, Bit_1007, Bit_1008, Bit_1009, Bit_1010, Bit_1011, Bit_1012, Bit_1013, Bit_1014, Bit_1015, Bit_1016, Bit_1017, Bit_1018, Bit_1019, Bit_1020, Bit_1021, Bit_1022, Bit_1023, Bit_1024, Bit_1025, Bit_1026, Bit_1027, Bit_1028, Bit_1029, Bit_1030, Bit_1031, Bit_1032, Bit_1033, Bit_1034, Bit_1035, Bit_1036, Bit_1037, Bit_1038, Bit_1039, Bit_1040, Bit_1041, Bit_1042, Bit_1043, Bit_1044, Bit_1045, Bit_1046, Bit_1047, Bit_1048, Bit_1049, Bit_1050, Bit_1051, Bit_1052, Bit_1053, Bit_1054, Bit_1055, Bit_1056, Bit_1057, Bit_1058, Bit_1059, Bit_1060, Bit_1061, Bit_1062, Bit_1063, Bit_1064, Bit_1065, Bit_1066, Bit_1067, Bit_1068, Bit_1069, Bit_1070, Bit_1071, Bit_1072, Bit_1073, Bit_1074, Bit_1075, Bit_1076, Bit_1077, Bit_1078, Bit_1079, Bit_1080, Bit_1081, Bit_1082, Bit_1083, Bit_1084, Bit_1085, Bit_1086, Bit_1087, Bit_1088, Bit_1089, Bit_1090, Bit_1091, Bit_1092, Bit_1093, Bit_1094, Bit_1095, Bit_1096, Bit_1097, Bit_1098, Bit_1099, Bit_1100, Bit_1101, Bit_1102, Bit_1103, Bit_1104, Bit_1105, Bit_1106, Bit_1107, Bit_1108, Bit_1109, Bit_1110, Bit_1111, Bit_1112, Bit_1113, Bit_1114, Bit_1115, Bit_1116, Bit_1117, Bit_1118, Bit_1119, Bit_1120, Bit_1121, Bit_1122, Bit_1123, Bit_1124, Bit_1125, Bit_1126, Bit_1127, Bit_1128, Bit_1129, Bit_1130, Bit_1131, Bit_1132, Bit_1133, Bit_1134, Bit_1135, Bit_1136, Bit_1137, Bit_1138, Bit_1139, Bit_1140, Bit_1141, Bit_1142, Bit_1143, Bit_1144, Bit_1145, Bit_1146, Bit_1147, Bit_1148, Bit_1149, Bit_1150, Bit_1151, Bit_1152, Bit_1153, Bit_1154, Bit_1155, Bit_1156, Bit_1157, Bit_1158, Bit_1159, Bit_1160, Bit_1161, Bit_1162, Bit_1163, Bit_1164, Bit_1165, Bit_1166, Bit_1167, Bit_1168, Bit_1169, Bit_1170, Bit_1171, Bit_1172, Bit_1173, Bit_1174, Bit_1175, Bit_1176, Bit_1177, Bit_1178, Bit_1179, Bit_1180, Bit_1181, Bit_1182, Bit_1183, Bit_1184, Bit_1185, Bit_1186, Bit_1187, Bit_1188, Bit_1189, Bit_1190, Bit_1191, Bit_1192, Bit_1193, Bit_1194, Bit_1195, Bit_1196, Bit_1197, Bit_1198, Bit_1199, Bit_1200, Bit_1201, Bit_1202, Bit_1203, Bit_1204, Bit_1205, Bit_1206, Bit_1207, Bit_1208, Bit_1209, Bit_1210, Bit_1211, Bit_1212, Bit_1213, Bit_1214, Bit_1215, Bit_1216, Bit_1217, Bit_1218, Bit_1219, Bit_1220, Bit_1221, Bit_1222, Bit_1223, Bit_1224, Bit_1225, Bit_1226, Bit_1227, Bit_1228, Bit_1229, Bit_1230, Bit_1231, Bit_1232, Bit_1233, Bit_1234, Bit_1235, Bit_1236, Bit_1237, Bit_1238, Bit_1239, Bit_1240, Bit_1241, Bit_1242, Bit_1243, Bit_1244, Bit_1245, Bit_1246, Bit_1247, Bit_1248, Bit_1249, Bit_1250, Bit_1251, Bit_1252, Bit_1253, Bit_1254, Bit_1255, Bit_1256, Bit_1257, Bit_1258, Bit_1259, Bit_1260, Bit_1261, Bit_1262, Bit_1263, Bit_1264, Bit_1265, Bit_1266, Bit_1267, Bit_1268, Bit_1269, Bit_1270, Bit_1271, Bit_1272, Bit_1273, Bit_1274, Bit_1275, Bit_1276, Bit_1277, Bit_1278, Bit_1279, Bit_1280, Bit_1281, Bit_1282, Bit_1283, Bit_1284, Bit_1285, Bit_1286, Bit_1287, Bit_1288, Bit_1289, Bit_1290, Bit_1291, Bit_1292, Bit_1293, Bit_1294, Bit_1295, Bit_1296, Bit_1297, Bit_1298, Bit_1299, Bit_1300, Bit_1301, Bit_1302, Bit_1303, Bit_1304, Bit_1305, Bit_1306, Bit_1307, Bit_1308, Bit_1309, Bit_1310, Bit_1311, Bit_1312, Bit_1313, Bit_1314, Bit_1315, Bit_1316, Bit_1317, Bit_1318, Bit_1319, Bit_1320, Bit_1321, Bit_1322, Bit_1323, Bit_1324, Bit_1325, Bit_1326, Bit_1327, Bit_1328, Bit_1329, Bit_1330, Bit_1331, Bit_1332, Bit_1333, Bit_1334, Bit_1335, Bit_1336, Bit_1337, Bit_1338, Bit_1339, Bit_1340, Bit_1341, Bit_1342, Bit_1343, Bit_1344, Bit_1345, Bit_1346, Bit_1347, Bit_1348, Bit_1349, Bit_1350, Bit_1351, Bit_1352, Bit_1353, Bit_1354, Bit_1355, Bit_1356, Bit_1357, Bit_1358, Bit_1359, Bit_1360, Bit_1361, Bit_1362, Bit_1363, Bit_1364, Bit_1365, Bit_1366, Bit_1367, Bit_1368, Bit_1369, Bit_1370, Bit_1371, Bit_1372, Bit_1373, Bit_1374, Bit_1375, Bit_1376, Bit_1377, Bit_1378, Bit_1379, Bit_1380, Bit_1381, Bit_1382, Bit_1383, Bit_1384, Bit_1385, Bit_1386, Bit_1387, Bit_1388, Bit_1389, Bit_1390, Bit_1391, Bit_1392, Bit_1393, Bit_1394, Bit_1395, Bit_1396, Bit_1397, Bit_1398, Bit_1399, Bit_1400, Bit_1401, Bit_1402, Bit_1403, Bit_1404, Bit_1405, Bit_1406, Bit_1407, Bit_1408, Bit_1409, Bit_1410, Bit_1411, Bit_1412, Bit_1413, Bit_1414, Bit_1415, Bit_1416, Bit_1417, Bit_1418, Bit_1419, Bit_1420, Bit_1421, Bit_1422, Bit_1423, Bit_1424, Bit_1425, Bit_1426, Bit_1427, Bit_1428, Bit_1429, Bit_1430, Bit_1431, Bit_1432, Bit_1433, Bit_1434, Bit_1435, Bit_1436, Bit_1437, Bit_1438, Bit_1439, Bit_1440;
reg  [7:0] cnt;
reg  [4:0] iter;
reg  Check_1, Check_2, Check_3, Check_4, Check_5, Check_6, Check_7, Check_8, Check_9, Check_10, Check_11, Check_12, Check_13, Check_14, Check_15, Check_16, Check_17, Check_18, Check_19, Check_20, Check_21, Check_22, Check_23, Check_24, Check_25, Check_26, Check_27, Check_28, Check_29, Check_30, Check_31, Check_32, Check_33, Check_34, Check_35, Check_36, Check_37, Check_38, Check_39, Check_40, Check_41, Check_42, Check_43, Check_44, Check_45, Check_46, Check_47, Check_48, Check_49, Check_50, Check_51, Check_52, Check_53, Check_54, Check_55, Check_56, Check_57, Check_58, Check_59, Check_60, Check_61, Check_62, Check_63, Check_64, Check_65, Check_66, Check_67, Check_68, Check_69, Check_70, Check_71, Check_72, Check_73, Check_74, Check_75, Check_76, Check_77, Check_78, Check_79, Check_80, Check_81, Check_82, Check_83, Check_84, Check_85, Check_86, Check_87, Check_88, Check_89, Check_90, Check_91, Check_92, Check_93, Check_94, Check_95, Check_96, Check_97, Check_98, Check_99, Check_100, Check_101, Check_102, Check_103, Check_104, Check_105, Check_106, Check_107, Check_108, Check_109, Check_110, Check_111, Check_112, Check_113, Check_114, Check_115, Check_116, Check_117, Check_118, Check_119, Check_120, Check_121, Check_122, Check_123, Check_124, Check_125, Check_126, Check_127, Check_128, Check_129, Check_130, Check_131, Check_132, Check_133, Check_134, Check_135, Check_136, Check_137, Check_138, Check_139, Check_140, Check_141, Check_142, Check_143, Check_144, Check_145, Check_146, Check_147, Check_148, Check_149, Check_150, Check_151, Check_152, Check_153, Check_154, Check_155, Check_156, Check_157, Check_158, Check_159, Check_160, Check_161, Check_162, Check_163, Check_164, Check_165, Check_166, Check_167, Check_168, Check_169, Check_170, Check_171, Check_172, Check_173, Check_174, Check_175, Check_176, Check_177, Check_178, Check_179, Check_180, Check_181, Check_182, Check_183, Check_184, Check_185, Check_186, Check_187, Check_188, Check_189, Check_190, Check_191, Check_192, Check_193, Check_194, Check_195, Check_196, Check_197, Check_198, Check_199, Check_200, Check_201, Check_202, Check_203, Check_204, Check_205, Check_206, Check_207, Check_208, Check_209, Check_210, Check_211, Check_212, Check_213, Check_214, Check_215, Check_216, Check_217, Check_218, Check_219, Check_220, Check_221, Check_222, Check_223, Check_224, Check_225, Check_226, Check_227, Check_228, Check_229, Check_230, Check_231, Check_232, Check_233, Check_234, Check_235, Check_236, Check_237, Check_238, Check_239, Check_240, Check_241, Check_242, Check_243, Check_244, Check_245, Check_246, Check_247, Check_248, Check_249, Check_250, Check_251, Check_252, Check_253, Check_254, Check_255, Check_256, Check_257, Check_258, Check_259, Check_260, Check_261, Check_262, Check_263, Check_264, Check_265, Check_266, Check_267, Check_268, Check_269, Check_270, Check_271, Check_272, Check_273, Check_274, Check_275, Check_276, Check_277, Check_278, Check_279, Check_280, Check_281, Check_282, Check_283, Check_284, Check_285, Check_286, Check_287, Check_288, Check_Sum;
reg  [quan_width - 1:0] L_1, L_2, L_3, L_4, L_5, L_6, L_7, L_8, L_9, L_10, L_11, L_12, L_13, L_14, L_15, L_16, L_17, L_18, L_19, L_20, L_21, L_22, L_23, L_24, L_25, L_26, L_27, L_28, L_29, L_30, L_31, L_32, L_33, L_34, L_35, L_36, L_37, L_38, L_39, L_40, L_41, L_42, L_43, L_44, L_45, L_46, L_47, L_48, L_49, L_50, L_51, L_52, L_53, L_54, L_55, L_56, L_57, L_58, L_59, L_60, L_61, L_62, L_63, L_64, L_65, L_66, L_67, L_68, L_69, L_70, L_71, L_72, L_73, L_74, L_75, L_76, L_77, L_78, L_79, L_80, L_81, L_82, L_83, L_84, L_85, L_86, L_87, L_88, L_89, L_90, L_91, L_92, L_93, L_94, L_95, L_96, L_97, L_98, L_99, L_100, L_101, L_102, L_103, L_104, L_105, L_106, L_107, L_108, L_109, L_110, L_111, L_112, L_113, L_114, L_115, L_116, L_117, L_118, L_119, L_120, L_121, L_122, L_123, L_124, L_125, L_126, L_127, L_128, L_129, L_130, L_131, L_132, L_133, L_134, L_135, L_136, L_137, L_138, L_139, L_140, L_141, L_142, L_143, L_144, L_145, L_146, L_147, L_148, L_149, L_150, L_151, L_152, L_153, L_154, L_155, L_156, L_157, L_158, L_159, L_160, L_161, L_162, L_163, L_164, L_165, L_166, L_167, L_168, L_169, L_170, L_171, L_172, L_173, L_174, L_175, L_176, L_177, L_178, L_179, L_180, L_181, L_182, L_183, L_184, L_185, L_186, L_187, L_188, L_189, L_190, L_191, L_192, L_193, L_194, L_195, L_196, L_197, L_198, L_199, L_200, L_201, L_202, L_203, L_204, L_205, L_206, L_207, L_208, L_209, L_210, L_211, L_212, L_213, L_214, L_215, L_216, L_217, L_218, L_219, L_220, L_221, L_222, L_223, L_224, L_225, L_226, L_227, L_228, L_229, L_230, L_231, L_232, L_233, L_234, L_235, L_236, L_237, L_238, L_239, L_240, L_241, L_242, L_243, L_244, L_245, L_246, L_247, L_248, L_249, L_250, L_251, L_252, L_253, L_254, L_255, L_256, L_257, L_258, L_259, L_260, L_261, L_262, L_263, L_264, L_265, L_266, L_267, L_268, L_269, L_270, L_271, L_272, L_273, L_274, L_275, L_276, L_277, L_278, L_279, L_280, L_281, L_282, L_283, L_284, L_285, L_286, L_287, L_288, L_289, L_290, L_291, L_292, L_293, L_294, L_295, L_296, L_297, L_298, L_299, L_300, L_301, L_302, L_303, L_304, L_305, L_306, L_307, L_308, L_309, L_310, L_311, L_312, L_313, L_314, L_315, L_316, L_317, L_318, L_319, L_320, L_321, L_322, L_323, L_324, L_325, L_326, L_327, L_328, L_329, L_330, L_331, L_332, L_333, L_334, L_335, L_336, L_337, L_338, L_339, L_340, L_341, L_342, L_343, L_344, L_345, L_346, L_347, L_348, L_349, L_350, L_351, L_352, L_353, L_354, L_355, L_356, L_357, L_358, L_359, L_360, L_361, L_362, L_363, L_364, L_365, L_366, L_367, L_368, L_369, L_370, L_371, L_372, L_373, L_374, L_375, L_376, L_377, L_378, L_379, L_380, L_381, L_382, L_383, L_384, L_385, L_386, L_387, L_388, L_389, L_390, L_391, L_392, L_393, L_394, L_395, L_396, L_397, L_398, L_399, L_400, L_401, L_402, L_403, L_404, L_405, L_406, L_407, L_408, L_409, L_410, L_411, L_412, L_413, L_414, L_415, L_416, L_417, L_418, L_419, L_420, L_421, L_422, L_423, L_424, L_425, L_426, L_427, L_428, L_429, L_430, L_431, L_432, L_433, L_434, L_435, L_436, L_437, L_438, L_439, L_440, L_441, L_442, L_443, L_444, L_445, L_446, L_447, L_448, L_449, L_450, L_451, L_452, L_453, L_454, L_455, L_456, L_457, L_458, L_459, L_460, L_461, L_462, L_463, L_464, L_465, L_466, L_467, L_468, L_469, L_470, L_471, L_472, L_473, L_474, L_475, L_476, L_477, L_478, L_479, L_480, L_481, L_482, L_483, L_484, L_485, L_486, L_487, L_488, L_489, L_490, L_491, L_492, L_493, L_494, L_495, L_496, L_497, L_498, L_499, L_500, L_501, L_502, L_503, L_504, L_505, L_506, L_507, L_508, L_509, L_510, L_511, L_512, L_513, L_514, L_515, L_516, L_517, L_518, L_519, L_520, L_521, L_522, L_523, L_524, L_525, L_526, L_527, L_528, L_529, L_530, L_531, L_532, L_533, L_534, L_535, L_536, L_537, L_538, L_539, L_540, L_541, L_542, L_543, L_544, L_545, L_546, L_547, L_548, L_549, L_550, L_551, L_552, L_553, L_554, L_555, L_556, L_557, L_558, L_559, L_560, L_561, L_562, L_563, L_564, L_565, L_566, L_567, L_568, L_569, L_570, L_571, L_572, L_573, L_574, L_575, L_576, L_577, L_578, L_579, L_580, L_581, L_582, L_583, L_584, L_585, L_586, L_587, L_588, L_589, L_590, L_591, L_592, L_593, L_594, L_595, L_596, L_597, L_598, L_599, L_600, L_601, L_602, L_603, L_604, L_605, L_606, L_607, L_608, L_609, L_610, L_611, L_612, L_613, L_614, L_615, L_616, L_617, L_618, L_619, L_620, L_621, L_622, L_623, L_624, L_625, L_626, L_627, L_628, L_629, L_630, L_631, L_632, L_633, L_634, L_635, L_636, L_637, L_638, L_639, L_640, L_641, L_642, L_643, L_644, L_645, L_646, L_647, L_648, L_649, L_650, L_651, L_652, L_653, L_654, L_655, L_656, L_657, L_658, L_659, L_660, L_661, L_662, L_663, L_664, L_665, L_666, L_667, L_668, L_669, L_670, L_671, L_672, L_673, L_674, L_675, L_676, L_677, L_678, L_679, L_680, L_681, L_682, L_683, L_684, L_685, L_686, L_687, L_688, L_689, L_690, L_691, L_692, L_693, L_694, L_695, L_696, L_697, L_698, L_699, L_700, L_701, L_702, L_703, L_704, L_705, L_706, L_707, L_708, L_709, L_710, L_711, L_712, L_713, L_714, L_715, L_716, L_717, L_718, L_719, L_720, L_721, L_722, L_723, L_724, L_725, L_726, L_727, L_728, L_729, L_730, L_731, L_732, L_733, L_734, L_735, L_736, L_737, L_738, L_739, L_740, L_741, L_742, L_743, L_744, L_745, L_746, L_747, L_748, L_749, L_750, L_751, L_752, L_753, L_754, L_755, L_756, L_757, L_758, L_759, L_760, L_761, L_762, L_763, L_764, L_765, L_766, L_767, L_768, L_769, L_770, L_771, L_772, L_773, L_774, L_775, L_776, L_777, L_778, L_779, L_780, L_781, L_782, L_783, L_784, L_785, L_786, L_787, L_788, L_789, L_790, L_791, L_792, L_793, L_794, L_795, L_796, L_797, L_798, L_799, L_800, L_801, L_802, L_803, L_804, L_805, L_806, L_807, L_808, L_809, L_810, L_811, L_812, L_813, L_814, L_815, L_816, L_817, L_818, L_819, L_820, L_821, L_822, L_823, L_824, L_825, L_826, L_827, L_828, L_829, L_830, L_831, L_832, L_833, L_834, L_835, L_836, L_837, L_838, L_839, L_840, L_841, L_842, L_843, L_844, L_845, L_846, L_847, L_848, L_849, L_850, L_851, L_852, L_853, L_854, L_855, L_856, L_857, L_858, L_859, L_860, L_861, L_862, L_863, L_864, L_865, L_866, L_867, L_868, L_869, L_870, L_871, L_872, L_873, L_874, L_875, L_876, L_877, L_878, L_879, L_880, L_881, L_882, L_883, L_884, L_885, L_886, L_887, L_888, L_889, L_890, L_891, L_892, L_893, L_894, L_895, L_896, L_897, L_898, L_899, L_900, L_901, L_902, L_903, L_904, L_905, L_906, L_907, L_908, L_909, L_910, L_911, L_912, L_913, L_914, L_915, L_916, L_917, L_918, L_919, L_920, L_921, L_922, L_923, L_924, L_925, L_926, L_927, L_928, L_929, L_930, L_931, L_932, L_933, L_934, L_935, L_936, L_937, L_938, L_939, L_940, L_941, L_942, L_943, L_944, L_945, L_946, L_947, L_948, L_949, L_950, L_951, L_952, L_953, L_954, L_955, L_956, L_957, L_958, L_959, L_960, L_961, L_962, L_963, L_964, L_965, L_966, L_967, L_968, L_969, L_970, L_971, L_972, L_973, L_974, L_975, L_976, L_977, L_978, L_979, L_980, L_981, L_982, L_983, L_984, L_985, L_986, L_987, L_988, L_989, L_990, L_991, L_992, L_993, L_994, L_995, L_996, L_997, L_998, L_999, L_1000, L_1001, L_1002, L_1003, L_1004, L_1005, L_1006, L_1007, L_1008, L_1009, L_1010, L_1011, L_1012, L_1013, L_1014, L_1015, L_1016, L_1017, L_1018, L_1019, L_1020, L_1021, L_1022, L_1023, L_1024, L_1025, L_1026, L_1027, L_1028, L_1029, L_1030, L_1031, L_1032, L_1033, L_1034, L_1035, L_1036, L_1037, L_1038, L_1039, L_1040, L_1041, L_1042, L_1043, L_1044, L_1045, L_1046, L_1047, L_1048, L_1049, L_1050, L_1051, L_1052, L_1053, L_1054, L_1055, L_1056, L_1057, L_1058, L_1059, L_1060, L_1061, L_1062, L_1063, L_1064, L_1065, L_1066, L_1067, L_1068, L_1069, L_1070, L_1071, L_1072, L_1073, L_1074, L_1075, L_1076, L_1077, L_1078, L_1079, L_1080, L_1081, L_1082, L_1083, L_1084, L_1085, L_1086, L_1087, L_1088, L_1089, L_1090, L_1091, L_1092, L_1093, L_1094, L_1095, L_1096, L_1097, L_1098, L_1099, L_1100, L_1101, L_1102, L_1103, L_1104, L_1105, L_1106, L_1107, L_1108, L_1109, L_1110, L_1111, L_1112, L_1113, L_1114, L_1115, L_1116, L_1117, L_1118, L_1119, L_1120, L_1121, L_1122, L_1123, L_1124, L_1125, L_1126, L_1127, L_1128, L_1129, L_1130, L_1131, L_1132, L_1133, L_1134, L_1135, L_1136, L_1137, L_1138, L_1139, L_1140, L_1141, L_1142, L_1143, L_1144, L_1145, L_1146, L_1147, L_1148, L_1149, L_1150, L_1151, L_1152, L_1153, L_1154, L_1155, L_1156, L_1157, L_1158, L_1159, L_1160, L_1161, L_1162, L_1163, L_1164, L_1165, L_1166, L_1167, L_1168, L_1169, L_1170, L_1171, L_1172, L_1173, L_1174, L_1175, L_1176, L_1177, L_1178, L_1179, L_1180, L_1181, L_1182, L_1183, L_1184, L_1185, L_1186, L_1187, L_1188, L_1189, L_1190, L_1191, L_1192, L_1193, L_1194, L_1195, L_1196, L_1197, L_1198, L_1199, L_1200, L_1201, L_1202, L_1203, L_1204, L_1205, L_1206, L_1207, L_1208, L_1209, L_1210, L_1211, L_1212, L_1213, L_1214, L_1215, L_1216, L_1217, L_1218, L_1219, L_1220, L_1221, L_1222, L_1223, L_1224, L_1225, L_1226, L_1227, L_1228, L_1229, L_1230, L_1231, L_1232, L_1233, L_1234, L_1235, L_1236, L_1237, L_1238, L_1239, L_1240, L_1241, L_1242, L_1243, L_1244, L_1245, L_1246, L_1247, L_1248, L_1249, L_1250, L_1251, L_1252, L_1253, L_1254, L_1255, L_1256, L_1257, L_1258, L_1259, L_1260, L_1261, L_1262, L_1263, L_1264, L_1265, L_1266, L_1267, L_1268, L_1269, L_1270, L_1271, L_1272, L_1273, L_1274, L_1275, L_1276, L_1277, L_1278, L_1279, L_1280, L_1281, L_1282, L_1283, L_1284, L_1285, L_1286, L_1287, L_1288, L_1289, L_1290, L_1291, L_1292, L_1293, L_1294, L_1295, L_1296, L_1297, L_1298, L_1299, L_1300, L_1301, L_1302, L_1303, L_1304, L_1305, L_1306, L_1307, L_1308, L_1309, L_1310, L_1311, L_1312, L_1313, L_1314, L_1315, L_1316, L_1317, L_1318, L_1319, L_1320, L_1321, L_1322, L_1323, L_1324, L_1325, L_1326, L_1327, L_1328, L_1329, L_1330, L_1331, L_1332, L_1333, L_1334, L_1335, L_1336, L_1337, L_1338, L_1339, L_1340, L_1341, L_1342, L_1343, L_1344, L_1345, L_1346, L_1347, L_1348, L_1349, L_1350, L_1351, L_1352, L_1353, L_1354, L_1355, L_1356, L_1357, L_1358, L_1359, L_1360, L_1361, L_1362, L_1363, L_1364, L_1365, L_1366, L_1367, L_1368, L_1369, L_1370, L_1371, L_1372, L_1373, L_1374, L_1375, L_1376, L_1377, L_1378, L_1379, L_1380, L_1381, L_1382, L_1383, L_1384, L_1385, L_1386, L_1387, L_1388, L_1389, L_1390, L_1391, L_1392, L_1393, L_1394, L_1395, L_1396, L_1397, L_1398, L_1399, L_1400, L_1401, L_1402, L_1403, L_1404, L_1405, L_1406, L_1407, L_1408, L_1409, L_1410, L_1411, L_1412, L_1413, L_1414, L_1415, L_1416, L_1417, L_1418, L_1419, L_1420, L_1421, L_1422, L_1423, L_1424, L_1425, L_1426, L_1427, L_1428, L_1429, L_1430, L_1431, L_1432, L_1433, L_1434, L_1435, L_1436, L_1437, L_1438, L_1439, L_1440;
wire [quan_width - 1:0] C2V_1_5, C2V_1_89, C2V_1_109, C2V_1_170, C2V_1_232, C2V_1_275, C2V_1_375, C2V_1_429, C2V_1_526, C2V_1_762, C2V_1_810, C2V_1_858, C2V_1_899, C2V_1_940, C2V_1_974, C2V_1_1013, C2V_1_1087, C2V_1_1146, C2V_1_1153, C2V_2_14, C2V_2_63, C2V_2_119, C2V_2_167, C2V_2_196, C2V_2_265, C2V_2_316, C2V_2_423, C2V_2_512, C2V_2_672, C2V_2_685, C2V_2_853, C2V_2_895, C2V_2_958, C2V_2_989, C2V_2_1021, C2V_2_1088, C2V_2_1119, C2V_2_1153, C2V_2_1154, C2V_3_9, C2V_3_84, C2V_3_101, C2V_3_183, C2V_3_201, C2V_3_268, C2V_3_365, C2V_3_420, C2V_3_531, C2V_3_588, C2V_3_664, C2V_3_768, C2V_3_899, C2V_3_943, C2V_3_968, C2V_3_1028, C2V_3_1058, C2V_3_1151, C2V_3_1154, C2V_3_1155, C2V_4_28, C2V_4_87, C2V_4_126, C2V_4_182, C2V_4_199, C2V_4_253, C2V_4_477, C2V_4_517, C2V_4_553, C2V_4_615, C2V_4_640, C2V_4_686, C2V_4_903, C2V_4_927, C2V_4_963, C2V_4_1041, C2V_4_1068, C2V_4_1132, C2V_4_1155, C2V_4_1156, C2V_5_47, C2V_5_57, C2V_5_140, C2V_5_163, C2V_5_227, C2V_5_245, C2V_5_294, C2V_5_361, C2V_5_440, C2V_5_674, C2V_5_738, C2V_5_792, C2V_5_870, C2V_5_918, C2V_5_961, C2V_5_1013, C2V_5_1062, C2V_5_1110, C2V_5_1156, C2V_5_1157, C2V_6_30, C2V_6_54, C2V_6_142, C2V_6_162, C2V_6_196, C2V_6_275, C2V_6_328, C2V_6_480, C2V_6_529, C2V_6_610, C2V_6_814, C2V_6_842, C2V_6_875, C2V_6_937, C2V_6_972, C2V_6_1039, C2V_6_1103, C2V_6_1105, C2V_6_1157, C2V_6_1158, C2V_7_6, C2V_7_90, C2V_7_110, C2V_7_171, C2V_7_233, C2V_7_276, C2V_7_376, C2V_7_430, C2V_7_527, C2V_7_763, C2V_7_811, C2V_7_859, C2V_7_900, C2V_7_941, C2V_7_975, C2V_7_1014, C2V_7_1088, C2V_7_1147, C2V_7_1158, C2V_7_1159, C2V_8_15, C2V_8_64, C2V_8_120, C2V_8_168, C2V_8_197, C2V_8_266, C2V_8_317, C2V_8_424, C2V_8_513, C2V_8_625, C2V_8_686, C2V_8_854, C2V_8_896, C2V_8_959, C2V_8_990, C2V_8_1022, C2V_8_1089, C2V_8_1120, C2V_8_1159, C2V_8_1160, C2V_9_10, C2V_9_85, C2V_9_102, C2V_9_184, C2V_9_202, C2V_9_269, C2V_9_366, C2V_9_421, C2V_9_532, C2V_9_589, C2V_9_665, C2V_9_721, C2V_9_900, C2V_9_944, C2V_9_969, C2V_9_1029, C2V_9_1059, C2V_9_1152, C2V_9_1160, C2V_9_1161, C2V_10_29, C2V_10_88, C2V_10_127, C2V_10_183, C2V_10_200, C2V_10_254, C2V_10_478, C2V_10_518, C2V_10_554, C2V_10_616, C2V_10_641, C2V_10_687, C2V_10_904, C2V_10_928, C2V_10_964, C2V_10_1042, C2V_10_1069, C2V_10_1133, C2V_10_1161, C2V_10_1162, C2V_11_48, C2V_11_58, C2V_11_141, C2V_11_164, C2V_11_228, C2V_11_246, C2V_11_295, C2V_11_362, C2V_11_441, C2V_11_675, C2V_11_739, C2V_11_793, C2V_11_871, C2V_11_919, C2V_11_962, C2V_11_1014, C2V_11_1063, C2V_11_1111, C2V_11_1162, C2V_11_1163, C2V_12_31, C2V_12_55, C2V_12_143, C2V_12_163, C2V_12_197, C2V_12_276, C2V_12_329, C2V_12_433, C2V_12_530, C2V_12_611, C2V_12_815, C2V_12_843, C2V_12_876, C2V_12_938, C2V_12_973, C2V_12_1040, C2V_12_1104, C2V_12_1106, C2V_12_1163, C2V_12_1164, C2V_13_7, C2V_13_91, C2V_13_111, C2V_13_172, C2V_13_234, C2V_13_277, C2V_13_377, C2V_13_431, C2V_13_528, C2V_13_764, C2V_13_812, C2V_13_860, C2V_13_901, C2V_13_942, C2V_13_976, C2V_13_1015, C2V_13_1089, C2V_13_1148, C2V_13_1164, C2V_13_1165, C2V_14_16, C2V_14_65, C2V_14_121, C2V_14_169, C2V_14_198, C2V_14_267, C2V_14_318, C2V_14_425, C2V_14_514, C2V_14_626, C2V_14_687, C2V_14_855, C2V_14_897, C2V_14_960, C2V_14_991, C2V_14_1023, C2V_14_1090, C2V_14_1121, C2V_14_1165, C2V_14_1166, C2V_15_11, C2V_15_86, C2V_15_103, C2V_15_185, C2V_15_203, C2V_15_270, C2V_15_367, C2V_15_422, C2V_15_533, C2V_15_590, C2V_15_666, C2V_15_722, C2V_15_901, C2V_15_945, C2V_15_970, C2V_15_1030, C2V_15_1060, C2V_15_1105, C2V_15_1166, C2V_15_1167, C2V_16_30, C2V_16_89, C2V_16_128, C2V_16_184, C2V_16_201, C2V_16_255, C2V_16_479, C2V_16_519, C2V_16_555, C2V_16_617, C2V_16_642, C2V_16_688, C2V_16_905, C2V_16_929, C2V_16_965, C2V_16_1043, C2V_16_1070, C2V_16_1134, C2V_16_1167, C2V_16_1168, C2V_17_1, C2V_17_59, C2V_17_142, C2V_17_165, C2V_17_229, C2V_17_247, C2V_17_296, C2V_17_363, C2V_17_442, C2V_17_676, C2V_17_740, C2V_17_794, C2V_17_872, C2V_17_920, C2V_17_963, C2V_17_1015, C2V_17_1064, C2V_17_1112, C2V_17_1168, C2V_17_1169, C2V_18_32, C2V_18_56, C2V_18_144, C2V_18_164, C2V_18_198, C2V_18_277, C2V_18_330, C2V_18_434, C2V_18_531, C2V_18_612, C2V_18_816, C2V_18_844, C2V_18_877, C2V_18_939, C2V_18_974, C2V_18_1041, C2V_18_1057, C2V_18_1107, C2V_18_1169, C2V_18_1170, C2V_19_8, C2V_19_92, C2V_19_112, C2V_19_173, C2V_19_235, C2V_19_278, C2V_19_378, C2V_19_432, C2V_19_481, C2V_19_765, C2V_19_813, C2V_19_861, C2V_19_902, C2V_19_943, C2V_19_977, C2V_19_1016, C2V_19_1090, C2V_19_1149, C2V_19_1170, C2V_19_1171, C2V_20_17, C2V_20_66, C2V_20_122, C2V_20_170, C2V_20_199, C2V_20_268, C2V_20_319, C2V_20_426, C2V_20_515, C2V_20_627, C2V_20_688, C2V_20_856, C2V_20_898, C2V_20_913, C2V_20_992, C2V_20_1024, C2V_20_1091, C2V_20_1122, C2V_20_1171, C2V_20_1172, C2V_21_12, C2V_21_87, C2V_21_104, C2V_21_186, C2V_21_204, C2V_21_271, C2V_21_368, C2V_21_423, C2V_21_534, C2V_21_591, C2V_21_667, C2V_21_723, C2V_21_902, C2V_21_946, C2V_21_971, C2V_21_1031, C2V_21_1061, C2V_21_1106, C2V_21_1172, C2V_21_1173, C2V_22_31, C2V_22_90, C2V_22_129, C2V_22_185, C2V_22_202, C2V_22_256, C2V_22_480, C2V_22_520, C2V_22_556, C2V_22_618, C2V_22_643, C2V_22_689, C2V_22_906, C2V_22_930, C2V_22_966, C2V_22_1044, C2V_22_1071, C2V_22_1135, C2V_22_1173, C2V_22_1174, C2V_23_2, C2V_23_60, C2V_23_143, C2V_23_166, C2V_23_230, C2V_23_248, C2V_23_297, C2V_23_364, C2V_23_443, C2V_23_677, C2V_23_741, C2V_23_795, C2V_23_873, C2V_23_921, C2V_23_964, C2V_23_1016, C2V_23_1065, C2V_23_1113, C2V_23_1174, C2V_23_1175, C2V_24_33, C2V_24_57, C2V_24_97, C2V_24_165, C2V_24_199, C2V_24_278, C2V_24_331, C2V_24_435, C2V_24_532, C2V_24_613, C2V_24_769, C2V_24_845, C2V_24_878, C2V_24_940, C2V_24_975, C2V_24_1042, C2V_24_1058, C2V_24_1108, C2V_24_1175, C2V_24_1176, C2V_25_9, C2V_25_93, C2V_25_113, C2V_25_174, C2V_25_236, C2V_25_279, C2V_25_379, C2V_25_385, C2V_25_482, C2V_25_766, C2V_25_814, C2V_25_862, C2V_25_903, C2V_25_944, C2V_25_978, C2V_25_1017, C2V_25_1091, C2V_25_1150, C2V_25_1176, C2V_25_1177, C2V_26_18, C2V_26_67, C2V_26_123, C2V_26_171, C2V_26_200, C2V_26_269, C2V_26_320, C2V_26_427, C2V_26_516, C2V_26_628, C2V_26_689, C2V_26_857, C2V_26_899, C2V_26_914, C2V_26_993, C2V_26_1025, C2V_26_1092, C2V_26_1123, C2V_26_1177, C2V_26_1178, C2V_27_13, C2V_27_88, C2V_27_105, C2V_27_187, C2V_27_205, C2V_27_272, C2V_27_369, C2V_27_424, C2V_27_535, C2V_27_592, C2V_27_668, C2V_27_724, C2V_27_903, C2V_27_947, C2V_27_972, C2V_27_1032, C2V_27_1062, C2V_27_1107, C2V_27_1178, C2V_27_1179, C2V_28_32, C2V_28_91, C2V_28_130, C2V_28_186, C2V_28_203, C2V_28_257, C2V_28_433, C2V_28_521, C2V_28_557, C2V_28_619, C2V_28_644, C2V_28_690, C2V_28_907, C2V_28_931, C2V_28_967, C2V_28_1045, C2V_28_1072, C2V_28_1136, C2V_28_1179, C2V_28_1180, C2V_29_3, C2V_29_61, C2V_29_144, C2V_29_167, C2V_29_231, C2V_29_249, C2V_29_298, C2V_29_365, C2V_29_444, C2V_29_678, C2V_29_742, C2V_29_796, C2V_29_874, C2V_29_922, C2V_29_965, C2V_29_1017, C2V_29_1066, C2V_29_1114, C2V_29_1180, C2V_29_1181, C2V_30_34, C2V_30_58, C2V_30_98, C2V_30_166, C2V_30_200, C2V_30_279, C2V_30_332, C2V_30_436, C2V_30_533, C2V_30_614, C2V_30_770, C2V_30_846, C2V_30_879, C2V_30_941, C2V_30_976, C2V_30_1043, C2V_30_1059, C2V_30_1109, C2V_30_1181, C2V_30_1182, C2V_31_10, C2V_31_94, C2V_31_114, C2V_31_175, C2V_31_237, C2V_31_280, C2V_31_380, C2V_31_386, C2V_31_483, C2V_31_767, C2V_31_815, C2V_31_863, C2V_31_904, C2V_31_945, C2V_31_979, C2V_31_1018, C2V_31_1092, C2V_31_1151, C2V_31_1182, C2V_31_1183, C2V_32_19, C2V_32_68, C2V_32_124, C2V_32_172, C2V_32_201, C2V_32_270, C2V_32_321, C2V_32_428, C2V_32_517, C2V_32_629, C2V_32_690, C2V_32_858, C2V_32_900, C2V_32_915, C2V_32_994, C2V_32_1026, C2V_32_1093, C2V_32_1124, C2V_32_1183, C2V_32_1184, C2V_33_14, C2V_33_89, C2V_33_106, C2V_33_188, C2V_33_206, C2V_33_273, C2V_33_370, C2V_33_425, C2V_33_536, C2V_33_593, C2V_33_669, C2V_33_725, C2V_33_904, C2V_33_948, C2V_33_973, C2V_33_1033, C2V_33_1063, C2V_33_1108, C2V_33_1184, C2V_33_1185, C2V_34_33, C2V_34_92, C2V_34_131, C2V_34_187, C2V_34_204, C2V_34_258, C2V_34_434, C2V_34_522, C2V_34_558, C2V_34_620, C2V_34_645, C2V_34_691, C2V_34_908, C2V_34_932, C2V_34_968, C2V_34_1046, C2V_34_1073, C2V_34_1137, C2V_34_1185, C2V_34_1186, C2V_35_4, C2V_35_62, C2V_35_97, C2V_35_168, C2V_35_232, C2V_35_250, C2V_35_299, C2V_35_366, C2V_35_445, C2V_35_679, C2V_35_743, C2V_35_797, C2V_35_875, C2V_35_923, C2V_35_966, C2V_35_1018, C2V_35_1067, C2V_35_1115, C2V_35_1186, C2V_35_1187, C2V_36_35, C2V_36_59, C2V_36_99, C2V_36_167, C2V_36_201, C2V_36_280, C2V_36_333, C2V_36_437, C2V_36_534, C2V_36_615, C2V_36_771, C2V_36_847, C2V_36_880, C2V_36_942, C2V_36_977, C2V_36_1044, C2V_36_1060, C2V_36_1110, C2V_36_1187, C2V_36_1188, C2V_37_11, C2V_37_95, C2V_37_115, C2V_37_176, C2V_37_238, C2V_37_281, C2V_37_381, C2V_37_387, C2V_37_484, C2V_37_768, C2V_37_816, C2V_37_864, C2V_37_905, C2V_37_946, C2V_37_980, C2V_37_1019, C2V_37_1093, C2V_37_1152, C2V_37_1188, C2V_37_1189, C2V_38_20, C2V_38_69, C2V_38_125, C2V_38_173, C2V_38_202, C2V_38_271, C2V_38_322, C2V_38_429, C2V_38_518, C2V_38_630, C2V_38_691, C2V_38_859, C2V_38_901, C2V_38_916, C2V_38_995, C2V_38_1027, C2V_38_1094, C2V_38_1125, C2V_38_1189, C2V_38_1190, C2V_39_15, C2V_39_90, C2V_39_107, C2V_39_189, C2V_39_207, C2V_39_274, C2V_39_371, C2V_39_426, C2V_39_537, C2V_39_594, C2V_39_670, C2V_39_726, C2V_39_905, C2V_39_949, C2V_39_974, C2V_39_1034, C2V_39_1064, C2V_39_1109, C2V_39_1190, C2V_39_1191, C2V_40_34, C2V_40_93, C2V_40_132, C2V_40_188, C2V_40_205, C2V_40_259, C2V_40_435, C2V_40_523, C2V_40_559, C2V_40_621, C2V_40_646, C2V_40_692, C2V_40_909, C2V_40_933, C2V_40_969, C2V_40_1047, C2V_40_1074, C2V_40_1138, C2V_40_1191, C2V_40_1192, C2V_41_5, C2V_41_63, C2V_41_98, C2V_41_169, C2V_41_233, C2V_41_251, C2V_41_300, C2V_41_367, C2V_41_446, C2V_41_680, C2V_41_744, C2V_41_798, C2V_41_876, C2V_41_924, C2V_41_967, C2V_41_1019, C2V_41_1068, C2V_41_1116, C2V_41_1192, C2V_41_1193, C2V_42_36, C2V_42_60, C2V_42_100, C2V_42_168, C2V_42_202, C2V_42_281, C2V_42_334, C2V_42_438, C2V_42_535, C2V_42_616, C2V_42_772, C2V_42_848, C2V_42_881, C2V_42_943, C2V_42_978, C2V_42_1045, C2V_42_1061, C2V_42_1111, C2V_42_1193, C2V_42_1194, C2V_43_12, C2V_43_96, C2V_43_116, C2V_43_177, C2V_43_239, C2V_43_282, C2V_43_382, C2V_43_388, C2V_43_485, C2V_43_721, C2V_43_769, C2V_43_817, C2V_43_906, C2V_43_947, C2V_43_981, C2V_43_1020, C2V_43_1094, C2V_43_1105, C2V_43_1194, C2V_43_1195, C2V_44_21, C2V_44_70, C2V_44_126, C2V_44_174, C2V_44_203, C2V_44_272, C2V_44_323, C2V_44_430, C2V_44_519, C2V_44_631, C2V_44_692, C2V_44_860, C2V_44_902, C2V_44_917, C2V_44_996, C2V_44_1028, C2V_44_1095, C2V_44_1126, C2V_44_1195, C2V_44_1196, C2V_45_16, C2V_45_91, C2V_45_108, C2V_45_190, C2V_45_208, C2V_45_275, C2V_45_372, C2V_45_427, C2V_45_538, C2V_45_595, C2V_45_671, C2V_45_727, C2V_45_906, C2V_45_950, C2V_45_975, C2V_45_1035, C2V_45_1065, C2V_45_1110, C2V_45_1196, C2V_45_1197, C2V_46_35, C2V_46_94, C2V_46_133, C2V_46_189, C2V_46_206, C2V_46_260, C2V_46_436, C2V_46_524, C2V_46_560, C2V_46_622, C2V_46_647, C2V_46_693, C2V_46_910, C2V_46_934, C2V_46_970, C2V_46_1048, C2V_46_1075, C2V_46_1139, C2V_46_1197, C2V_46_1198, C2V_47_6, C2V_47_64, C2V_47_99, C2V_47_170, C2V_47_234, C2V_47_252, C2V_47_301, C2V_47_368, C2V_47_447, C2V_47_681, C2V_47_745, C2V_47_799, C2V_47_877, C2V_47_925, C2V_47_968, C2V_47_1020, C2V_47_1069, C2V_47_1117, C2V_47_1198, C2V_47_1199, C2V_48_37, C2V_48_61, C2V_48_101, C2V_48_169, C2V_48_203, C2V_48_282, C2V_48_335, C2V_48_439, C2V_48_536, C2V_48_617, C2V_48_773, C2V_48_849, C2V_48_882, C2V_48_944, C2V_48_979, C2V_48_1046, C2V_48_1062, C2V_48_1112, C2V_48_1199, C2V_48_1200, C2V_49_13, C2V_49_49, C2V_49_117, C2V_49_178, C2V_49_240, C2V_49_283, C2V_49_383, C2V_49_389, C2V_49_486, C2V_49_722, C2V_49_770, C2V_49_818, C2V_49_907, C2V_49_948, C2V_49_982, C2V_49_1021, C2V_49_1095, C2V_49_1106, C2V_49_1200, C2V_49_1201, C2V_50_22, C2V_50_71, C2V_50_127, C2V_50_175, C2V_50_204, C2V_50_273, C2V_50_324, C2V_50_431, C2V_50_520, C2V_50_632, C2V_50_693, C2V_50_861, C2V_50_903, C2V_50_918, C2V_50_997, C2V_50_1029, C2V_50_1096, C2V_50_1127, C2V_50_1201, C2V_50_1202, C2V_51_17, C2V_51_92, C2V_51_109, C2V_51_191, C2V_51_209, C2V_51_276, C2V_51_373, C2V_51_428, C2V_51_539, C2V_51_596, C2V_51_672, C2V_51_728, C2V_51_907, C2V_51_951, C2V_51_976, C2V_51_1036, C2V_51_1066, C2V_51_1111, C2V_51_1202, C2V_51_1203, C2V_52_36, C2V_52_95, C2V_52_134, C2V_52_190, C2V_52_207, C2V_52_261, C2V_52_437, C2V_52_525, C2V_52_561, C2V_52_623, C2V_52_648, C2V_52_694, C2V_52_911, C2V_52_935, C2V_52_971, C2V_52_1049, C2V_52_1076, C2V_52_1140, C2V_52_1203, C2V_52_1204, C2V_53_7, C2V_53_65, C2V_53_100, C2V_53_171, C2V_53_235, C2V_53_253, C2V_53_302, C2V_53_369, C2V_53_448, C2V_53_682, C2V_53_746, C2V_53_800, C2V_53_878, C2V_53_926, C2V_53_969, C2V_53_1021, C2V_53_1070, C2V_53_1118, C2V_53_1204, C2V_53_1205, C2V_54_38, C2V_54_62, C2V_54_102, C2V_54_170, C2V_54_204, C2V_54_283, C2V_54_336, C2V_54_440, C2V_54_537, C2V_54_618, C2V_54_774, C2V_54_850, C2V_54_883, C2V_54_945, C2V_54_980, C2V_54_1047, C2V_54_1063, C2V_54_1113, C2V_54_1205, C2V_54_1206, C2V_55_14, C2V_55_50, C2V_55_118, C2V_55_179, C2V_55_193, C2V_55_284, C2V_55_384, C2V_55_390, C2V_55_487, C2V_55_723, C2V_55_771, C2V_55_819, C2V_55_908, C2V_55_949, C2V_55_983, C2V_55_1022, C2V_55_1096, C2V_55_1107, C2V_55_1206, C2V_55_1207, C2V_56_23, C2V_56_72, C2V_56_128, C2V_56_176, C2V_56_205, C2V_56_274, C2V_56_325, C2V_56_432, C2V_56_521, C2V_56_633, C2V_56_694, C2V_56_862, C2V_56_904, C2V_56_919, C2V_56_998, C2V_56_1030, C2V_56_1097, C2V_56_1128, C2V_56_1207, C2V_56_1208, C2V_57_18, C2V_57_93, C2V_57_110, C2V_57_192, C2V_57_210, C2V_57_277, C2V_57_374, C2V_57_429, C2V_57_540, C2V_57_597, C2V_57_625, C2V_57_729, C2V_57_908, C2V_57_952, C2V_57_977, C2V_57_1037, C2V_57_1067, C2V_57_1112, C2V_57_1208, C2V_57_1209, C2V_58_37, C2V_58_96, C2V_58_135, C2V_58_191, C2V_58_208, C2V_58_262, C2V_58_438, C2V_58_526, C2V_58_562, C2V_58_624, C2V_58_649, C2V_58_695, C2V_58_912, C2V_58_936, C2V_58_972, C2V_58_1050, C2V_58_1077, C2V_58_1141, C2V_58_1209, C2V_58_1210, C2V_59_8, C2V_59_66, C2V_59_101, C2V_59_172, C2V_59_236, C2V_59_254, C2V_59_303, C2V_59_370, C2V_59_449, C2V_59_683, C2V_59_747, C2V_59_801, C2V_59_879, C2V_59_927, C2V_59_970, C2V_59_1022, C2V_59_1071, C2V_59_1119, C2V_59_1210, C2V_59_1211, C2V_60_39, C2V_60_63, C2V_60_103, C2V_60_171, C2V_60_205, C2V_60_284, C2V_60_289, C2V_60_441, C2V_60_538, C2V_60_619, C2V_60_775, C2V_60_851, C2V_60_884, C2V_60_946, C2V_60_981, C2V_60_1048, C2V_60_1064, C2V_60_1114, C2V_60_1211, C2V_60_1212, C2V_61_15, C2V_61_51, C2V_61_119, C2V_61_180, C2V_61_194, C2V_61_285, C2V_61_337, C2V_61_391, C2V_61_488, C2V_61_724, C2V_61_772, C2V_61_820, C2V_61_909, C2V_61_950, C2V_61_984, C2V_61_1023, C2V_61_1097, C2V_61_1108, C2V_61_1212, C2V_61_1213, C2V_62_24, C2V_62_73, C2V_62_129, C2V_62_177, C2V_62_206, C2V_62_275, C2V_62_326, C2V_62_385, C2V_62_522, C2V_62_634, C2V_62_695, C2V_62_863, C2V_62_905, C2V_62_920, C2V_62_999, C2V_62_1031, C2V_62_1098, C2V_62_1129, C2V_62_1213, C2V_62_1214, C2V_63_19, C2V_63_94, C2V_63_111, C2V_63_145, C2V_63_211, C2V_63_278, C2V_63_375, C2V_63_430, C2V_63_541, C2V_63_598, C2V_63_626, C2V_63_730, C2V_63_909, C2V_63_953, C2V_63_978, C2V_63_1038, C2V_63_1068, C2V_63_1113, C2V_63_1214, C2V_63_1215, C2V_64_38, C2V_64_49, C2V_64_136, C2V_64_192, C2V_64_209, C2V_64_263, C2V_64_439, C2V_64_527, C2V_64_563, C2V_64_577, C2V_64_650, C2V_64_696, C2V_64_865, C2V_64_937, C2V_64_973, C2V_64_1051, C2V_64_1078, C2V_64_1142, C2V_64_1215, C2V_64_1216, C2V_65_9, C2V_65_67, C2V_65_102, C2V_65_173, C2V_65_237, C2V_65_255, C2V_65_304, C2V_65_371, C2V_65_450, C2V_65_684, C2V_65_748, C2V_65_802, C2V_65_880, C2V_65_928, C2V_65_971, C2V_65_1023, C2V_65_1072, C2V_65_1120, C2V_65_1216, C2V_65_1217, C2V_66_40, C2V_66_64, C2V_66_104, C2V_66_172, C2V_66_206, C2V_66_285, C2V_66_290, C2V_66_442, C2V_66_539, C2V_66_620, C2V_66_776, C2V_66_852, C2V_66_885, C2V_66_947, C2V_66_982, C2V_66_1049, C2V_66_1065, C2V_66_1115, C2V_66_1217, C2V_66_1218, C2V_67_16, C2V_67_52, C2V_67_120, C2V_67_181, C2V_67_195, C2V_67_286, C2V_67_338, C2V_67_392, C2V_67_489, C2V_67_725, C2V_67_773, C2V_67_821, C2V_67_910, C2V_67_951, C2V_67_985, C2V_67_1024, C2V_67_1098, C2V_67_1109, C2V_67_1218, C2V_67_1219, C2V_68_25, C2V_68_74, C2V_68_130, C2V_68_178, C2V_68_207, C2V_68_276, C2V_68_327, C2V_68_386, C2V_68_523, C2V_68_635, C2V_68_696, C2V_68_864, C2V_68_906, C2V_68_921, C2V_68_1000, C2V_68_1032, C2V_68_1099, C2V_68_1130, C2V_68_1219, C2V_68_1220, C2V_69_20, C2V_69_95, C2V_69_112, C2V_69_146, C2V_69_212, C2V_69_279, C2V_69_376, C2V_69_431, C2V_69_542, C2V_69_599, C2V_69_627, C2V_69_731, C2V_69_910, C2V_69_954, C2V_69_979, C2V_69_1039, C2V_69_1069, C2V_69_1114, C2V_69_1220, C2V_69_1221, C2V_70_39, C2V_70_50, C2V_70_137, C2V_70_145, C2V_70_210, C2V_70_264, C2V_70_440, C2V_70_528, C2V_70_564, C2V_70_578, C2V_70_651, C2V_70_697, C2V_70_866, C2V_70_938, C2V_70_974, C2V_70_1052, C2V_70_1079, C2V_70_1143, C2V_70_1221, C2V_70_1222, C2V_71_10, C2V_71_68, C2V_71_103, C2V_71_174, C2V_71_238, C2V_71_256, C2V_71_305, C2V_71_372, C2V_71_451, C2V_71_685, C2V_71_749, C2V_71_803, C2V_71_881, C2V_71_929, C2V_71_972, C2V_71_1024, C2V_71_1073, C2V_71_1121, C2V_71_1222, C2V_71_1223, C2V_72_41, C2V_72_65, C2V_72_105, C2V_72_173, C2V_72_207, C2V_72_286, C2V_72_291, C2V_72_443, C2V_72_540, C2V_72_621, C2V_72_777, C2V_72_853, C2V_72_886, C2V_72_948, C2V_72_983, C2V_72_1050, C2V_72_1066, C2V_72_1116, C2V_72_1223, C2V_72_1224, C2V_73_17, C2V_73_53, C2V_73_121, C2V_73_182, C2V_73_196, C2V_73_287, C2V_73_339, C2V_73_393, C2V_73_490, C2V_73_726, C2V_73_774, C2V_73_822, C2V_73_911, C2V_73_952, C2V_73_986, C2V_73_1025, C2V_73_1099, C2V_73_1110, C2V_73_1224, C2V_73_1225, C2V_74_26, C2V_74_75, C2V_74_131, C2V_74_179, C2V_74_208, C2V_74_277, C2V_74_328, C2V_74_387, C2V_74_524, C2V_74_636, C2V_74_697, C2V_74_817, C2V_74_907, C2V_74_922, C2V_74_1001, C2V_74_1033, C2V_74_1100, C2V_74_1131, C2V_74_1225, C2V_74_1226, C2V_75_21, C2V_75_96, C2V_75_113, C2V_75_147, C2V_75_213, C2V_75_280, C2V_75_377, C2V_75_432, C2V_75_543, C2V_75_600, C2V_75_628, C2V_75_732, C2V_75_911, C2V_75_955, C2V_75_980, C2V_75_1040, C2V_75_1070, C2V_75_1115, C2V_75_1226, C2V_75_1227, C2V_76_40, C2V_76_51, C2V_76_138, C2V_76_146, C2V_76_211, C2V_76_265, C2V_76_441, C2V_76_481, C2V_76_565, C2V_76_579, C2V_76_652, C2V_76_698, C2V_76_867, C2V_76_939, C2V_76_975, C2V_76_1053, C2V_76_1080, C2V_76_1144, C2V_76_1227, C2V_76_1228, C2V_77_11, C2V_77_69, C2V_77_104, C2V_77_175, C2V_77_239, C2V_77_257, C2V_77_306, C2V_77_373, C2V_77_452, C2V_77_686, C2V_77_750, C2V_77_804, C2V_77_882, C2V_77_930, C2V_77_973, C2V_77_1025, C2V_77_1074, C2V_77_1122, C2V_77_1228, C2V_77_1229, C2V_78_42, C2V_78_66, C2V_78_106, C2V_78_174, C2V_78_208, C2V_78_287, C2V_78_292, C2V_78_444, C2V_78_541, C2V_78_622, C2V_78_778, C2V_78_854, C2V_78_887, C2V_78_949, C2V_78_984, C2V_78_1051, C2V_78_1067, C2V_78_1117, C2V_78_1229, C2V_78_1230, C2V_79_18, C2V_79_54, C2V_79_122, C2V_79_183, C2V_79_197, C2V_79_288, C2V_79_340, C2V_79_394, C2V_79_491, C2V_79_727, C2V_79_775, C2V_79_823, C2V_79_912, C2V_79_953, C2V_79_987, C2V_79_1026, C2V_79_1100, C2V_79_1111, C2V_79_1230, C2V_79_1231, C2V_80_27, C2V_80_76, C2V_80_132, C2V_80_180, C2V_80_209, C2V_80_278, C2V_80_329, C2V_80_388, C2V_80_525, C2V_80_637, C2V_80_698, C2V_80_818, C2V_80_908, C2V_80_923, C2V_80_1002, C2V_80_1034, C2V_80_1101, C2V_80_1132, C2V_80_1231, C2V_80_1232, C2V_81_22, C2V_81_49, C2V_81_114, C2V_81_148, C2V_81_214, C2V_81_281, C2V_81_378, C2V_81_385, C2V_81_544, C2V_81_601, C2V_81_629, C2V_81_733, C2V_81_912, C2V_81_956, C2V_81_981, C2V_81_1041, C2V_81_1071, C2V_81_1116, C2V_81_1232, C2V_81_1233, C2V_82_41, C2V_82_52, C2V_82_139, C2V_82_147, C2V_82_212, C2V_82_266, C2V_82_442, C2V_82_482, C2V_82_566, C2V_82_580, C2V_82_653, C2V_82_699, C2V_82_868, C2V_82_940, C2V_82_976, C2V_82_1054, C2V_82_1081, C2V_82_1145, C2V_82_1233, C2V_82_1234, C2V_83_12, C2V_83_70, C2V_83_105, C2V_83_176, C2V_83_240, C2V_83_258, C2V_83_307, C2V_83_374, C2V_83_453, C2V_83_687, C2V_83_751, C2V_83_805, C2V_83_883, C2V_83_931, C2V_83_974, C2V_83_1026, C2V_83_1075, C2V_83_1123, C2V_83_1234, C2V_83_1235, C2V_84_43, C2V_84_67, C2V_84_107, C2V_84_175, C2V_84_209, C2V_84_288, C2V_84_293, C2V_84_445, C2V_84_542, C2V_84_623, C2V_84_779, C2V_84_855, C2V_84_888, C2V_84_950, C2V_84_985, C2V_84_1052, C2V_84_1068, C2V_84_1118, C2V_84_1235, C2V_84_1236, C2V_85_19, C2V_85_55, C2V_85_123, C2V_85_184, C2V_85_198, C2V_85_241, C2V_85_341, C2V_85_395, C2V_85_492, C2V_85_728, C2V_85_776, C2V_85_824, C2V_85_865, C2V_85_954, C2V_85_988, C2V_85_1027, C2V_85_1101, C2V_85_1112, C2V_85_1236, C2V_85_1237, C2V_86_28, C2V_86_77, C2V_86_133, C2V_86_181, C2V_86_210, C2V_86_279, C2V_86_330, C2V_86_389, C2V_86_526, C2V_86_638, C2V_86_699, C2V_86_819, C2V_86_909, C2V_86_924, C2V_86_1003, C2V_86_1035, C2V_86_1102, C2V_86_1133, C2V_86_1237, C2V_86_1238, C2V_87_23, C2V_87_50, C2V_87_115, C2V_87_149, C2V_87_215, C2V_87_282, C2V_87_379, C2V_87_386, C2V_87_545, C2V_87_602, C2V_87_630, C2V_87_734, C2V_87_865, C2V_87_957, C2V_87_982, C2V_87_1042, C2V_87_1072, C2V_87_1117, C2V_87_1238, C2V_87_1239, C2V_88_42, C2V_88_53, C2V_88_140, C2V_88_148, C2V_88_213, C2V_88_267, C2V_88_443, C2V_88_483, C2V_88_567, C2V_88_581, C2V_88_654, C2V_88_700, C2V_88_869, C2V_88_941, C2V_88_977, C2V_88_1055, C2V_88_1082, C2V_88_1146, C2V_88_1239, C2V_88_1240, C2V_89_13, C2V_89_71, C2V_89_106, C2V_89_177, C2V_89_193, C2V_89_259, C2V_89_308, C2V_89_375, C2V_89_454, C2V_89_688, C2V_89_752, C2V_89_806, C2V_89_884, C2V_89_932, C2V_89_975, C2V_89_1027, C2V_89_1076, C2V_89_1124, C2V_89_1240, C2V_89_1241, C2V_90_44, C2V_90_68, C2V_90_108, C2V_90_176, C2V_90_210, C2V_90_241, C2V_90_294, C2V_90_446, C2V_90_543, C2V_90_624, C2V_90_780, C2V_90_856, C2V_90_889, C2V_90_951, C2V_90_986, C2V_90_1053, C2V_90_1069, C2V_90_1119, C2V_90_1241, C2V_90_1242, C2V_91_20, C2V_91_56, C2V_91_124, C2V_91_185, C2V_91_199, C2V_91_242, C2V_91_342, C2V_91_396, C2V_91_493, C2V_91_729, C2V_91_777, C2V_91_825, C2V_91_866, C2V_91_955, C2V_91_989, C2V_91_1028, C2V_91_1102, C2V_91_1113, C2V_91_1242, C2V_91_1243, C2V_92_29, C2V_92_78, C2V_92_134, C2V_92_182, C2V_92_211, C2V_92_280, C2V_92_331, C2V_92_390, C2V_92_527, C2V_92_639, C2V_92_700, C2V_92_820, C2V_92_910, C2V_92_925, C2V_92_1004, C2V_92_1036, C2V_92_1103, C2V_92_1134, C2V_92_1243, C2V_92_1244, C2V_93_24, C2V_93_51, C2V_93_116, C2V_93_150, C2V_93_216, C2V_93_283, C2V_93_380, C2V_93_387, C2V_93_546, C2V_93_603, C2V_93_631, C2V_93_735, C2V_93_866, C2V_93_958, C2V_93_983, C2V_93_1043, C2V_93_1073, C2V_93_1118, C2V_93_1244, C2V_93_1245, C2V_94_43, C2V_94_54, C2V_94_141, C2V_94_149, C2V_94_214, C2V_94_268, C2V_94_444, C2V_94_484, C2V_94_568, C2V_94_582, C2V_94_655, C2V_94_701, C2V_94_870, C2V_94_942, C2V_94_978, C2V_94_1056, C2V_94_1083, C2V_94_1147, C2V_94_1245, C2V_94_1246, C2V_95_14, C2V_95_72, C2V_95_107, C2V_95_178, C2V_95_194, C2V_95_260, C2V_95_309, C2V_95_376, C2V_95_455, C2V_95_689, C2V_95_753, C2V_95_807, C2V_95_885, C2V_95_933, C2V_95_976, C2V_95_1028, C2V_95_1077, C2V_95_1125, C2V_95_1246, C2V_95_1247, C2V_96_45, C2V_96_69, C2V_96_109, C2V_96_177, C2V_96_211, C2V_96_242, C2V_96_295, C2V_96_447, C2V_96_544, C2V_96_577, C2V_96_781, C2V_96_857, C2V_96_890, C2V_96_952, C2V_96_987, C2V_96_1054, C2V_96_1070, C2V_96_1120, C2V_96_1247, C2V_96_1248, C2V_97_21, C2V_97_57, C2V_97_125, C2V_97_186, C2V_97_200, C2V_97_243, C2V_97_343, C2V_97_397, C2V_97_494, C2V_97_730, C2V_97_778, C2V_97_826, C2V_97_867, C2V_97_956, C2V_97_990, C2V_97_1029, C2V_97_1103, C2V_97_1114, C2V_97_1248, C2V_97_1249, C2V_98_30, C2V_98_79, C2V_98_135, C2V_98_183, C2V_98_212, C2V_98_281, C2V_98_332, C2V_98_391, C2V_98_528, C2V_98_640, C2V_98_701, C2V_98_821, C2V_98_911, C2V_98_926, C2V_98_1005, C2V_98_1037, C2V_98_1104, C2V_98_1135, C2V_98_1249, C2V_98_1250, C2V_99_25, C2V_99_52, C2V_99_117, C2V_99_151, C2V_99_217, C2V_99_284, C2V_99_381, C2V_99_388, C2V_99_547, C2V_99_604, C2V_99_632, C2V_99_736, C2V_99_867, C2V_99_959, C2V_99_984, C2V_99_1044, C2V_99_1074, C2V_99_1119, C2V_99_1250, C2V_99_1251, C2V_100_44, C2V_100_55, C2V_100_142, C2V_100_150, C2V_100_215, C2V_100_269, C2V_100_445, C2V_100_485, C2V_100_569, C2V_100_583, C2V_100_656, C2V_100_702, C2V_100_871, C2V_100_943, C2V_100_979, C2V_100_1009, C2V_100_1084, C2V_100_1148, C2V_100_1251, C2V_100_1252, C2V_101_15, C2V_101_73, C2V_101_108, C2V_101_179, C2V_101_195, C2V_101_261, C2V_101_310, C2V_101_377, C2V_101_456, C2V_101_690, C2V_101_754, C2V_101_808, C2V_101_886, C2V_101_934, C2V_101_977, C2V_101_1029, C2V_101_1078, C2V_101_1126, C2V_101_1252, C2V_101_1253, C2V_102_46, C2V_102_70, C2V_102_110, C2V_102_178, C2V_102_212, C2V_102_243, C2V_102_296, C2V_102_448, C2V_102_545, C2V_102_578, C2V_102_782, C2V_102_858, C2V_102_891, C2V_102_953, C2V_102_988, C2V_102_1055, C2V_102_1071, C2V_102_1121, C2V_102_1253, C2V_102_1254, C2V_103_22, C2V_103_58, C2V_103_126, C2V_103_187, C2V_103_201, C2V_103_244, C2V_103_344, C2V_103_398, C2V_103_495, C2V_103_731, C2V_103_779, C2V_103_827, C2V_103_868, C2V_103_957, C2V_103_991, C2V_103_1030, C2V_103_1104, C2V_103_1115, C2V_103_1254, C2V_103_1255, C2V_104_31, C2V_104_80, C2V_104_136, C2V_104_184, C2V_104_213, C2V_104_282, C2V_104_333, C2V_104_392, C2V_104_481, C2V_104_641, C2V_104_702, C2V_104_822, C2V_104_912, C2V_104_927, C2V_104_1006, C2V_104_1038, C2V_104_1057, C2V_104_1136, C2V_104_1255, C2V_104_1256, C2V_105_26, C2V_105_53, C2V_105_118, C2V_105_152, C2V_105_218, C2V_105_285, C2V_105_382, C2V_105_389, C2V_105_548, C2V_105_605, C2V_105_633, C2V_105_737, C2V_105_868, C2V_105_960, C2V_105_985, C2V_105_1045, C2V_105_1075, C2V_105_1120, C2V_105_1256, C2V_105_1257, C2V_106_45, C2V_106_56, C2V_106_143, C2V_106_151, C2V_106_216, C2V_106_270, C2V_106_446, C2V_106_486, C2V_106_570, C2V_106_584, C2V_106_657, C2V_106_703, C2V_106_872, C2V_106_944, C2V_106_980, C2V_106_1010, C2V_106_1085, C2V_106_1149, C2V_106_1257, C2V_106_1258, C2V_107_16, C2V_107_74, C2V_107_109, C2V_107_180, C2V_107_196, C2V_107_262, C2V_107_311, C2V_107_378, C2V_107_457, C2V_107_691, C2V_107_755, C2V_107_809, C2V_107_887, C2V_107_935, C2V_107_978, C2V_107_1030, C2V_107_1079, C2V_107_1127, C2V_107_1258, C2V_107_1259, C2V_108_47, C2V_108_71, C2V_108_111, C2V_108_179, C2V_108_213, C2V_108_244, C2V_108_297, C2V_108_449, C2V_108_546, C2V_108_579, C2V_108_783, C2V_108_859, C2V_108_892, C2V_108_954, C2V_108_989, C2V_108_1056, C2V_108_1072, C2V_108_1122, C2V_108_1259, C2V_108_1260, C2V_109_23, C2V_109_59, C2V_109_127, C2V_109_188, C2V_109_202, C2V_109_245, C2V_109_345, C2V_109_399, C2V_109_496, C2V_109_732, C2V_109_780, C2V_109_828, C2V_109_869, C2V_109_958, C2V_109_992, C2V_109_1031, C2V_109_1057, C2V_109_1116, C2V_109_1260, C2V_109_1261, C2V_110_32, C2V_110_81, C2V_110_137, C2V_110_185, C2V_110_214, C2V_110_283, C2V_110_334, C2V_110_393, C2V_110_482, C2V_110_642, C2V_110_703, C2V_110_823, C2V_110_865, C2V_110_928, C2V_110_1007, C2V_110_1039, C2V_110_1058, C2V_110_1137, C2V_110_1261, C2V_110_1262, C2V_111_27, C2V_111_54, C2V_111_119, C2V_111_153, C2V_111_219, C2V_111_286, C2V_111_383, C2V_111_390, C2V_111_549, C2V_111_606, C2V_111_634, C2V_111_738, C2V_111_869, C2V_111_913, C2V_111_986, C2V_111_1046, C2V_111_1076, C2V_111_1121, C2V_111_1262, C2V_111_1263, C2V_112_46, C2V_112_57, C2V_112_144, C2V_112_152, C2V_112_217, C2V_112_271, C2V_112_447, C2V_112_487, C2V_112_571, C2V_112_585, C2V_112_658, C2V_112_704, C2V_112_873, C2V_112_945, C2V_112_981, C2V_112_1011, C2V_112_1086, C2V_112_1150, C2V_112_1263, C2V_112_1264, C2V_113_17, C2V_113_75, C2V_113_110, C2V_113_181, C2V_113_197, C2V_113_263, C2V_113_312, C2V_113_379, C2V_113_458, C2V_113_692, C2V_113_756, C2V_113_810, C2V_113_888, C2V_113_936, C2V_113_979, C2V_113_1031, C2V_113_1080, C2V_113_1128, C2V_113_1264, C2V_113_1265, C2V_114_48, C2V_114_72, C2V_114_112, C2V_114_180, C2V_114_214, C2V_114_245, C2V_114_298, C2V_114_450, C2V_114_547, C2V_114_580, C2V_114_784, C2V_114_860, C2V_114_893, C2V_114_955, C2V_114_990, C2V_114_1009, C2V_114_1073, C2V_114_1123, C2V_114_1265, C2V_114_1266, C2V_115_24, C2V_115_60, C2V_115_128, C2V_115_189, C2V_115_203, C2V_115_246, C2V_115_346, C2V_115_400, C2V_115_497, C2V_115_733, C2V_115_781, C2V_115_829, C2V_115_870, C2V_115_959, C2V_115_993, C2V_115_1032, C2V_115_1058, C2V_115_1117, C2V_115_1266, C2V_115_1267, C2V_116_33, C2V_116_82, C2V_116_138, C2V_116_186, C2V_116_215, C2V_116_284, C2V_116_335, C2V_116_394, C2V_116_483, C2V_116_643, C2V_116_704, C2V_116_824, C2V_116_866, C2V_116_929, C2V_116_1008, C2V_116_1040, C2V_116_1059, C2V_116_1138, C2V_116_1267, C2V_116_1268, C2V_117_28, C2V_117_55, C2V_117_120, C2V_117_154, C2V_117_220, C2V_117_287, C2V_117_384, C2V_117_391, C2V_117_550, C2V_117_607, C2V_117_635, C2V_117_739, C2V_117_870, C2V_117_914, C2V_117_987, C2V_117_1047, C2V_117_1077, C2V_117_1122, C2V_117_1268, C2V_117_1269, C2V_118_47, C2V_118_58, C2V_118_97, C2V_118_153, C2V_118_218, C2V_118_272, C2V_118_448, C2V_118_488, C2V_118_572, C2V_118_586, C2V_118_659, C2V_118_705, C2V_118_874, C2V_118_946, C2V_118_982, C2V_118_1012, C2V_118_1087, C2V_118_1151, C2V_118_1269, C2V_118_1270, C2V_119_18, C2V_119_76, C2V_119_111, C2V_119_182, C2V_119_198, C2V_119_264, C2V_119_313, C2V_119_380, C2V_119_459, C2V_119_693, C2V_119_757, C2V_119_811, C2V_119_889, C2V_119_937, C2V_119_980, C2V_119_1032, C2V_119_1081, C2V_119_1129, C2V_119_1270, C2V_119_1271, C2V_120_1, C2V_120_73, C2V_120_113, C2V_120_181, C2V_120_215, C2V_120_246, C2V_120_299, C2V_120_451, C2V_120_548, C2V_120_581, C2V_120_785, C2V_120_861, C2V_120_894, C2V_120_956, C2V_120_991, C2V_120_1010, C2V_120_1074, C2V_120_1124, C2V_120_1271, C2V_120_1272, C2V_121_25, C2V_121_61, C2V_121_129, C2V_121_190, C2V_121_204, C2V_121_247, C2V_121_347, C2V_121_401, C2V_121_498, C2V_121_734, C2V_121_782, C2V_121_830, C2V_121_871, C2V_121_960, C2V_121_994, C2V_121_1033, C2V_121_1059, C2V_121_1118, C2V_121_1272, C2V_121_1273, C2V_122_34, C2V_122_83, C2V_122_139, C2V_122_187, C2V_122_216, C2V_122_285, C2V_122_336, C2V_122_395, C2V_122_484, C2V_122_644, C2V_122_705, C2V_122_825, C2V_122_867, C2V_122_930, C2V_122_961, C2V_122_1041, C2V_122_1060, C2V_122_1139, C2V_122_1273, C2V_122_1274, C2V_123_29, C2V_123_56, C2V_123_121, C2V_123_155, C2V_123_221, C2V_123_288, C2V_123_337, C2V_123_392, C2V_123_551, C2V_123_608, C2V_123_636, C2V_123_740, C2V_123_871, C2V_123_915, C2V_123_988, C2V_123_1048, C2V_123_1078, C2V_123_1123, C2V_123_1274, C2V_123_1275, C2V_124_48, C2V_124_59, C2V_124_98, C2V_124_154, C2V_124_219, C2V_124_273, C2V_124_449, C2V_124_489, C2V_124_573, C2V_124_587, C2V_124_660, C2V_124_706, C2V_124_875, C2V_124_947, C2V_124_983, C2V_124_1013, C2V_124_1088, C2V_124_1152, C2V_124_1275, C2V_124_1276, C2V_125_19, C2V_125_77, C2V_125_112, C2V_125_183, C2V_125_199, C2V_125_265, C2V_125_314, C2V_125_381, C2V_125_460, C2V_125_694, C2V_125_758, C2V_125_812, C2V_125_890, C2V_125_938, C2V_125_981, C2V_125_1033, C2V_125_1082, C2V_125_1130, C2V_125_1276, C2V_125_1277, C2V_126_2, C2V_126_74, C2V_126_114, C2V_126_182, C2V_126_216, C2V_126_247, C2V_126_300, C2V_126_452, C2V_126_549, C2V_126_582, C2V_126_786, C2V_126_862, C2V_126_895, C2V_126_957, C2V_126_992, C2V_126_1011, C2V_126_1075, C2V_126_1125, C2V_126_1277, C2V_126_1278, C2V_127_26, C2V_127_62, C2V_127_130, C2V_127_191, C2V_127_205, C2V_127_248, C2V_127_348, C2V_127_402, C2V_127_499, C2V_127_735, C2V_127_783, C2V_127_831, C2V_127_872, C2V_127_913, C2V_127_995, C2V_127_1034, C2V_127_1060, C2V_127_1119, C2V_127_1278, C2V_127_1279, C2V_128_35, C2V_128_84, C2V_128_140, C2V_128_188, C2V_128_217, C2V_128_286, C2V_128_289, C2V_128_396, C2V_128_485, C2V_128_645, C2V_128_706, C2V_128_826, C2V_128_868, C2V_128_931, C2V_128_962, C2V_128_1042, C2V_128_1061, C2V_128_1140, C2V_128_1279, C2V_128_1280, C2V_129_30, C2V_129_57, C2V_129_122, C2V_129_156, C2V_129_222, C2V_129_241, C2V_129_338, C2V_129_393, C2V_129_552, C2V_129_609, C2V_129_637, C2V_129_741, C2V_129_872, C2V_129_916, C2V_129_989, C2V_129_1049, C2V_129_1079, C2V_129_1124, C2V_129_1280, C2V_129_1281, C2V_130_1, C2V_130_60, C2V_130_99, C2V_130_155, C2V_130_220, C2V_130_274, C2V_130_450, C2V_130_490, C2V_130_574, C2V_130_588, C2V_130_661, C2V_130_707, C2V_130_876, C2V_130_948, C2V_130_984, C2V_130_1014, C2V_130_1089, C2V_130_1105, C2V_130_1281, C2V_130_1282, C2V_131_20, C2V_131_78, C2V_131_113, C2V_131_184, C2V_131_200, C2V_131_266, C2V_131_315, C2V_131_382, C2V_131_461, C2V_131_695, C2V_131_759, C2V_131_813, C2V_131_891, C2V_131_939, C2V_131_982, C2V_131_1034, C2V_131_1083, C2V_131_1131, C2V_131_1282, C2V_131_1283, C2V_132_3, C2V_132_75, C2V_132_115, C2V_132_183, C2V_132_217, C2V_132_248, C2V_132_301, C2V_132_453, C2V_132_550, C2V_132_583, C2V_132_787, C2V_132_863, C2V_132_896, C2V_132_958, C2V_132_993, C2V_132_1012, C2V_132_1076, C2V_132_1126, C2V_132_1283, C2V_132_1284, C2V_133_27, C2V_133_63, C2V_133_131, C2V_133_192, C2V_133_206, C2V_133_249, C2V_133_349, C2V_133_403, C2V_133_500, C2V_133_736, C2V_133_784, C2V_133_832, C2V_133_873, C2V_133_914, C2V_133_996, C2V_133_1035, C2V_133_1061, C2V_133_1120, C2V_133_1284, C2V_133_1285, C2V_134_36, C2V_134_85, C2V_134_141, C2V_134_189, C2V_134_218, C2V_134_287, C2V_134_290, C2V_134_397, C2V_134_486, C2V_134_646, C2V_134_707, C2V_134_827, C2V_134_869, C2V_134_932, C2V_134_963, C2V_134_1043, C2V_134_1062, C2V_134_1141, C2V_134_1285, C2V_134_1286, C2V_135_31, C2V_135_58, C2V_135_123, C2V_135_157, C2V_135_223, C2V_135_242, C2V_135_339, C2V_135_394, C2V_135_553, C2V_135_610, C2V_135_638, C2V_135_742, C2V_135_873, C2V_135_917, C2V_135_990, C2V_135_1050, C2V_135_1080, C2V_135_1125, C2V_135_1286, C2V_135_1287, C2V_136_2, C2V_136_61, C2V_136_100, C2V_136_156, C2V_136_221, C2V_136_275, C2V_136_451, C2V_136_491, C2V_136_575, C2V_136_589, C2V_136_662, C2V_136_708, C2V_136_877, C2V_136_949, C2V_136_985, C2V_136_1015, C2V_136_1090, C2V_136_1106, C2V_136_1287, C2V_136_1288, C2V_137_21, C2V_137_79, C2V_137_114, C2V_137_185, C2V_137_201, C2V_137_267, C2V_137_316, C2V_137_383, C2V_137_462, C2V_137_696, C2V_137_760, C2V_137_814, C2V_137_892, C2V_137_940, C2V_137_983, C2V_137_1035, C2V_137_1084, C2V_137_1132, C2V_137_1288, C2V_137_1289, C2V_138_4, C2V_138_76, C2V_138_116, C2V_138_184, C2V_138_218, C2V_138_249, C2V_138_302, C2V_138_454, C2V_138_551, C2V_138_584, C2V_138_788, C2V_138_864, C2V_138_897, C2V_138_959, C2V_138_994, C2V_138_1013, C2V_138_1077, C2V_138_1127, C2V_138_1289, C2V_138_1290, C2V_139_28, C2V_139_64, C2V_139_132, C2V_139_145, C2V_139_207, C2V_139_250, C2V_139_350, C2V_139_404, C2V_139_501, C2V_139_737, C2V_139_785, C2V_139_833, C2V_139_874, C2V_139_915, C2V_139_997, C2V_139_1036, C2V_139_1062, C2V_139_1121, C2V_139_1290, C2V_139_1291, C2V_140_37, C2V_140_86, C2V_140_142, C2V_140_190, C2V_140_219, C2V_140_288, C2V_140_291, C2V_140_398, C2V_140_487, C2V_140_647, C2V_140_708, C2V_140_828, C2V_140_870, C2V_140_933, C2V_140_964, C2V_140_1044, C2V_140_1063, C2V_140_1142, C2V_140_1291, C2V_140_1292, C2V_141_32, C2V_141_59, C2V_141_124, C2V_141_158, C2V_141_224, C2V_141_243, C2V_141_340, C2V_141_395, C2V_141_554, C2V_141_611, C2V_141_639, C2V_141_743, C2V_141_874, C2V_141_918, C2V_141_991, C2V_141_1051, C2V_141_1081, C2V_141_1126, C2V_141_1292, C2V_141_1293, C2V_142_3, C2V_142_62, C2V_142_101, C2V_142_157, C2V_142_222, C2V_142_276, C2V_142_452, C2V_142_492, C2V_142_576, C2V_142_590, C2V_142_663, C2V_142_709, C2V_142_878, C2V_142_950, C2V_142_986, C2V_142_1016, C2V_142_1091, C2V_142_1107, C2V_142_1293, C2V_142_1294, C2V_143_22, C2V_143_80, C2V_143_115, C2V_143_186, C2V_143_202, C2V_143_268, C2V_143_317, C2V_143_384, C2V_143_463, C2V_143_697, C2V_143_761, C2V_143_815, C2V_143_893, C2V_143_941, C2V_143_984, C2V_143_1036, C2V_143_1085, C2V_143_1133, C2V_143_1294, C2V_143_1295, C2V_144_5, C2V_144_77, C2V_144_117, C2V_144_185, C2V_144_219, C2V_144_250, C2V_144_303, C2V_144_455, C2V_144_552, C2V_144_585, C2V_144_789, C2V_144_817, C2V_144_898, C2V_144_960, C2V_144_995, C2V_144_1014, C2V_144_1078, C2V_144_1128, C2V_144_1295, C2V_144_1296, C2V_145_29, C2V_145_65, C2V_145_133, C2V_145_146, C2V_145_208, C2V_145_251, C2V_145_351, C2V_145_405, C2V_145_502, C2V_145_738, C2V_145_786, C2V_145_834, C2V_145_875, C2V_145_916, C2V_145_998, C2V_145_1037, C2V_145_1063, C2V_145_1122, C2V_145_1296, C2V_145_1297, C2V_146_38, C2V_146_87, C2V_146_143, C2V_146_191, C2V_146_220, C2V_146_241, C2V_146_292, C2V_146_399, C2V_146_488, C2V_146_648, C2V_146_709, C2V_146_829, C2V_146_871, C2V_146_934, C2V_146_965, C2V_146_1045, C2V_146_1064, C2V_146_1143, C2V_146_1297, C2V_146_1298, C2V_147_33, C2V_147_60, C2V_147_125, C2V_147_159, C2V_147_225, C2V_147_244, C2V_147_341, C2V_147_396, C2V_147_555, C2V_147_612, C2V_147_640, C2V_147_744, C2V_147_875, C2V_147_919, C2V_147_992, C2V_147_1052, C2V_147_1082, C2V_147_1127, C2V_147_1298, C2V_147_1299, C2V_148_4, C2V_148_63, C2V_148_102, C2V_148_158, C2V_148_223, C2V_148_277, C2V_148_453, C2V_148_493, C2V_148_529, C2V_148_591, C2V_148_664, C2V_148_710, C2V_148_879, C2V_148_951, C2V_148_987, C2V_148_1017, C2V_148_1092, C2V_148_1108, C2V_148_1299, C2V_148_1300, C2V_149_23, C2V_149_81, C2V_149_116, C2V_149_187, C2V_149_203, C2V_149_269, C2V_149_318, C2V_149_337, C2V_149_464, C2V_149_698, C2V_149_762, C2V_149_816, C2V_149_894, C2V_149_942, C2V_149_985, C2V_149_1037, C2V_149_1086, C2V_149_1134, C2V_149_1300, C2V_149_1301, C2V_150_6, C2V_150_78, C2V_150_118, C2V_150_186, C2V_150_220, C2V_150_251, C2V_150_304, C2V_150_456, C2V_150_553, C2V_150_586, C2V_150_790, C2V_150_818, C2V_150_899, C2V_150_913, C2V_150_996, C2V_150_1015, C2V_150_1079, C2V_150_1129, C2V_150_1301, C2V_150_1302, C2V_151_30, C2V_151_66, C2V_151_134, C2V_151_147, C2V_151_209, C2V_151_252, C2V_151_352, C2V_151_406, C2V_151_503, C2V_151_739, C2V_151_787, C2V_151_835, C2V_151_876, C2V_151_917, C2V_151_999, C2V_151_1038, C2V_151_1064, C2V_151_1123, C2V_151_1302, C2V_151_1303, C2V_152_39, C2V_152_88, C2V_152_144, C2V_152_192, C2V_152_221, C2V_152_242, C2V_152_293, C2V_152_400, C2V_152_489, C2V_152_649, C2V_152_710, C2V_152_830, C2V_152_872, C2V_152_935, C2V_152_966, C2V_152_1046, C2V_152_1065, C2V_152_1144, C2V_152_1303, C2V_152_1304, C2V_153_34, C2V_153_61, C2V_153_126, C2V_153_160, C2V_153_226, C2V_153_245, C2V_153_342, C2V_153_397, C2V_153_556, C2V_153_613, C2V_153_641, C2V_153_745, C2V_153_876, C2V_153_920, C2V_153_993, C2V_153_1053, C2V_153_1083, C2V_153_1128, C2V_153_1304, C2V_153_1305, C2V_154_5, C2V_154_64, C2V_154_103, C2V_154_159, C2V_154_224, C2V_154_278, C2V_154_454, C2V_154_494, C2V_154_530, C2V_154_592, C2V_154_665, C2V_154_711, C2V_154_880, C2V_154_952, C2V_154_988, C2V_154_1018, C2V_154_1093, C2V_154_1109, C2V_154_1305, C2V_154_1306, C2V_155_24, C2V_155_82, C2V_155_117, C2V_155_188, C2V_155_204, C2V_155_270, C2V_155_319, C2V_155_338, C2V_155_465, C2V_155_699, C2V_155_763, C2V_155_769, C2V_155_895, C2V_155_943, C2V_155_986, C2V_155_1038, C2V_155_1087, C2V_155_1135, C2V_155_1306, C2V_155_1307, C2V_156_7, C2V_156_79, C2V_156_119, C2V_156_187, C2V_156_221, C2V_156_252, C2V_156_305, C2V_156_457, C2V_156_554, C2V_156_587, C2V_156_791, C2V_156_819, C2V_156_900, C2V_156_914, C2V_156_997, C2V_156_1016, C2V_156_1080, C2V_156_1130, C2V_156_1307, C2V_156_1308, C2V_157_31, C2V_157_67, C2V_157_135, C2V_157_148, C2V_157_210, C2V_157_253, C2V_157_353, C2V_157_407, C2V_157_504, C2V_157_740, C2V_157_788, C2V_157_836, C2V_157_877, C2V_157_918, C2V_157_1000, C2V_157_1039, C2V_157_1065, C2V_157_1124, C2V_157_1308, C2V_157_1309, C2V_158_40, C2V_158_89, C2V_158_97, C2V_158_145, C2V_158_222, C2V_158_243, C2V_158_294, C2V_158_401, C2V_158_490, C2V_158_650, C2V_158_711, C2V_158_831, C2V_158_873, C2V_158_936, C2V_158_967, C2V_158_1047, C2V_158_1066, C2V_158_1145, C2V_158_1309, C2V_158_1310, C2V_159_35, C2V_159_62, C2V_159_127, C2V_159_161, C2V_159_227, C2V_159_246, C2V_159_343, C2V_159_398, C2V_159_557, C2V_159_614, C2V_159_642, C2V_159_746, C2V_159_877, C2V_159_921, C2V_159_994, C2V_159_1054, C2V_159_1084, C2V_159_1129, C2V_159_1310, C2V_159_1311, C2V_160_6, C2V_160_65, C2V_160_104, C2V_160_160, C2V_160_225, C2V_160_279, C2V_160_455, C2V_160_495, C2V_160_531, C2V_160_593, C2V_160_666, C2V_160_712, C2V_160_881, C2V_160_953, C2V_160_989, C2V_160_1019, C2V_160_1094, C2V_160_1110, C2V_160_1311, C2V_160_1312, C2V_161_25, C2V_161_83, C2V_161_118, C2V_161_189, C2V_161_205, C2V_161_271, C2V_161_320, C2V_161_339, C2V_161_466, C2V_161_700, C2V_161_764, C2V_161_770, C2V_161_896, C2V_161_944, C2V_161_987, C2V_161_1039, C2V_161_1088, C2V_161_1136, C2V_161_1312, C2V_161_1313, C2V_162_8, C2V_162_80, C2V_162_120, C2V_162_188, C2V_162_222, C2V_162_253, C2V_162_306, C2V_162_458, C2V_162_555, C2V_162_588, C2V_162_792, C2V_162_820, C2V_162_901, C2V_162_915, C2V_162_998, C2V_162_1017, C2V_162_1081, C2V_162_1131, C2V_162_1313, C2V_162_1314, C2V_163_32, C2V_163_68, C2V_163_136, C2V_163_149, C2V_163_211, C2V_163_254, C2V_163_354, C2V_163_408, C2V_163_505, C2V_163_741, C2V_163_789, C2V_163_837, C2V_163_878, C2V_163_919, C2V_163_1001, C2V_163_1040, C2V_163_1066, C2V_163_1125, C2V_163_1314, C2V_163_1315, C2V_164_41, C2V_164_90, C2V_164_98, C2V_164_146, C2V_164_223, C2V_164_244, C2V_164_295, C2V_164_402, C2V_164_491, C2V_164_651, C2V_164_712, C2V_164_832, C2V_164_874, C2V_164_937, C2V_164_968, C2V_164_1048, C2V_164_1067, C2V_164_1146, C2V_164_1315, C2V_164_1316, C2V_165_36, C2V_165_63, C2V_165_128, C2V_165_162, C2V_165_228, C2V_165_247, C2V_165_344, C2V_165_399, C2V_165_558, C2V_165_615, C2V_165_643, C2V_165_747, C2V_165_878, C2V_165_922, C2V_165_995, C2V_165_1055, C2V_165_1085, C2V_165_1130, C2V_165_1316, C2V_165_1317, C2V_166_7, C2V_166_66, C2V_166_105, C2V_166_161, C2V_166_226, C2V_166_280, C2V_166_456, C2V_166_496, C2V_166_532, C2V_166_594, C2V_166_667, C2V_166_713, C2V_166_882, C2V_166_954, C2V_166_990, C2V_166_1020, C2V_166_1095, C2V_166_1111, C2V_166_1317, C2V_166_1318, C2V_167_26, C2V_167_84, C2V_167_119, C2V_167_190, C2V_167_206, C2V_167_272, C2V_167_321, C2V_167_340, C2V_167_467, C2V_167_701, C2V_167_765, C2V_167_771, C2V_167_897, C2V_167_945, C2V_167_988, C2V_167_1040, C2V_167_1089, C2V_167_1137, C2V_167_1318, C2V_167_1319, C2V_168_9, C2V_168_81, C2V_168_121, C2V_168_189, C2V_168_223, C2V_168_254, C2V_168_307, C2V_168_459, C2V_168_556, C2V_168_589, C2V_168_793, C2V_168_821, C2V_168_902, C2V_168_916, C2V_168_999, C2V_168_1018, C2V_168_1082, C2V_168_1132, C2V_168_1319, C2V_168_1320, C2V_169_33, C2V_169_69, C2V_169_137, C2V_169_150, C2V_169_212, C2V_169_255, C2V_169_355, C2V_169_409, C2V_169_506, C2V_169_742, C2V_169_790, C2V_169_838, C2V_169_879, C2V_169_920, C2V_169_1002, C2V_169_1041, C2V_169_1067, C2V_169_1126, C2V_169_1320, C2V_169_1321, C2V_170_42, C2V_170_91, C2V_170_99, C2V_170_147, C2V_170_224, C2V_170_245, C2V_170_296, C2V_170_403, C2V_170_492, C2V_170_652, C2V_170_713, C2V_170_833, C2V_170_875, C2V_170_938, C2V_170_969, C2V_170_1049, C2V_170_1068, C2V_170_1147, C2V_170_1321, C2V_170_1322, C2V_171_37, C2V_171_64, C2V_171_129, C2V_171_163, C2V_171_229, C2V_171_248, C2V_171_345, C2V_171_400, C2V_171_559, C2V_171_616, C2V_171_644, C2V_171_748, C2V_171_879, C2V_171_923, C2V_171_996, C2V_171_1056, C2V_171_1086, C2V_171_1131, C2V_171_1322, C2V_171_1323, C2V_172_8, C2V_172_67, C2V_172_106, C2V_172_162, C2V_172_227, C2V_172_281, C2V_172_457, C2V_172_497, C2V_172_533, C2V_172_595, C2V_172_668, C2V_172_714, C2V_172_883, C2V_172_955, C2V_172_991, C2V_172_1021, C2V_172_1096, C2V_172_1112, C2V_172_1323, C2V_172_1324, C2V_173_27, C2V_173_85, C2V_173_120, C2V_173_191, C2V_173_207, C2V_173_273, C2V_173_322, C2V_173_341, C2V_173_468, C2V_173_702, C2V_173_766, C2V_173_772, C2V_173_898, C2V_173_946, C2V_173_989, C2V_173_1041, C2V_173_1090, C2V_173_1138, C2V_173_1324, C2V_173_1325, C2V_174_10, C2V_174_82, C2V_174_122, C2V_174_190, C2V_174_224, C2V_174_255, C2V_174_308, C2V_174_460, C2V_174_557, C2V_174_590, C2V_174_794, C2V_174_822, C2V_174_903, C2V_174_917, C2V_174_1000, C2V_174_1019, C2V_174_1083, C2V_174_1133, C2V_174_1325, C2V_174_1326, C2V_175_34, C2V_175_70, C2V_175_138, C2V_175_151, C2V_175_213, C2V_175_256, C2V_175_356, C2V_175_410, C2V_175_507, C2V_175_743, C2V_175_791, C2V_175_839, C2V_175_880, C2V_175_921, C2V_175_1003, C2V_175_1042, C2V_175_1068, C2V_175_1127, C2V_175_1326, C2V_175_1327, C2V_176_43, C2V_176_92, C2V_176_100, C2V_176_148, C2V_176_225, C2V_176_246, C2V_176_297, C2V_176_404, C2V_176_493, C2V_176_653, C2V_176_714, C2V_176_834, C2V_176_876, C2V_176_939, C2V_176_970, C2V_176_1050, C2V_176_1069, C2V_176_1148, C2V_176_1327, C2V_176_1328, C2V_177_38, C2V_177_65, C2V_177_130, C2V_177_164, C2V_177_230, C2V_177_249, C2V_177_346, C2V_177_401, C2V_177_560, C2V_177_617, C2V_177_645, C2V_177_749, C2V_177_880, C2V_177_924, C2V_177_997, C2V_177_1009, C2V_177_1087, C2V_177_1132, C2V_177_1328, C2V_177_1329, C2V_178_9, C2V_178_68, C2V_178_107, C2V_178_163, C2V_178_228, C2V_178_282, C2V_178_458, C2V_178_498, C2V_178_534, C2V_178_596, C2V_178_669, C2V_178_715, C2V_178_884, C2V_178_956, C2V_178_992, C2V_178_1022, C2V_178_1097, C2V_178_1113, C2V_178_1329, C2V_178_1330, C2V_179_28, C2V_179_86, C2V_179_121, C2V_179_192, C2V_179_208, C2V_179_274, C2V_179_323, C2V_179_342, C2V_179_469, C2V_179_703, C2V_179_767, C2V_179_773, C2V_179_899, C2V_179_947, C2V_179_990, C2V_179_1042, C2V_179_1091, C2V_179_1139, C2V_179_1330, C2V_179_1331, C2V_180_11, C2V_180_83, C2V_180_123, C2V_180_191, C2V_180_225, C2V_180_256, C2V_180_309, C2V_180_461, C2V_180_558, C2V_180_591, C2V_180_795, C2V_180_823, C2V_180_904, C2V_180_918, C2V_180_1001, C2V_180_1020, C2V_180_1084, C2V_180_1134, C2V_180_1331, C2V_180_1332, C2V_181_35, C2V_181_71, C2V_181_139, C2V_181_152, C2V_181_214, C2V_181_257, C2V_181_357, C2V_181_411, C2V_181_508, C2V_181_744, C2V_181_792, C2V_181_840, C2V_181_881, C2V_181_922, C2V_181_1004, C2V_181_1043, C2V_181_1069, C2V_181_1128, C2V_181_1332, C2V_181_1333, C2V_182_44, C2V_182_93, C2V_182_101, C2V_182_149, C2V_182_226, C2V_182_247, C2V_182_298, C2V_182_405, C2V_182_494, C2V_182_654, C2V_182_715, C2V_182_835, C2V_182_877, C2V_182_940, C2V_182_971, C2V_182_1051, C2V_182_1070, C2V_182_1149, C2V_182_1333, C2V_182_1334, C2V_183_39, C2V_183_66, C2V_183_131, C2V_183_165, C2V_183_231, C2V_183_250, C2V_183_347, C2V_183_402, C2V_183_561, C2V_183_618, C2V_183_646, C2V_183_750, C2V_183_881, C2V_183_925, C2V_183_998, C2V_183_1010, C2V_183_1088, C2V_183_1133, C2V_183_1334, C2V_183_1335, C2V_184_10, C2V_184_69, C2V_184_108, C2V_184_164, C2V_184_229, C2V_184_283, C2V_184_459, C2V_184_499, C2V_184_535, C2V_184_597, C2V_184_670, C2V_184_716, C2V_184_885, C2V_184_957, C2V_184_993, C2V_184_1023, C2V_184_1098, C2V_184_1114, C2V_184_1335, C2V_184_1336, C2V_185_29, C2V_185_87, C2V_185_122, C2V_185_145, C2V_185_209, C2V_185_275, C2V_185_324, C2V_185_343, C2V_185_470, C2V_185_704, C2V_185_768, C2V_185_774, C2V_185_900, C2V_185_948, C2V_185_991, C2V_185_1043, C2V_185_1092, C2V_185_1140, C2V_185_1336, C2V_185_1337, C2V_186_12, C2V_186_84, C2V_186_124, C2V_186_192, C2V_186_226, C2V_186_257, C2V_186_310, C2V_186_462, C2V_186_559, C2V_186_592, C2V_186_796, C2V_186_824, C2V_186_905, C2V_186_919, C2V_186_1002, C2V_186_1021, C2V_186_1085, C2V_186_1135, C2V_186_1337, C2V_186_1338, C2V_187_36, C2V_187_72, C2V_187_140, C2V_187_153, C2V_187_215, C2V_187_258, C2V_187_358, C2V_187_412, C2V_187_509, C2V_187_745, C2V_187_793, C2V_187_841, C2V_187_882, C2V_187_923, C2V_187_1005, C2V_187_1044, C2V_187_1070, C2V_187_1129, C2V_187_1338, C2V_187_1339, C2V_188_45, C2V_188_94, C2V_188_102, C2V_188_150, C2V_188_227, C2V_188_248, C2V_188_299, C2V_188_406, C2V_188_495, C2V_188_655, C2V_188_716, C2V_188_836, C2V_188_878, C2V_188_941, C2V_188_972, C2V_188_1052, C2V_188_1071, C2V_188_1150, C2V_188_1339, C2V_188_1340, C2V_189_40, C2V_189_67, C2V_189_132, C2V_189_166, C2V_189_232, C2V_189_251, C2V_189_348, C2V_189_403, C2V_189_562, C2V_189_619, C2V_189_647, C2V_189_751, C2V_189_882, C2V_189_926, C2V_189_999, C2V_189_1011, C2V_189_1089, C2V_189_1134, C2V_189_1340, C2V_189_1341, C2V_190_11, C2V_190_70, C2V_190_109, C2V_190_165, C2V_190_230, C2V_190_284, C2V_190_460, C2V_190_500, C2V_190_536, C2V_190_598, C2V_190_671, C2V_190_717, C2V_190_886, C2V_190_958, C2V_190_994, C2V_190_1024, C2V_190_1099, C2V_190_1115, C2V_190_1341, C2V_190_1342, C2V_191_30, C2V_191_88, C2V_191_123, C2V_191_146, C2V_191_210, C2V_191_276, C2V_191_325, C2V_191_344, C2V_191_471, C2V_191_705, C2V_191_721, C2V_191_775, C2V_191_901, C2V_191_949, C2V_191_992, C2V_191_1044, C2V_191_1093, C2V_191_1141, C2V_191_1342, C2V_191_1343, C2V_192_13, C2V_192_85, C2V_192_125, C2V_192_145, C2V_192_227, C2V_192_258, C2V_192_311, C2V_192_463, C2V_192_560, C2V_192_593, C2V_192_797, C2V_192_825, C2V_192_906, C2V_192_920, C2V_192_1003, C2V_192_1022, C2V_192_1086, C2V_192_1136, C2V_192_1343, C2V_192_1344, C2V_193_37, C2V_193_73, C2V_193_141, C2V_193_154, C2V_193_216, C2V_193_259, C2V_193_359, C2V_193_413, C2V_193_510, C2V_193_746, C2V_193_794, C2V_193_842, C2V_193_883, C2V_193_924, C2V_193_1006, C2V_193_1045, C2V_193_1071, C2V_193_1130, C2V_193_1344, C2V_193_1345, C2V_194_46, C2V_194_95, C2V_194_103, C2V_194_151, C2V_194_228, C2V_194_249, C2V_194_300, C2V_194_407, C2V_194_496, C2V_194_656, C2V_194_717, C2V_194_837, C2V_194_879, C2V_194_942, C2V_194_973, C2V_194_1053, C2V_194_1072, C2V_194_1151, C2V_194_1345, C2V_194_1346, C2V_195_41, C2V_195_68, C2V_195_133, C2V_195_167, C2V_195_233, C2V_195_252, C2V_195_349, C2V_195_404, C2V_195_563, C2V_195_620, C2V_195_648, C2V_195_752, C2V_195_883, C2V_195_927, C2V_195_1000, C2V_195_1012, C2V_195_1090, C2V_195_1135, C2V_195_1346, C2V_195_1347, C2V_196_12, C2V_196_71, C2V_196_110, C2V_196_166, C2V_196_231, C2V_196_285, C2V_196_461, C2V_196_501, C2V_196_537, C2V_196_599, C2V_196_672, C2V_196_718, C2V_196_887, C2V_196_959, C2V_196_995, C2V_196_1025, C2V_196_1100, C2V_196_1116, C2V_196_1347, C2V_196_1348, C2V_197_31, C2V_197_89, C2V_197_124, C2V_197_147, C2V_197_211, C2V_197_277, C2V_197_326, C2V_197_345, C2V_197_472, C2V_197_706, C2V_197_722, C2V_197_776, C2V_197_902, C2V_197_950, C2V_197_993, C2V_197_1045, C2V_197_1094, C2V_197_1142, C2V_197_1348, C2V_197_1349, C2V_198_14, C2V_198_86, C2V_198_126, C2V_198_146, C2V_198_228, C2V_198_259, C2V_198_312, C2V_198_464, C2V_198_561, C2V_198_594, C2V_198_798, C2V_198_826, C2V_198_907, C2V_198_921, C2V_198_1004, C2V_198_1023, C2V_198_1087, C2V_198_1137, C2V_198_1349, C2V_198_1350, C2V_199_38, C2V_199_74, C2V_199_142, C2V_199_155, C2V_199_217, C2V_199_260, C2V_199_360, C2V_199_414, C2V_199_511, C2V_199_747, C2V_199_795, C2V_199_843, C2V_199_884, C2V_199_925, C2V_199_1007, C2V_199_1046, C2V_199_1072, C2V_199_1131, C2V_199_1350, C2V_199_1351, C2V_200_47, C2V_200_96, C2V_200_104, C2V_200_152, C2V_200_229, C2V_200_250, C2V_200_301, C2V_200_408, C2V_200_497, C2V_200_657, C2V_200_718, C2V_200_838, C2V_200_880, C2V_200_943, C2V_200_974, C2V_200_1054, C2V_200_1073, C2V_200_1152, C2V_200_1351, C2V_200_1352, C2V_201_42, C2V_201_69, C2V_201_134, C2V_201_168, C2V_201_234, C2V_201_253, C2V_201_350, C2V_201_405, C2V_201_564, C2V_201_621, C2V_201_649, C2V_201_753, C2V_201_884, C2V_201_928, C2V_201_1001, C2V_201_1013, C2V_201_1091, C2V_201_1136, C2V_201_1352, C2V_201_1353, C2V_202_13, C2V_202_72, C2V_202_111, C2V_202_167, C2V_202_232, C2V_202_286, C2V_202_462, C2V_202_502, C2V_202_538, C2V_202_600, C2V_202_625, C2V_202_719, C2V_202_888, C2V_202_960, C2V_202_996, C2V_202_1026, C2V_202_1101, C2V_202_1117, C2V_202_1353, C2V_202_1354, C2V_203_32, C2V_203_90, C2V_203_125, C2V_203_148, C2V_203_212, C2V_203_278, C2V_203_327, C2V_203_346, C2V_203_473, C2V_203_707, C2V_203_723, C2V_203_777, C2V_203_903, C2V_203_951, C2V_203_994, C2V_203_1046, C2V_203_1095, C2V_203_1143, C2V_203_1354, C2V_203_1355, C2V_204_15, C2V_204_87, C2V_204_127, C2V_204_147, C2V_204_229, C2V_204_260, C2V_204_313, C2V_204_465, C2V_204_562, C2V_204_595, C2V_204_799, C2V_204_827, C2V_204_908, C2V_204_922, C2V_204_1005, C2V_204_1024, C2V_204_1088, C2V_204_1138, C2V_204_1355, C2V_204_1356, C2V_205_39, C2V_205_75, C2V_205_143, C2V_205_156, C2V_205_218, C2V_205_261, C2V_205_361, C2V_205_415, C2V_205_512, C2V_205_748, C2V_205_796, C2V_205_844, C2V_205_885, C2V_205_926, C2V_205_1008, C2V_205_1047, C2V_205_1073, C2V_205_1132, C2V_205_1356, C2V_205_1357, C2V_206_48, C2V_206_49, C2V_206_105, C2V_206_153, C2V_206_230, C2V_206_251, C2V_206_302, C2V_206_409, C2V_206_498, C2V_206_658, C2V_206_719, C2V_206_839, C2V_206_881, C2V_206_944, C2V_206_975, C2V_206_1055, C2V_206_1074, C2V_206_1105, C2V_206_1357, C2V_206_1358, C2V_207_43, C2V_207_70, C2V_207_135, C2V_207_169, C2V_207_235, C2V_207_254, C2V_207_351, C2V_207_406, C2V_207_565, C2V_207_622, C2V_207_650, C2V_207_754, C2V_207_885, C2V_207_929, C2V_207_1002, C2V_207_1014, C2V_207_1092, C2V_207_1137, C2V_207_1358, C2V_207_1359, C2V_208_14, C2V_208_73, C2V_208_112, C2V_208_168, C2V_208_233, C2V_208_287, C2V_208_463, C2V_208_503, C2V_208_539, C2V_208_601, C2V_208_626, C2V_208_720, C2V_208_889, C2V_208_913, C2V_208_997, C2V_208_1027, C2V_208_1102, C2V_208_1118, C2V_208_1359, C2V_208_1360, C2V_209_33, C2V_209_91, C2V_209_126, C2V_209_149, C2V_209_213, C2V_209_279, C2V_209_328, C2V_209_347, C2V_209_474, C2V_209_708, C2V_209_724, C2V_209_778, C2V_209_904, C2V_209_952, C2V_209_995, C2V_209_1047, C2V_209_1096, C2V_209_1144, C2V_209_1360, C2V_209_1361, C2V_210_16, C2V_210_88, C2V_210_128, C2V_210_148, C2V_210_230, C2V_210_261, C2V_210_314, C2V_210_466, C2V_210_563, C2V_210_596, C2V_210_800, C2V_210_828, C2V_210_909, C2V_210_923, C2V_210_1006, C2V_210_1025, C2V_210_1089, C2V_210_1139, C2V_210_1361, C2V_210_1362, C2V_211_40, C2V_211_76, C2V_211_144, C2V_211_157, C2V_211_219, C2V_211_262, C2V_211_362, C2V_211_416, C2V_211_513, C2V_211_749, C2V_211_797, C2V_211_845, C2V_211_886, C2V_211_927, C2V_211_961, C2V_211_1048, C2V_211_1074, C2V_211_1133, C2V_211_1362, C2V_211_1363, C2V_212_1, C2V_212_50, C2V_212_106, C2V_212_154, C2V_212_231, C2V_212_252, C2V_212_303, C2V_212_410, C2V_212_499, C2V_212_659, C2V_212_720, C2V_212_840, C2V_212_882, C2V_212_945, C2V_212_976, C2V_212_1056, C2V_212_1075, C2V_212_1106, C2V_212_1363, C2V_212_1364, C2V_213_44, C2V_213_71, C2V_213_136, C2V_213_170, C2V_213_236, C2V_213_255, C2V_213_352, C2V_213_407, C2V_213_566, C2V_213_623, C2V_213_651, C2V_213_755, C2V_213_886, C2V_213_930, C2V_213_1003, C2V_213_1015, C2V_213_1093, C2V_213_1138, C2V_213_1364, C2V_213_1365, C2V_214_15, C2V_214_74, C2V_214_113, C2V_214_169, C2V_214_234, C2V_214_288, C2V_214_464, C2V_214_504, C2V_214_540, C2V_214_602, C2V_214_627, C2V_214_673, C2V_214_890, C2V_214_914, C2V_214_998, C2V_214_1028, C2V_214_1103, C2V_214_1119, C2V_214_1365, C2V_214_1366, C2V_215_34, C2V_215_92, C2V_215_127, C2V_215_150, C2V_215_214, C2V_215_280, C2V_215_329, C2V_215_348, C2V_215_475, C2V_215_709, C2V_215_725, C2V_215_779, C2V_215_905, C2V_215_953, C2V_215_996, C2V_215_1048, C2V_215_1097, C2V_215_1145, C2V_215_1366, C2V_215_1367, C2V_216_17, C2V_216_89, C2V_216_129, C2V_216_149, C2V_216_231, C2V_216_262, C2V_216_315, C2V_216_467, C2V_216_564, C2V_216_597, C2V_216_801, C2V_216_829, C2V_216_910, C2V_216_924, C2V_216_1007, C2V_216_1026, C2V_216_1090, C2V_216_1140, C2V_216_1367, C2V_216_1368, C2V_217_41, C2V_217_77, C2V_217_97, C2V_217_158, C2V_217_220, C2V_217_263, C2V_217_363, C2V_217_417, C2V_217_514, C2V_217_750, C2V_217_798, C2V_217_846, C2V_217_887, C2V_217_928, C2V_217_962, C2V_217_1049, C2V_217_1075, C2V_217_1134, C2V_217_1368, C2V_217_1369, C2V_218_2, C2V_218_51, C2V_218_107, C2V_218_155, C2V_218_232, C2V_218_253, C2V_218_304, C2V_218_411, C2V_218_500, C2V_218_660, C2V_218_673, C2V_218_841, C2V_218_883, C2V_218_946, C2V_218_977, C2V_218_1009, C2V_218_1076, C2V_218_1107, C2V_218_1369, C2V_218_1370, C2V_219_45, C2V_219_72, C2V_219_137, C2V_219_171, C2V_219_237, C2V_219_256, C2V_219_353, C2V_219_408, C2V_219_567, C2V_219_624, C2V_219_652, C2V_219_756, C2V_219_887, C2V_219_931, C2V_219_1004, C2V_219_1016, C2V_219_1094, C2V_219_1139, C2V_219_1370, C2V_219_1371, C2V_220_16, C2V_220_75, C2V_220_114, C2V_220_170, C2V_220_235, C2V_220_241, C2V_220_465, C2V_220_505, C2V_220_541, C2V_220_603, C2V_220_628, C2V_220_674, C2V_220_891, C2V_220_915, C2V_220_999, C2V_220_1029, C2V_220_1104, C2V_220_1120, C2V_220_1371, C2V_220_1372, C2V_221_35, C2V_221_93, C2V_221_128, C2V_221_151, C2V_221_215, C2V_221_281, C2V_221_330, C2V_221_349, C2V_221_476, C2V_221_710, C2V_221_726, C2V_221_780, C2V_221_906, C2V_221_954, C2V_221_997, C2V_221_1049, C2V_221_1098, C2V_221_1146, C2V_221_1372, C2V_221_1373, C2V_222_18, C2V_222_90, C2V_222_130, C2V_222_150, C2V_222_232, C2V_222_263, C2V_222_316, C2V_222_468, C2V_222_565, C2V_222_598, C2V_222_802, C2V_222_830, C2V_222_911, C2V_222_925, C2V_222_1008, C2V_222_1027, C2V_222_1091, C2V_222_1141, C2V_222_1373, C2V_222_1374, C2V_223_42, C2V_223_78, C2V_223_98, C2V_223_159, C2V_223_221, C2V_223_264, C2V_223_364, C2V_223_418, C2V_223_515, C2V_223_751, C2V_223_799, C2V_223_847, C2V_223_888, C2V_223_929, C2V_223_963, C2V_223_1050, C2V_223_1076, C2V_223_1135, C2V_223_1374, C2V_223_1375, C2V_224_3, C2V_224_52, C2V_224_108, C2V_224_156, C2V_224_233, C2V_224_254, C2V_224_305, C2V_224_412, C2V_224_501, C2V_224_661, C2V_224_674, C2V_224_842, C2V_224_884, C2V_224_947, C2V_224_978, C2V_224_1010, C2V_224_1077, C2V_224_1108, C2V_224_1375, C2V_224_1376, C2V_225_46, C2V_225_73, C2V_225_138, C2V_225_172, C2V_225_238, C2V_225_257, C2V_225_354, C2V_225_409, C2V_225_568, C2V_225_577, C2V_225_653, C2V_225_757, C2V_225_888, C2V_225_932, C2V_225_1005, C2V_225_1017, C2V_225_1095, C2V_225_1140, C2V_225_1376, C2V_225_1377, C2V_226_17, C2V_226_76, C2V_226_115, C2V_226_171, C2V_226_236, C2V_226_242, C2V_226_466, C2V_226_506, C2V_226_542, C2V_226_604, C2V_226_629, C2V_226_675, C2V_226_892, C2V_226_916, C2V_226_1000, C2V_226_1030, C2V_226_1057, C2V_226_1121, C2V_226_1377, C2V_226_1378, C2V_227_36, C2V_227_94, C2V_227_129, C2V_227_152, C2V_227_216, C2V_227_282, C2V_227_331, C2V_227_350, C2V_227_477, C2V_227_711, C2V_227_727, C2V_227_781, C2V_227_907, C2V_227_955, C2V_227_998, C2V_227_1050, C2V_227_1099, C2V_227_1147, C2V_227_1378, C2V_227_1379, C2V_228_19, C2V_228_91, C2V_228_131, C2V_228_151, C2V_228_233, C2V_228_264, C2V_228_317, C2V_228_469, C2V_228_566, C2V_228_599, C2V_228_803, C2V_228_831, C2V_228_912, C2V_228_926, C2V_228_961, C2V_228_1028, C2V_228_1092, C2V_228_1142, C2V_228_1379, C2V_228_1380, C2V_229_43, C2V_229_79, C2V_229_99, C2V_229_160, C2V_229_222, C2V_229_265, C2V_229_365, C2V_229_419, C2V_229_516, C2V_229_752, C2V_229_800, C2V_229_848, C2V_229_889, C2V_229_930, C2V_229_964, C2V_229_1051, C2V_229_1077, C2V_229_1136, C2V_229_1380, C2V_229_1381, C2V_230_4, C2V_230_53, C2V_230_109, C2V_230_157, C2V_230_234, C2V_230_255, C2V_230_306, C2V_230_413, C2V_230_502, C2V_230_662, C2V_230_675, C2V_230_843, C2V_230_885, C2V_230_948, C2V_230_979, C2V_230_1011, C2V_230_1078, C2V_230_1109, C2V_230_1381, C2V_230_1382, C2V_231_47, C2V_231_74, C2V_231_139, C2V_231_173, C2V_231_239, C2V_231_258, C2V_231_355, C2V_231_410, C2V_231_569, C2V_231_578, C2V_231_654, C2V_231_758, C2V_231_889, C2V_231_933, C2V_231_1006, C2V_231_1018, C2V_231_1096, C2V_231_1141, C2V_231_1382, C2V_231_1383, C2V_232_18, C2V_232_77, C2V_232_116, C2V_232_172, C2V_232_237, C2V_232_243, C2V_232_467, C2V_232_507, C2V_232_543, C2V_232_605, C2V_232_630, C2V_232_676, C2V_232_893, C2V_232_917, C2V_232_1001, C2V_232_1031, C2V_232_1058, C2V_232_1122, C2V_232_1383, C2V_232_1384, C2V_233_37, C2V_233_95, C2V_233_130, C2V_233_153, C2V_233_217, C2V_233_283, C2V_233_332, C2V_233_351, C2V_233_478, C2V_233_712, C2V_233_728, C2V_233_782, C2V_233_908, C2V_233_956, C2V_233_999, C2V_233_1051, C2V_233_1100, C2V_233_1148, C2V_233_1384, C2V_233_1385, C2V_234_20, C2V_234_92, C2V_234_132, C2V_234_152, C2V_234_234, C2V_234_265, C2V_234_318, C2V_234_470, C2V_234_567, C2V_234_600, C2V_234_804, C2V_234_832, C2V_234_865, C2V_234_927, C2V_234_962, C2V_234_1029, C2V_234_1093, C2V_234_1143, C2V_234_1385, C2V_234_1386, C2V_235_44, C2V_235_80, C2V_235_100, C2V_235_161, C2V_235_223, C2V_235_266, C2V_235_366, C2V_235_420, C2V_235_517, C2V_235_753, C2V_235_801, C2V_235_849, C2V_235_890, C2V_235_931, C2V_235_965, C2V_235_1052, C2V_235_1078, C2V_235_1137, C2V_235_1386, C2V_235_1387, C2V_236_5, C2V_236_54, C2V_236_110, C2V_236_158, C2V_236_235, C2V_236_256, C2V_236_307, C2V_236_414, C2V_236_503, C2V_236_663, C2V_236_676, C2V_236_844, C2V_236_886, C2V_236_949, C2V_236_980, C2V_236_1012, C2V_236_1079, C2V_236_1110, C2V_236_1387, C2V_236_1388, C2V_237_48, C2V_237_75, C2V_237_140, C2V_237_174, C2V_237_240, C2V_237_259, C2V_237_356, C2V_237_411, C2V_237_570, C2V_237_579, C2V_237_655, C2V_237_759, C2V_237_890, C2V_237_934, C2V_237_1007, C2V_237_1019, C2V_237_1097, C2V_237_1142, C2V_237_1388, C2V_237_1389, C2V_238_19, C2V_238_78, C2V_238_117, C2V_238_173, C2V_238_238, C2V_238_244, C2V_238_468, C2V_238_508, C2V_238_544, C2V_238_606, C2V_238_631, C2V_238_677, C2V_238_894, C2V_238_918, C2V_238_1002, C2V_238_1032, C2V_238_1059, C2V_238_1123, C2V_238_1389, C2V_238_1390, C2V_239_38, C2V_239_96, C2V_239_131, C2V_239_154, C2V_239_218, C2V_239_284, C2V_239_333, C2V_239_352, C2V_239_479, C2V_239_713, C2V_239_729, C2V_239_783, C2V_239_909, C2V_239_957, C2V_239_1000, C2V_239_1052, C2V_239_1101, C2V_239_1149, C2V_239_1390, C2V_239_1391, C2V_240_21, C2V_240_93, C2V_240_133, C2V_240_153, C2V_240_235, C2V_240_266, C2V_240_319, C2V_240_471, C2V_240_568, C2V_240_601, C2V_240_805, C2V_240_833, C2V_240_866, C2V_240_928, C2V_240_963, C2V_240_1030, C2V_240_1094, C2V_240_1144, C2V_240_1391, C2V_240_1392, C2V_241_45, C2V_241_81, C2V_241_101, C2V_241_162, C2V_241_224, C2V_241_267, C2V_241_367, C2V_241_421, C2V_241_518, C2V_241_754, C2V_241_802, C2V_241_850, C2V_241_891, C2V_241_932, C2V_241_966, C2V_241_1053, C2V_241_1079, C2V_241_1138, C2V_241_1392, C2V_241_1393, C2V_242_6, C2V_242_55, C2V_242_111, C2V_242_159, C2V_242_236, C2V_242_257, C2V_242_308, C2V_242_415, C2V_242_504, C2V_242_664, C2V_242_677, C2V_242_845, C2V_242_887, C2V_242_950, C2V_242_981, C2V_242_1013, C2V_242_1080, C2V_242_1111, C2V_242_1393, C2V_242_1394, C2V_243_1, C2V_243_76, C2V_243_141, C2V_243_175, C2V_243_193, C2V_243_260, C2V_243_357, C2V_243_412, C2V_243_571, C2V_243_580, C2V_243_656, C2V_243_760, C2V_243_891, C2V_243_935, C2V_243_1008, C2V_243_1020, C2V_243_1098, C2V_243_1143, C2V_243_1394, C2V_243_1395, C2V_244_20, C2V_244_79, C2V_244_118, C2V_244_174, C2V_244_239, C2V_244_245, C2V_244_469, C2V_244_509, C2V_244_545, C2V_244_607, C2V_244_632, C2V_244_678, C2V_244_895, C2V_244_919, C2V_244_1003, C2V_244_1033, C2V_244_1060, C2V_244_1124, C2V_244_1395, C2V_244_1396, C2V_245_39, C2V_245_49, C2V_245_132, C2V_245_155, C2V_245_219, C2V_245_285, C2V_245_334, C2V_245_353, C2V_245_480, C2V_245_714, C2V_245_730, C2V_245_784, C2V_245_910, C2V_245_958, C2V_245_1001, C2V_245_1053, C2V_245_1102, C2V_245_1150, C2V_245_1396, C2V_245_1397, C2V_246_22, C2V_246_94, C2V_246_134, C2V_246_154, C2V_246_236, C2V_246_267, C2V_246_320, C2V_246_472, C2V_246_569, C2V_246_602, C2V_246_806, C2V_246_834, C2V_246_867, C2V_246_929, C2V_246_964, C2V_246_1031, C2V_246_1095, C2V_246_1145, C2V_246_1397, C2V_246_1398, C2V_247_46, C2V_247_82, C2V_247_102, C2V_247_163, C2V_247_225, C2V_247_268, C2V_247_368, C2V_247_422, C2V_247_519, C2V_247_755, C2V_247_803, C2V_247_851, C2V_247_892, C2V_247_933, C2V_247_967, C2V_247_1054, C2V_247_1080, C2V_247_1139, C2V_247_1398, C2V_247_1399, C2V_248_7, C2V_248_56, C2V_248_112, C2V_248_160, C2V_248_237, C2V_248_258, C2V_248_309, C2V_248_416, C2V_248_505, C2V_248_665, C2V_248_678, C2V_248_846, C2V_248_888, C2V_248_951, C2V_248_982, C2V_248_1014, C2V_248_1081, C2V_248_1112, C2V_248_1399, C2V_248_1400, C2V_249_2, C2V_249_77, C2V_249_142, C2V_249_176, C2V_249_194, C2V_249_261, C2V_249_358, C2V_249_413, C2V_249_572, C2V_249_581, C2V_249_657, C2V_249_761, C2V_249_892, C2V_249_936, C2V_249_961, C2V_249_1021, C2V_249_1099, C2V_249_1144, C2V_249_1400, C2V_249_1401, C2V_250_21, C2V_250_80, C2V_250_119, C2V_250_175, C2V_250_240, C2V_250_246, C2V_250_470, C2V_250_510, C2V_250_546, C2V_250_608, C2V_250_633, C2V_250_679, C2V_250_896, C2V_250_920, C2V_250_1004, C2V_250_1034, C2V_250_1061, C2V_250_1125, C2V_250_1401, C2V_250_1402, C2V_251_40, C2V_251_50, C2V_251_133, C2V_251_156, C2V_251_220, C2V_251_286, C2V_251_335, C2V_251_354, C2V_251_433, C2V_251_715, C2V_251_731, C2V_251_785, C2V_251_911, C2V_251_959, C2V_251_1002, C2V_251_1054, C2V_251_1103, C2V_251_1151, C2V_251_1402, C2V_251_1403, C2V_252_23, C2V_252_95, C2V_252_135, C2V_252_155, C2V_252_237, C2V_252_268, C2V_252_321, C2V_252_473, C2V_252_570, C2V_252_603, C2V_252_807, C2V_252_835, C2V_252_868, C2V_252_930, C2V_252_965, C2V_252_1032, C2V_252_1096, C2V_252_1146, C2V_252_1403, C2V_252_1404, C2V_253_47, C2V_253_83, C2V_253_103, C2V_253_164, C2V_253_226, C2V_253_269, C2V_253_369, C2V_253_423, C2V_253_520, C2V_253_756, C2V_253_804, C2V_253_852, C2V_253_893, C2V_253_934, C2V_253_968, C2V_253_1055, C2V_253_1081, C2V_253_1140, C2V_253_1404, C2V_253_1405, C2V_254_8, C2V_254_57, C2V_254_113, C2V_254_161, C2V_254_238, C2V_254_259, C2V_254_310, C2V_254_417, C2V_254_506, C2V_254_666, C2V_254_679, C2V_254_847, C2V_254_889, C2V_254_952, C2V_254_983, C2V_254_1015, C2V_254_1082, C2V_254_1113, C2V_254_1405, C2V_254_1406, C2V_255_3, C2V_255_78, C2V_255_143, C2V_255_177, C2V_255_195, C2V_255_262, C2V_255_359, C2V_255_414, C2V_255_573, C2V_255_582, C2V_255_658, C2V_255_762, C2V_255_893, C2V_255_937, C2V_255_962, C2V_255_1022, C2V_255_1100, C2V_255_1145, C2V_255_1406, C2V_255_1407, C2V_256_22, C2V_256_81, C2V_256_120, C2V_256_176, C2V_256_193, C2V_256_247, C2V_256_471, C2V_256_511, C2V_256_547, C2V_256_609, C2V_256_634, C2V_256_680, C2V_256_897, C2V_256_921, C2V_256_1005, C2V_256_1035, C2V_256_1062, C2V_256_1126, C2V_256_1407, C2V_256_1408, C2V_257_41, C2V_257_51, C2V_257_134, C2V_257_157, C2V_257_221, C2V_257_287, C2V_257_336, C2V_257_355, C2V_257_434, C2V_257_716, C2V_257_732, C2V_257_786, C2V_257_912, C2V_257_960, C2V_257_1003, C2V_257_1055, C2V_257_1104, C2V_257_1152, C2V_257_1408, C2V_257_1409, C2V_258_24, C2V_258_96, C2V_258_136, C2V_258_156, C2V_258_238, C2V_258_269, C2V_258_322, C2V_258_474, C2V_258_571, C2V_258_604, C2V_258_808, C2V_258_836, C2V_258_869, C2V_258_931, C2V_258_966, C2V_258_1033, C2V_258_1097, C2V_258_1147, C2V_258_1409, C2V_258_1410, C2V_259_48, C2V_259_84, C2V_259_104, C2V_259_165, C2V_259_227, C2V_259_270, C2V_259_370, C2V_259_424, C2V_259_521, C2V_259_757, C2V_259_805, C2V_259_853, C2V_259_894, C2V_259_935, C2V_259_969, C2V_259_1056, C2V_259_1082, C2V_259_1141, C2V_259_1410, C2V_259_1411, C2V_260_9, C2V_260_58, C2V_260_114, C2V_260_162, C2V_260_239, C2V_260_260, C2V_260_311, C2V_260_418, C2V_260_507, C2V_260_667, C2V_260_680, C2V_260_848, C2V_260_890, C2V_260_953, C2V_260_984, C2V_260_1016, C2V_260_1083, C2V_260_1114, C2V_260_1411, C2V_260_1412, C2V_261_4, C2V_261_79, C2V_261_144, C2V_261_178, C2V_261_196, C2V_261_263, C2V_261_360, C2V_261_415, C2V_261_574, C2V_261_583, C2V_261_659, C2V_261_763, C2V_261_894, C2V_261_938, C2V_261_963, C2V_261_1023, C2V_261_1101, C2V_261_1146, C2V_261_1412, C2V_261_1413, C2V_262_23, C2V_262_82, C2V_262_121, C2V_262_177, C2V_262_194, C2V_262_248, C2V_262_472, C2V_262_512, C2V_262_548, C2V_262_610, C2V_262_635, C2V_262_681, C2V_262_898, C2V_262_922, C2V_262_1006, C2V_262_1036, C2V_262_1063, C2V_262_1127, C2V_262_1413, C2V_262_1414, C2V_263_42, C2V_263_52, C2V_263_135, C2V_263_158, C2V_263_222, C2V_263_288, C2V_263_289, C2V_263_356, C2V_263_435, C2V_263_717, C2V_263_733, C2V_263_787, C2V_263_865, C2V_263_913, C2V_263_1004, C2V_263_1056, C2V_263_1057, C2V_263_1105, C2V_263_1414, C2V_263_1415, C2V_264_25, C2V_264_49, C2V_264_137, C2V_264_157, C2V_264_239, C2V_264_270, C2V_264_323, C2V_264_475, C2V_264_572, C2V_264_605, C2V_264_809, C2V_264_837, C2V_264_870, C2V_264_932, C2V_264_967, C2V_264_1034, C2V_264_1098, C2V_264_1148, C2V_264_1415, C2V_264_1416, C2V_265_1, C2V_265_85, C2V_265_105, C2V_265_166, C2V_265_228, C2V_265_271, C2V_265_371, C2V_265_425, C2V_265_522, C2V_265_758, C2V_265_806, C2V_265_854, C2V_265_895, C2V_265_936, C2V_265_970, C2V_265_1009, C2V_265_1083, C2V_265_1142, C2V_265_1416, C2V_265_1417, C2V_266_10, C2V_266_59, C2V_266_115, C2V_266_163, C2V_266_240, C2V_266_261, C2V_266_312, C2V_266_419, C2V_266_508, C2V_266_668, C2V_266_681, C2V_266_849, C2V_266_891, C2V_266_954, C2V_266_985, C2V_266_1017, C2V_266_1084, C2V_266_1115, C2V_266_1417, C2V_266_1418, C2V_267_5, C2V_267_80, C2V_267_97, C2V_267_179, C2V_267_197, C2V_267_264, C2V_267_361, C2V_267_416, C2V_267_575, C2V_267_584, C2V_267_660, C2V_267_764, C2V_267_895, C2V_267_939, C2V_267_964, C2V_267_1024, C2V_267_1102, C2V_267_1147, C2V_267_1418, C2V_267_1419, C2V_268_24, C2V_268_83, C2V_268_122, C2V_268_178, C2V_268_195, C2V_268_249, C2V_268_473, C2V_268_513, C2V_268_549, C2V_268_611, C2V_268_636, C2V_268_682, C2V_268_899, C2V_268_923, C2V_268_1007, C2V_268_1037, C2V_268_1064, C2V_268_1128, C2V_268_1419, C2V_268_1420, C2V_269_43, C2V_269_53, C2V_269_136, C2V_269_159, C2V_269_223, C2V_269_241, C2V_269_290, C2V_269_357, C2V_269_436, C2V_269_718, C2V_269_734, C2V_269_788, C2V_269_866, C2V_269_914, C2V_269_1005, C2V_269_1009, C2V_269_1058, C2V_269_1106, C2V_269_1420, C2V_269_1421, C2V_270_26, C2V_270_50, C2V_270_138, C2V_270_158, C2V_270_240, C2V_270_271, C2V_270_324, C2V_270_476, C2V_270_573, C2V_270_606, C2V_270_810, C2V_270_838, C2V_270_871, C2V_270_933, C2V_270_968, C2V_270_1035, C2V_270_1099, C2V_270_1149, C2V_270_1421, C2V_270_1422, C2V_271_2, C2V_271_86, C2V_271_106, C2V_271_167, C2V_271_229, C2V_271_272, C2V_271_372, C2V_271_426, C2V_271_523, C2V_271_759, C2V_271_807, C2V_271_855, C2V_271_896, C2V_271_937, C2V_271_971, C2V_271_1010, C2V_271_1084, C2V_271_1143, C2V_271_1422, C2V_271_1423, C2V_272_11, C2V_272_60, C2V_272_116, C2V_272_164, C2V_272_193, C2V_272_262, C2V_272_313, C2V_272_420, C2V_272_509, C2V_272_669, C2V_272_682, C2V_272_850, C2V_272_892, C2V_272_955, C2V_272_986, C2V_272_1018, C2V_272_1085, C2V_272_1116, C2V_272_1423, C2V_272_1424, C2V_273_6, C2V_273_81, C2V_273_98, C2V_273_180, C2V_273_198, C2V_273_265, C2V_273_362, C2V_273_417, C2V_273_576, C2V_273_585, C2V_273_661, C2V_273_765, C2V_273_896, C2V_273_940, C2V_273_965, C2V_273_1025, C2V_273_1103, C2V_273_1148, C2V_273_1424, C2V_273_1425, C2V_274_25, C2V_274_84, C2V_274_123, C2V_274_179, C2V_274_196, C2V_274_250, C2V_274_474, C2V_274_514, C2V_274_550, C2V_274_612, C2V_274_637, C2V_274_683, C2V_274_900, C2V_274_924, C2V_274_1008, C2V_274_1038, C2V_274_1065, C2V_274_1129, C2V_274_1425, C2V_274_1426, C2V_275_44, C2V_275_54, C2V_275_137, C2V_275_160, C2V_275_224, C2V_275_242, C2V_275_291, C2V_275_358, C2V_275_437, C2V_275_719, C2V_275_735, C2V_275_789, C2V_275_867, C2V_275_915, C2V_275_1006, C2V_275_1010, C2V_275_1059, C2V_275_1107, C2V_275_1426, C2V_275_1427, C2V_276_27, C2V_276_51, C2V_276_139, C2V_276_159, C2V_276_193, C2V_276_272, C2V_276_325, C2V_276_477, C2V_276_574, C2V_276_607, C2V_276_811, C2V_276_839, C2V_276_872, C2V_276_934, C2V_276_969, C2V_276_1036, C2V_276_1100, C2V_276_1150, C2V_276_1427, C2V_276_1428, C2V_277_3, C2V_277_87, C2V_277_107, C2V_277_168, C2V_277_230, C2V_277_273, C2V_277_373, C2V_277_427, C2V_277_524, C2V_277_760, C2V_277_808, C2V_277_856, C2V_277_897, C2V_277_938, C2V_277_972, C2V_277_1011, C2V_277_1085, C2V_277_1144, C2V_277_1428, C2V_277_1429, C2V_278_12, C2V_278_61, C2V_278_117, C2V_278_165, C2V_278_194, C2V_278_263, C2V_278_314, C2V_278_421, C2V_278_510, C2V_278_670, C2V_278_683, C2V_278_851, C2V_278_893, C2V_278_956, C2V_278_987, C2V_278_1019, C2V_278_1086, C2V_278_1117, C2V_278_1429, C2V_278_1430, C2V_279_7, C2V_279_82, C2V_279_99, C2V_279_181, C2V_279_199, C2V_279_266, C2V_279_363, C2V_279_418, C2V_279_529, C2V_279_586, C2V_279_662, C2V_279_766, C2V_279_897, C2V_279_941, C2V_279_966, C2V_279_1026, C2V_279_1104, C2V_279_1149, C2V_279_1430, C2V_279_1431, C2V_280_26, C2V_280_85, C2V_280_124, C2V_280_180, C2V_280_197, C2V_280_251, C2V_280_475, C2V_280_515, C2V_280_551, C2V_280_613, C2V_280_638, C2V_280_684, C2V_280_901, C2V_280_925, C2V_280_961, C2V_280_1039, C2V_280_1066, C2V_280_1130, C2V_280_1431, C2V_280_1432, C2V_281_45, C2V_281_55, C2V_281_138, C2V_281_161, C2V_281_225, C2V_281_243, C2V_281_292, C2V_281_359, C2V_281_438, C2V_281_720, C2V_281_736, C2V_281_790, C2V_281_868, C2V_281_916, C2V_281_1007, C2V_281_1011, C2V_281_1060, C2V_281_1108, C2V_281_1432, C2V_281_1433, C2V_282_28, C2V_282_52, C2V_282_140, C2V_282_160, C2V_282_194, C2V_282_273, C2V_282_326, C2V_282_478, C2V_282_575, C2V_282_608, C2V_282_812, C2V_282_840, C2V_282_873, C2V_282_935, C2V_282_970, C2V_282_1037, C2V_282_1101, C2V_282_1151, C2V_282_1433, C2V_282_1434, C2V_283_4, C2V_283_88, C2V_283_108, C2V_283_169, C2V_283_231, C2V_283_274, C2V_283_374, C2V_283_428, C2V_283_525, C2V_283_761, C2V_283_809, C2V_283_857, C2V_283_898, C2V_283_939, C2V_283_973, C2V_283_1012, C2V_283_1086, C2V_283_1145, C2V_283_1434, C2V_283_1435, C2V_284_13, C2V_284_62, C2V_284_118, C2V_284_166, C2V_284_195, C2V_284_264, C2V_284_315, C2V_284_422, C2V_284_511, C2V_284_671, C2V_284_684, C2V_284_852, C2V_284_894, C2V_284_957, C2V_284_988, C2V_284_1020, C2V_284_1087, C2V_284_1118, C2V_284_1435, C2V_284_1436, C2V_285_8, C2V_285_83, C2V_285_100, C2V_285_182, C2V_285_200, C2V_285_267, C2V_285_364, C2V_285_419, C2V_285_530, C2V_285_587, C2V_285_663, C2V_285_767, C2V_285_898, C2V_285_942, C2V_285_967, C2V_285_1027, C2V_285_1057, C2V_285_1150, C2V_285_1436, C2V_285_1437, C2V_286_27, C2V_286_86, C2V_286_125, C2V_286_181, C2V_286_198, C2V_286_252, C2V_286_476, C2V_286_516, C2V_286_552, C2V_286_614, C2V_286_639, C2V_286_685, C2V_286_902, C2V_286_926, C2V_286_962, C2V_286_1040, C2V_286_1067, C2V_286_1131, C2V_286_1437, C2V_286_1438, C2V_287_46, C2V_287_56, C2V_287_139, C2V_287_162, C2V_287_226, C2V_287_244, C2V_287_293, C2V_287_360, C2V_287_439, C2V_287_673, C2V_287_737, C2V_287_791, C2V_287_869, C2V_287_917, C2V_287_1008, C2V_287_1012, C2V_287_1061, C2V_287_1109, C2V_287_1438, C2V_287_1439, C2V_288_29, C2V_288_53, C2V_288_141, C2V_288_161, C2V_288_195, C2V_288_274, C2V_288_327, C2V_288_479, C2V_288_576, C2V_288_609, C2V_288_813, C2V_288_841, C2V_288_874, C2V_288_936, C2V_288_971, C2V_288_1038, C2V_288_1102, C2V_288_1152, C2V_288_1439, C2V_288_1440, C2V_0_0;
wire [quan_width - 1:0] V2C_5_1, V2C_89_1, V2C_109_1, V2C_170_1, V2C_232_1, V2C_275_1, V2C_375_1, V2C_429_1, V2C_526_1, V2C_762_1, V2C_810_1, V2C_858_1, V2C_899_1, V2C_940_1, V2C_974_1, V2C_1013_1, V2C_1087_1, V2C_1146_1, V2C_1153_1, V2C_14_2, V2C_63_2, V2C_119_2, V2C_167_2, V2C_196_2, V2C_265_2, V2C_316_2, V2C_423_2, V2C_512_2, V2C_672_2, V2C_685_2, V2C_853_2, V2C_895_2, V2C_958_2, V2C_989_2, V2C_1021_2, V2C_1088_2, V2C_1119_2, V2C_1153_2, V2C_1154_2, V2C_9_3, V2C_84_3, V2C_101_3, V2C_183_3, V2C_201_3, V2C_268_3, V2C_365_3, V2C_420_3, V2C_531_3, V2C_588_3, V2C_664_3, V2C_768_3, V2C_899_3, V2C_943_3, V2C_968_3, V2C_1028_3, V2C_1058_3, V2C_1151_3, V2C_1154_3, V2C_1155_3, V2C_28_4, V2C_87_4, V2C_126_4, V2C_182_4, V2C_199_4, V2C_253_4, V2C_477_4, V2C_517_4, V2C_553_4, V2C_615_4, V2C_640_4, V2C_686_4, V2C_903_4, V2C_927_4, V2C_963_4, V2C_1041_4, V2C_1068_4, V2C_1132_4, V2C_1155_4, V2C_1156_4, V2C_47_5, V2C_57_5, V2C_140_5, V2C_163_5, V2C_227_5, V2C_245_5, V2C_294_5, V2C_361_5, V2C_440_5, V2C_674_5, V2C_738_5, V2C_792_5, V2C_870_5, V2C_918_5, V2C_961_5, V2C_1013_5, V2C_1062_5, V2C_1110_5, V2C_1156_5, V2C_1157_5, V2C_30_6, V2C_54_6, V2C_142_6, V2C_162_6, V2C_196_6, V2C_275_6, V2C_328_6, V2C_480_6, V2C_529_6, V2C_610_6, V2C_814_6, V2C_842_6, V2C_875_6, V2C_937_6, V2C_972_6, V2C_1039_6, V2C_1103_6, V2C_1105_6, V2C_1157_6, V2C_1158_6, V2C_6_7, V2C_90_7, V2C_110_7, V2C_171_7, V2C_233_7, V2C_276_7, V2C_376_7, V2C_430_7, V2C_527_7, V2C_763_7, V2C_811_7, V2C_859_7, V2C_900_7, V2C_941_7, V2C_975_7, V2C_1014_7, V2C_1088_7, V2C_1147_7, V2C_1158_7, V2C_1159_7, V2C_15_8, V2C_64_8, V2C_120_8, V2C_168_8, V2C_197_8, V2C_266_8, V2C_317_8, V2C_424_8, V2C_513_8, V2C_625_8, V2C_686_8, V2C_854_8, V2C_896_8, V2C_959_8, V2C_990_8, V2C_1022_8, V2C_1089_8, V2C_1120_8, V2C_1159_8, V2C_1160_8, V2C_10_9, V2C_85_9, V2C_102_9, V2C_184_9, V2C_202_9, V2C_269_9, V2C_366_9, V2C_421_9, V2C_532_9, V2C_589_9, V2C_665_9, V2C_721_9, V2C_900_9, V2C_944_9, V2C_969_9, V2C_1029_9, V2C_1059_9, V2C_1152_9, V2C_1160_9, V2C_1161_9, V2C_29_10, V2C_88_10, V2C_127_10, V2C_183_10, V2C_200_10, V2C_254_10, V2C_478_10, V2C_518_10, V2C_554_10, V2C_616_10, V2C_641_10, V2C_687_10, V2C_904_10, V2C_928_10, V2C_964_10, V2C_1042_10, V2C_1069_10, V2C_1133_10, V2C_1161_10, V2C_1162_10, V2C_48_11, V2C_58_11, V2C_141_11, V2C_164_11, V2C_228_11, V2C_246_11, V2C_295_11, V2C_362_11, V2C_441_11, V2C_675_11, V2C_739_11, V2C_793_11, V2C_871_11, V2C_919_11, V2C_962_11, V2C_1014_11, V2C_1063_11, V2C_1111_11, V2C_1162_11, V2C_1163_11, V2C_31_12, V2C_55_12, V2C_143_12, V2C_163_12, V2C_197_12, V2C_276_12, V2C_329_12, V2C_433_12, V2C_530_12, V2C_611_12, V2C_815_12, V2C_843_12, V2C_876_12, V2C_938_12, V2C_973_12, V2C_1040_12, V2C_1104_12, V2C_1106_12, V2C_1163_12, V2C_1164_12, V2C_7_13, V2C_91_13, V2C_111_13, V2C_172_13, V2C_234_13, V2C_277_13, V2C_377_13, V2C_431_13, V2C_528_13, V2C_764_13, V2C_812_13, V2C_860_13, V2C_901_13, V2C_942_13, V2C_976_13, V2C_1015_13, V2C_1089_13, V2C_1148_13, V2C_1164_13, V2C_1165_13, V2C_16_14, V2C_65_14, V2C_121_14, V2C_169_14, V2C_198_14, V2C_267_14, V2C_318_14, V2C_425_14, V2C_514_14, V2C_626_14, V2C_687_14, V2C_855_14, V2C_897_14, V2C_960_14, V2C_991_14, V2C_1023_14, V2C_1090_14, V2C_1121_14, V2C_1165_14, V2C_1166_14, V2C_11_15, V2C_86_15, V2C_103_15, V2C_185_15, V2C_203_15, V2C_270_15, V2C_367_15, V2C_422_15, V2C_533_15, V2C_590_15, V2C_666_15, V2C_722_15, V2C_901_15, V2C_945_15, V2C_970_15, V2C_1030_15, V2C_1060_15, V2C_1105_15, V2C_1166_15, V2C_1167_15, V2C_30_16, V2C_89_16, V2C_128_16, V2C_184_16, V2C_201_16, V2C_255_16, V2C_479_16, V2C_519_16, V2C_555_16, V2C_617_16, V2C_642_16, V2C_688_16, V2C_905_16, V2C_929_16, V2C_965_16, V2C_1043_16, V2C_1070_16, V2C_1134_16, V2C_1167_16, V2C_1168_16, V2C_1_17, V2C_59_17, V2C_142_17, V2C_165_17, V2C_229_17, V2C_247_17, V2C_296_17, V2C_363_17, V2C_442_17, V2C_676_17, V2C_740_17, V2C_794_17, V2C_872_17, V2C_920_17, V2C_963_17, V2C_1015_17, V2C_1064_17, V2C_1112_17, V2C_1168_17, V2C_1169_17, V2C_32_18, V2C_56_18, V2C_144_18, V2C_164_18, V2C_198_18, V2C_277_18, V2C_330_18, V2C_434_18, V2C_531_18, V2C_612_18, V2C_816_18, V2C_844_18, V2C_877_18, V2C_939_18, V2C_974_18, V2C_1041_18, V2C_1057_18, V2C_1107_18, V2C_1169_18, V2C_1170_18, V2C_8_19, V2C_92_19, V2C_112_19, V2C_173_19, V2C_235_19, V2C_278_19, V2C_378_19, V2C_432_19, V2C_481_19, V2C_765_19, V2C_813_19, V2C_861_19, V2C_902_19, V2C_943_19, V2C_977_19, V2C_1016_19, V2C_1090_19, V2C_1149_19, V2C_1170_19, V2C_1171_19, V2C_17_20, V2C_66_20, V2C_122_20, V2C_170_20, V2C_199_20, V2C_268_20, V2C_319_20, V2C_426_20, V2C_515_20, V2C_627_20, V2C_688_20, V2C_856_20, V2C_898_20, V2C_913_20, V2C_992_20, V2C_1024_20, V2C_1091_20, V2C_1122_20, V2C_1171_20, V2C_1172_20, V2C_12_21, V2C_87_21, V2C_104_21, V2C_186_21, V2C_204_21, V2C_271_21, V2C_368_21, V2C_423_21, V2C_534_21, V2C_591_21, V2C_667_21, V2C_723_21, V2C_902_21, V2C_946_21, V2C_971_21, V2C_1031_21, V2C_1061_21, V2C_1106_21, V2C_1172_21, V2C_1173_21, V2C_31_22, V2C_90_22, V2C_129_22, V2C_185_22, V2C_202_22, V2C_256_22, V2C_480_22, V2C_520_22, V2C_556_22, V2C_618_22, V2C_643_22, V2C_689_22, V2C_906_22, V2C_930_22, V2C_966_22, V2C_1044_22, V2C_1071_22, V2C_1135_22, V2C_1173_22, V2C_1174_22, V2C_2_23, V2C_60_23, V2C_143_23, V2C_166_23, V2C_230_23, V2C_248_23, V2C_297_23, V2C_364_23, V2C_443_23, V2C_677_23, V2C_741_23, V2C_795_23, V2C_873_23, V2C_921_23, V2C_964_23, V2C_1016_23, V2C_1065_23, V2C_1113_23, V2C_1174_23, V2C_1175_23, V2C_33_24, V2C_57_24, V2C_97_24, V2C_165_24, V2C_199_24, V2C_278_24, V2C_331_24, V2C_435_24, V2C_532_24, V2C_613_24, V2C_769_24, V2C_845_24, V2C_878_24, V2C_940_24, V2C_975_24, V2C_1042_24, V2C_1058_24, V2C_1108_24, V2C_1175_24, V2C_1176_24, V2C_9_25, V2C_93_25, V2C_113_25, V2C_174_25, V2C_236_25, V2C_279_25, V2C_379_25, V2C_385_25, V2C_482_25, V2C_766_25, V2C_814_25, V2C_862_25, V2C_903_25, V2C_944_25, V2C_978_25, V2C_1017_25, V2C_1091_25, V2C_1150_25, V2C_1176_25, V2C_1177_25, V2C_18_26, V2C_67_26, V2C_123_26, V2C_171_26, V2C_200_26, V2C_269_26, V2C_320_26, V2C_427_26, V2C_516_26, V2C_628_26, V2C_689_26, V2C_857_26, V2C_899_26, V2C_914_26, V2C_993_26, V2C_1025_26, V2C_1092_26, V2C_1123_26, V2C_1177_26, V2C_1178_26, V2C_13_27, V2C_88_27, V2C_105_27, V2C_187_27, V2C_205_27, V2C_272_27, V2C_369_27, V2C_424_27, V2C_535_27, V2C_592_27, V2C_668_27, V2C_724_27, V2C_903_27, V2C_947_27, V2C_972_27, V2C_1032_27, V2C_1062_27, V2C_1107_27, V2C_1178_27, V2C_1179_27, V2C_32_28, V2C_91_28, V2C_130_28, V2C_186_28, V2C_203_28, V2C_257_28, V2C_433_28, V2C_521_28, V2C_557_28, V2C_619_28, V2C_644_28, V2C_690_28, V2C_907_28, V2C_931_28, V2C_967_28, V2C_1045_28, V2C_1072_28, V2C_1136_28, V2C_1179_28, V2C_1180_28, V2C_3_29, V2C_61_29, V2C_144_29, V2C_167_29, V2C_231_29, V2C_249_29, V2C_298_29, V2C_365_29, V2C_444_29, V2C_678_29, V2C_742_29, V2C_796_29, V2C_874_29, V2C_922_29, V2C_965_29, V2C_1017_29, V2C_1066_29, V2C_1114_29, V2C_1180_29, V2C_1181_29, V2C_34_30, V2C_58_30, V2C_98_30, V2C_166_30, V2C_200_30, V2C_279_30, V2C_332_30, V2C_436_30, V2C_533_30, V2C_614_30, V2C_770_30, V2C_846_30, V2C_879_30, V2C_941_30, V2C_976_30, V2C_1043_30, V2C_1059_30, V2C_1109_30, V2C_1181_30, V2C_1182_30, V2C_10_31, V2C_94_31, V2C_114_31, V2C_175_31, V2C_237_31, V2C_280_31, V2C_380_31, V2C_386_31, V2C_483_31, V2C_767_31, V2C_815_31, V2C_863_31, V2C_904_31, V2C_945_31, V2C_979_31, V2C_1018_31, V2C_1092_31, V2C_1151_31, V2C_1182_31, V2C_1183_31, V2C_19_32, V2C_68_32, V2C_124_32, V2C_172_32, V2C_201_32, V2C_270_32, V2C_321_32, V2C_428_32, V2C_517_32, V2C_629_32, V2C_690_32, V2C_858_32, V2C_900_32, V2C_915_32, V2C_994_32, V2C_1026_32, V2C_1093_32, V2C_1124_32, V2C_1183_32, V2C_1184_32, V2C_14_33, V2C_89_33, V2C_106_33, V2C_188_33, V2C_206_33, V2C_273_33, V2C_370_33, V2C_425_33, V2C_536_33, V2C_593_33, V2C_669_33, V2C_725_33, V2C_904_33, V2C_948_33, V2C_973_33, V2C_1033_33, V2C_1063_33, V2C_1108_33, V2C_1184_33, V2C_1185_33, V2C_33_34, V2C_92_34, V2C_131_34, V2C_187_34, V2C_204_34, V2C_258_34, V2C_434_34, V2C_522_34, V2C_558_34, V2C_620_34, V2C_645_34, V2C_691_34, V2C_908_34, V2C_932_34, V2C_968_34, V2C_1046_34, V2C_1073_34, V2C_1137_34, V2C_1185_34, V2C_1186_34, V2C_4_35, V2C_62_35, V2C_97_35, V2C_168_35, V2C_232_35, V2C_250_35, V2C_299_35, V2C_366_35, V2C_445_35, V2C_679_35, V2C_743_35, V2C_797_35, V2C_875_35, V2C_923_35, V2C_966_35, V2C_1018_35, V2C_1067_35, V2C_1115_35, V2C_1186_35, V2C_1187_35, V2C_35_36, V2C_59_36, V2C_99_36, V2C_167_36, V2C_201_36, V2C_280_36, V2C_333_36, V2C_437_36, V2C_534_36, V2C_615_36, V2C_771_36, V2C_847_36, V2C_880_36, V2C_942_36, V2C_977_36, V2C_1044_36, V2C_1060_36, V2C_1110_36, V2C_1187_36, V2C_1188_36, V2C_11_37, V2C_95_37, V2C_115_37, V2C_176_37, V2C_238_37, V2C_281_37, V2C_381_37, V2C_387_37, V2C_484_37, V2C_768_37, V2C_816_37, V2C_864_37, V2C_905_37, V2C_946_37, V2C_980_37, V2C_1019_37, V2C_1093_37, V2C_1152_37, V2C_1188_37, V2C_1189_37, V2C_20_38, V2C_69_38, V2C_125_38, V2C_173_38, V2C_202_38, V2C_271_38, V2C_322_38, V2C_429_38, V2C_518_38, V2C_630_38, V2C_691_38, V2C_859_38, V2C_901_38, V2C_916_38, V2C_995_38, V2C_1027_38, V2C_1094_38, V2C_1125_38, V2C_1189_38, V2C_1190_38, V2C_15_39, V2C_90_39, V2C_107_39, V2C_189_39, V2C_207_39, V2C_274_39, V2C_371_39, V2C_426_39, V2C_537_39, V2C_594_39, V2C_670_39, V2C_726_39, V2C_905_39, V2C_949_39, V2C_974_39, V2C_1034_39, V2C_1064_39, V2C_1109_39, V2C_1190_39, V2C_1191_39, V2C_34_40, V2C_93_40, V2C_132_40, V2C_188_40, V2C_205_40, V2C_259_40, V2C_435_40, V2C_523_40, V2C_559_40, V2C_621_40, V2C_646_40, V2C_692_40, V2C_909_40, V2C_933_40, V2C_969_40, V2C_1047_40, V2C_1074_40, V2C_1138_40, V2C_1191_40, V2C_1192_40, V2C_5_41, V2C_63_41, V2C_98_41, V2C_169_41, V2C_233_41, V2C_251_41, V2C_300_41, V2C_367_41, V2C_446_41, V2C_680_41, V2C_744_41, V2C_798_41, V2C_876_41, V2C_924_41, V2C_967_41, V2C_1019_41, V2C_1068_41, V2C_1116_41, V2C_1192_41, V2C_1193_41, V2C_36_42, V2C_60_42, V2C_100_42, V2C_168_42, V2C_202_42, V2C_281_42, V2C_334_42, V2C_438_42, V2C_535_42, V2C_616_42, V2C_772_42, V2C_848_42, V2C_881_42, V2C_943_42, V2C_978_42, V2C_1045_42, V2C_1061_42, V2C_1111_42, V2C_1193_42, V2C_1194_42, V2C_12_43, V2C_96_43, V2C_116_43, V2C_177_43, V2C_239_43, V2C_282_43, V2C_382_43, V2C_388_43, V2C_485_43, V2C_721_43, V2C_769_43, V2C_817_43, V2C_906_43, V2C_947_43, V2C_981_43, V2C_1020_43, V2C_1094_43, V2C_1105_43, V2C_1194_43, V2C_1195_43, V2C_21_44, V2C_70_44, V2C_126_44, V2C_174_44, V2C_203_44, V2C_272_44, V2C_323_44, V2C_430_44, V2C_519_44, V2C_631_44, V2C_692_44, V2C_860_44, V2C_902_44, V2C_917_44, V2C_996_44, V2C_1028_44, V2C_1095_44, V2C_1126_44, V2C_1195_44, V2C_1196_44, V2C_16_45, V2C_91_45, V2C_108_45, V2C_190_45, V2C_208_45, V2C_275_45, V2C_372_45, V2C_427_45, V2C_538_45, V2C_595_45, V2C_671_45, V2C_727_45, V2C_906_45, V2C_950_45, V2C_975_45, V2C_1035_45, V2C_1065_45, V2C_1110_45, V2C_1196_45, V2C_1197_45, V2C_35_46, V2C_94_46, V2C_133_46, V2C_189_46, V2C_206_46, V2C_260_46, V2C_436_46, V2C_524_46, V2C_560_46, V2C_622_46, V2C_647_46, V2C_693_46, V2C_910_46, V2C_934_46, V2C_970_46, V2C_1048_46, V2C_1075_46, V2C_1139_46, V2C_1197_46, V2C_1198_46, V2C_6_47, V2C_64_47, V2C_99_47, V2C_170_47, V2C_234_47, V2C_252_47, V2C_301_47, V2C_368_47, V2C_447_47, V2C_681_47, V2C_745_47, V2C_799_47, V2C_877_47, V2C_925_47, V2C_968_47, V2C_1020_47, V2C_1069_47, V2C_1117_47, V2C_1198_47, V2C_1199_47, V2C_37_48, V2C_61_48, V2C_101_48, V2C_169_48, V2C_203_48, V2C_282_48, V2C_335_48, V2C_439_48, V2C_536_48, V2C_617_48, V2C_773_48, V2C_849_48, V2C_882_48, V2C_944_48, V2C_979_48, V2C_1046_48, V2C_1062_48, V2C_1112_48, V2C_1199_48, V2C_1200_48, V2C_13_49, V2C_49_49, V2C_117_49, V2C_178_49, V2C_240_49, V2C_283_49, V2C_383_49, V2C_389_49, V2C_486_49, V2C_722_49, V2C_770_49, V2C_818_49, V2C_907_49, V2C_948_49, V2C_982_49, V2C_1021_49, V2C_1095_49, V2C_1106_49, V2C_1200_49, V2C_1201_49, V2C_22_50, V2C_71_50, V2C_127_50, V2C_175_50, V2C_204_50, V2C_273_50, V2C_324_50, V2C_431_50, V2C_520_50, V2C_632_50, V2C_693_50, V2C_861_50, V2C_903_50, V2C_918_50, V2C_997_50, V2C_1029_50, V2C_1096_50, V2C_1127_50, V2C_1201_50, V2C_1202_50, V2C_17_51, V2C_92_51, V2C_109_51, V2C_191_51, V2C_209_51, V2C_276_51, V2C_373_51, V2C_428_51, V2C_539_51, V2C_596_51, V2C_672_51, V2C_728_51, V2C_907_51, V2C_951_51, V2C_976_51, V2C_1036_51, V2C_1066_51, V2C_1111_51, V2C_1202_51, V2C_1203_51, V2C_36_52, V2C_95_52, V2C_134_52, V2C_190_52, V2C_207_52, V2C_261_52, V2C_437_52, V2C_525_52, V2C_561_52, V2C_623_52, V2C_648_52, V2C_694_52, V2C_911_52, V2C_935_52, V2C_971_52, V2C_1049_52, V2C_1076_52, V2C_1140_52, V2C_1203_52, V2C_1204_52, V2C_7_53, V2C_65_53, V2C_100_53, V2C_171_53, V2C_235_53, V2C_253_53, V2C_302_53, V2C_369_53, V2C_448_53, V2C_682_53, V2C_746_53, V2C_800_53, V2C_878_53, V2C_926_53, V2C_969_53, V2C_1021_53, V2C_1070_53, V2C_1118_53, V2C_1204_53, V2C_1205_53, V2C_38_54, V2C_62_54, V2C_102_54, V2C_170_54, V2C_204_54, V2C_283_54, V2C_336_54, V2C_440_54, V2C_537_54, V2C_618_54, V2C_774_54, V2C_850_54, V2C_883_54, V2C_945_54, V2C_980_54, V2C_1047_54, V2C_1063_54, V2C_1113_54, V2C_1205_54, V2C_1206_54, V2C_14_55, V2C_50_55, V2C_118_55, V2C_179_55, V2C_193_55, V2C_284_55, V2C_384_55, V2C_390_55, V2C_487_55, V2C_723_55, V2C_771_55, V2C_819_55, V2C_908_55, V2C_949_55, V2C_983_55, V2C_1022_55, V2C_1096_55, V2C_1107_55, V2C_1206_55, V2C_1207_55, V2C_23_56, V2C_72_56, V2C_128_56, V2C_176_56, V2C_205_56, V2C_274_56, V2C_325_56, V2C_432_56, V2C_521_56, V2C_633_56, V2C_694_56, V2C_862_56, V2C_904_56, V2C_919_56, V2C_998_56, V2C_1030_56, V2C_1097_56, V2C_1128_56, V2C_1207_56, V2C_1208_56, V2C_18_57, V2C_93_57, V2C_110_57, V2C_192_57, V2C_210_57, V2C_277_57, V2C_374_57, V2C_429_57, V2C_540_57, V2C_597_57, V2C_625_57, V2C_729_57, V2C_908_57, V2C_952_57, V2C_977_57, V2C_1037_57, V2C_1067_57, V2C_1112_57, V2C_1208_57, V2C_1209_57, V2C_37_58, V2C_96_58, V2C_135_58, V2C_191_58, V2C_208_58, V2C_262_58, V2C_438_58, V2C_526_58, V2C_562_58, V2C_624_58, V2C_649_58, V2C_695_58, V2C_912_58, V2C_936_58, V2C_972_58, V2C_1050_58, V2C_1077_58, V2C_1141_58, V2C_1209_58, V2C_1210_58, V2C_8_59, V2C_66_59, V2C_101_59, V2C_172_59, V2C_236_59, V2C_254_59, V2C_303_59, V2C_370_59, V2C_449_59, V2C_683_59, V2C_747_59, V2C_801_59, V2C_879_59, V2C_927_59, V2C_970_59, V2C_1022_59, V2C_1071_59, V2C_1119_59, V2C_1210_59, V2C_1211_59, V2C_39_60, V2C_63_60, V2C_103_60, V2C_171_60, V2C_205_60, V2C_284_60, V2C_289_60, V2C_441_60, V2C_538_60, V2C_619_60, V2C_775_60, V2C_851_60, V2C_884_60, V2C_946_60, V2C_981_60, V2C_1048_60, V2C_1064_60, V2C_1114_60, V2C_1211_60, V2C_1212_60, V2C_15_61, V2C_51_61, V2C_119_61, V2C_180_61, V2C_194_61, V2C_285_61, V2C_337_61, V2C_391_61, V2C_488_61, V2C_724_61, V2C_772_61, V2C_820_61, V2C_909_61, V2C_950_61, V2C_984_61, V2C_1023_61, V2C_1097_61, V2C_1108_61, V2C_1212_61, V2C_1213_61, V2C_24_62, V2C_73_62, V2C_129_62, V2C_177_62, V2C_206_62, V2C_275_62, V2C_326_62, V2C_385_62, V2C_522_62, V2C_634_62, V2C_695_62, V2C_863_62, V2C_905_62, V2C_920_62, V2C_999_62, V2C_1031_62, V2C_1098_62, V2C_1129_62, V2C_1213_62, V2C_1214_62, V2C_19_63, V2C_94_63, V2C_111_63, V2C_145_63, V2C_211_63, V2C_278_63, V2C_375_63, V2C_430_63, V2C_541_63, V2C_598_63, V2C_626_63, V2C_730_63, V2C_909_63, V2C_953_63, V2C_978_63, V2C_1038_63, V2C_1068_63, V2C_1113_63, V2C_1214_63, V2C_1215_63, V2C_38_64, V2C_49_64, V2C_136_64, V2C_192_64, V2C_209_64, V2C_263_64, V2C_439_64, V2C_527_64, V2C_563_64, V2C_577_64, V2C_650_64, V2C_696_64, V2C_865_64, V2C_937_64, V2C_973_64, V2C_1051_64, V2C_1078_64, V2C_1142_64, V2C_1215_64, V2C_1216_64, V2C_9_65, V2C_67_65, V2C_102_65, V2C_173_65, V2C_237_65, V2C_255_65, V2C_304_65, V2C_371_65, V2C_450_65, V2C_684_65, V2C_748_65, V2C_802_65, V2C_880_65, V2C_928_65, V2C_971_65, V2C_1023_65, V2C_1072_65, V2C_1120_65, V2C_1216_65, V2C_1217_65, V2C_40_66, V2C_64_66, V2C_104_66, V2C_172_66, V2C_206_66, V2C_285_66, V2C_290_66, V2C_442_66, V2C_539_66, V2C_620_66, V2C_776_66, V2C_852_66, V2C_885_66, V2C_947_66, V2C_982_66, V2C_1049_66, V2C_1065_66, V2C_1115_66, V2C_1217_66, V2C_1218_66, V2C_16_67, V2C_52_67, V2C_120_67, V2C_181_67, V2C_195_67, V2C_286_67, V2C_338_67, V2C_392_67, V2C_489_67, V2C_725_67, V2C_773_67, V2C_821_67, V2C_910_67, V2C_951_67, V2C_985_67, V2C_1024_67, V2C_1098_67, V2C_1109_67, V2C_1218_67, V2C_1219_67, V2C_25_68, V2C_74_68, V2C_130_68, V2C_178_68, V2C_207_68, V2C_276_68, V2C_327_68, V2C_386_68, V2C_523_68, V2C_635_68, V2C_696_68, V2C_864_68, V2C_906_68, V2C_921_68, V2C_1000_68, V2C_1032_68, V2C_1099_68, V2C_1130_68, V2C_1219_68, V2C_1220_68, V2C_20_69, V2C_95_69, V2C_112_69, V2C_146_69, V2C_212_69, V2C_279_69, V2C_376_69, V2C_431_69, V2C_542_69, V2C_599_69, V2C_627_69, V2C_731_69, V2C_910_69, V2C_954_69, V2C_979_69, V2C_1039_69, V2C_1069_69, V2C_1114_69, V2C_1220_69, V2C_1221_69, V2C_39_70, V2C_50_70, V2C_137_70, V2C_145_70, V2C_210_70, V2C_264_70, V2C_440_70, V2C_528_70, V2C_564_70, V2C_578_70, V2C_651_70, V2C_697_70, V2C_866_70, V2C_938_70, V2C_974_70, V2C_1052_70, V2C_1079_70, V2C_1143_70, V2C_1221_70, V2C_1222_70, V2C_10_71, V2C_68_71, V2C_103_71, V2C_174_71, V2C_238_71, V2C_256_71, V2C_305_71, V2C_372_71, V2C_451_71, V2C_685_71, V2C_749_71, V2C_803_71, V2C_881_71, V2C_929_71, V2C_972_71, V2C_1024_71, V2C_1073_71, V2C_1121_71, V2C_1222_71, V2C_1223_71, V2C_41_72, V2C_65_72, V2C_105_72, V2C_173_72, V2C_207_72, V2C_286_72, V2C_291_72, V2C_443_72, V2C_540_72, V2C_621_72, V2C_777_72, V2C_853_72, V2C_886_72, V2C_948_72, V2C_983_72, V2C_1050_72, V2C_1066_72, V2C_1116_72, V2C_1223_72, V2C_1224_72, V2C_17_73, V2C_53_73, V2C_121_73, V2C_182_73, V2C_196_73, V2C_287_73, V2C_339_73, V2C_393_73, V2C_490_73, V2C_726_73, V2C_774_73, V2C_822_73, V2C_911_73, V2C_952_73, V2C_986_73, V2C_1025_73, V2C_1099_73, V2C_1110_73, V2C_1224_73, V2C_1225_73, V2C_26_74, V2C_75_74, V2C_131_74, V2C_179_74, V2C_208_74, V2C_277_74, V2C_328_74, V2C_387_74, V2C_524_74, V2C_636_74, V2C_697_74, V2C_817_74, V2C_907_74, V2C_922_74, V2C_1001_74, V2C_1033_74, V2C_1100_74, V2C_1131_74, V2C_1225_74, V2C_1226_74, V2C_21_75, V2C_96_75, V2C_113_75, V2C_147_75, V2C_213_75, V2C_280_75, V2C_377_75, V2C_432_75, V2C_543_75, V2C_600_75, V2C_628_75, V2C_732_75, V2C_911_75, V2C_955_75, V2C_980_75, V2C_1040_75, V2C_1070_75, V2C_1115_75, V2C_1226_75, V2C_1227_75, V2C_40_76, V2C_51_76, V2C_138_76, V2C_146_76, V2C_211_76, V2C_265_76, V2C_441_76, V2C_481_76, V2C_565_76, V2C_579_76, V2C_652_76, V2C_698_76, V2C_867_76, V2C_939_76, V2C_975_76, V2C_1053_76, V2C_1080_76, V2C_1144_76, V2C_1227_76, V2C_1228_76, V2C_11_77, V2C_69_77, V2C_104_77, V2C_175_77, V2C_239_77, V2C_257_77, V2C_306_77, V2C_373_77, V2C_452_77, V2C_686_77, V2C_750_77, V2C_804_77, V2C_882_77, V2C_930_77, V2C_973_77, V2C_1025_77, V2C_1074_77, V2C_1122_77, V2C_1228_77, V2C_1229_77, V2C_42_78, V2C_66_78, V2C_106_78, V2C_174_78, V2C_208_78, V2C_287_78, V2C_292_78, V2C_444_78, V2C_541_78, V2C_622_78, V2C_778_78, V2C_854_78, V2C_887_78, V2C_949_78, V2C_984_78, V2C_1051_78, V2C_1067_78, V2C_1117_78, V2C_1229_78, V2C_1230_78, V2C_18_79, V2C_54_79, V2C_122_79, V2C_183_79, V2C_197_79, V2C_288_79, V2C_340_79, V2C_394_79, V2C_491_79, V2C_727_79, V2C_775_79, V2C_823_79, V2C_912_79, V2C_953_79, V2C_987_79, V2C_1026_79, V2C_1100_79, V2C_1111_79, V2C_1230_79, V2C_1231_79, V2C_27_80, V2C_76_80, V2C_132_80, V2C_180_80, V2C_209_80, V2C_278_80, V2C_329_80, V2C_388_80, V2C_525_80, V2C_637_80, V2C_698_80, V2C_818_80, V2C_908_80, V2C_923_80, V2C_1002_80, V2C_1034_80, V2C_1101_80, V2C_1132_80, V2C_1231_80, V2C_1232_80, V2C_22_81, V2C_49_81, V2C_114_81, V2C_148_81, V2C_214_81, V2C_281_81, V2C_378_81, V2C_385_81, V2C_544_81, V2C_601_81, V2C_629_81, V2C_733_81, V2C_912_81, V2C_956_81, V2C_981_81, V2C_1041_81, V2C_1071_81, V2C_1116_81, V2C_1232_81, V2C_1233_81, V2C_41_82, V2C_52_82, V2C_139_82, V2C_147_82, V2C_212_82, V2C_266_82, V2C_442_82, V2C_482_82, V2C_566_82, V2C_580_82, V2C_653_82, V2C_699_82, V2C_868_82, V2C_940_82, V2C_976_82, V2C_1054_82, V2C_1081_82, V2C_1145_82, V2C_1233_82, V2C_1234_82, V2C_12_83, V2C_70_83, V2C_105_83, V2C_176_83, V2C_240_83, V2C_258_83, V2C_307_83, V2C_374_83, V2C_453_83, V2C_687_83, V2C_751_83, V2C_805_83, V2C_883_83, V2C_931_83, V2C_974_83, V2C_1026_83, V2C_1075_83, V2C_1123_83, V2C_1234_83, V2C_1235_83, V2C_43_84, V2C_67_84, V2C_107_84, V2C_175_84, V2C_209_84, V2C_288_84, V2C_293_84, V2C_445_84, V2C_542_84, V2C_623_84, V2C_779_84, V2C_855_84, V2C_888_84, V2C_950_84, V2C_985_84, V2C_1052_84, V2C_1068_84, V2C_1118_84, V2C_1235_84, V2C_1236_84, V2C_19_85, V2C_55_85, V2C_123_85, V2C_184_85, V2C_198_85, V2C_241_85, V2C_341_85, V2C_395_85, V2C_492_85, V2C_728_85, V2C_776_85, V2C_824_85, V2C_865_85, V2C_954_85, V2C_988_85, V2C_1027_85, V2C_1101_85, V2C_1112_85, V2C_1236_85, V2C_1237_85, V2C_28_86, V2C_77_86, V2C_133_86, V2C_181_86, V2C_210_86, V2C_279_86, V2C_330_86, V2C_389_86, V2C_526_86, V2C_638_86, V2C_699_86, V2C_819_86, V2C_909_86, V2C_924_86, V2C_1003_86, V2C_1035_86, V2C_1102_86, V2C_1133_86, V2C_1237_86, V2C_1238_86, V2C_23_87, V2C_50_87, V2C_115_87, V2C_149_87, V2C_215_87, V2C_282_87, V2C_379_87, V2C_386_87, V2C_545_87, V2C_602_87, V2C_630_87, V2C_734_87, V2C_865_87, V2C_957_87, V2C_982_87, V2C_1042_87, V2C_1072_87, V2C_1117_87, V2C_1238_87, V2C_1239_87, V2C_42_88, V2C_53_88, V2C_140_88, V2C_148_88, V2C_213_88, V2C_267_88, V2C_443_88, V2C_483_88, V2C_567_88, V2C_581_88, V2C_654_88, V2C_700_88, V2C_869_88, V2C_941_88, V2C_977_88, V2C_1055_88, V2C_1082_88, V2C_1146_88, V2C_1239_88, V2C_1240_88, V2C_13_89, V2C_71_89, V2C_106_89, V2C_177_89, V2C_193_89, V2C_259_89, V2C_308_89, V2C_375_89, V2C_454_89, V2C_688_89, V2C_752_89, V2C_806_89, V2C_884_89, V2C_932_89, V2C_975_89, V2C_1027_89, V2C_1076_89, V2C_1124_89, V2C_1240_89, V2C_1241_89, V2C_44_90, V2C_68_90, V2C_108_90, V2C_176_90, V2C_210_90, V2C_241_90, V2C_294_90, V2C_446_90, V2C_543_90, V2C_624_90, V2C_780_90, V2C_856_90, V2C_889_90, V2C_951_90, V2C_986_90, V2C_1053_90, V2C_1069_90, V2C_1119_90, V2C_1241_90, V2C_1242_90, V2C_20_91, V2C_56_91, V2C_124_91, V2C_185_91, V2C_199_91, V2C_242_91, V2C_342_91, V2C_396_91, V2C_493_91, V2C_729_91, V2C_777_91, V2C_825_91, V2C_866_91, V2C_955_91, V2C_989_91, V2C_1028_91, V2C_1102_91, V2C_1113_91, V2C_1242_91, V2C_1243_91, V2C_29_92, V2C_78_92, V2C_134_92, V2C_182_92, V2C_211_92, V2C_280_92, V2C_331_92, V2C_390_92, V2C_527_92, V2C_639_92, V2C_700_92, V2C_820_92, V2C_910_92, V2C_925_92, V2C_1004_92, V2C_1036_92, V2C_1103_92, V2C_1134_92, V2C_1243_92, V2C_1244_92, V2C_24_93, V2C_51_93, V2C_116_93, V2C_150_93, V2C_216_93, V2C_283_93, V2C_380_93, V2C_387_93, V2C_546_93, V2C_603_93, V2C_631_93, V2C_735_93, V2C_866_93, V2C_958_93, V2C_983_93, V2C_1043_93, V2C_1073_93, V2C_1118_93, V2C_1244_93, V2C_1245_93, V2C_43_94, V2C_54_94, V2C_141_94, V2C_149_94, V2C_214_94, V2C_268_94, V2C_444_94, V2C_484_94, V2C_568_94, V2C_582_94, V2C_655_94, V2C_701_94, V2C_870_94, V2C_942_94, V2C_978_94, V2C_1056_94, V2C_1083_94, V2C_1147_94, V2C_1245_94, V2C_1246_94, V2C_14_95, V2C_72_95, V2C_107_95, V2C_178_95, V2C_194_95, V2C_260_95, V2C_309_95, V2C_376_95, V2C_455_95, V2C_689_95, V2C_753_95, V2C_807_95, V2C_885_95, V2C_933_95, V2C_976_95, V2C_1028_95, V2C_1077_95, V2C_1125_95, V2C_1246_95, V2C_1247_95, V2C_45_96, V2C_69_96, V2C_109_96, V2C_177_96, V2C_211_96, V2C_242_96, V2C_295_96, V2C_447_96, V2C_544_96, V2C_577_96, V2C_781_96, V2C_857_96, V2C_890_96, V2C_952_96, V2C_987_96, V2C_1054_96, V2C_1070_96, V2C_1120_96, V2C_1247_96, V2C_1248_96, V2C_21_97, V2C_57_97, V2C_125_97, V2C_186_97, V2C_200_97, V2C_243_97, V2C_343_97, V2C_397_97, V2C_494_97, V2C_730_97, V2C_778_97, V2C_826_97, V2C_867_97, V2C_956_97, V2C_990_97, V2C_1029_97, V2C_1103_97, V2C_1114_97, V2C_1248_97, V2C_1249_97, V2C_30_98, V2C_79_98, V2C_135_98, V2C_183_98, V2C_212_98, V2C_281_98, V2C_332_98, V2C_391_98, V2C_528_98, V2C_640_98, V2C_701_98, V2C_821_98, V2C_911_98, V2C_926_98, V2C_1005_98, V2C_1037_98, V2C_1104_98, V2C_1135_98, V2C_1249_98, V2C_1250_98, V2C_25_99, V2C_52_99, V2C_117_99, V2C_151_99, V2C_217_99, V2C_284_99, V2C_381_99, V2C_388_99, V2C_547_99, V2C_604_99, V2C_632_99, V2C_736_99, V2C_867_99, V2C_959_99, V2C_984_99, V2C_1044_99, V2C_1074_99, V2C_1119_99, V2C_1250_99, V2C_1251_99, V2C_44_100, V2C_55_100, V2C_142_100, V2C_150_100, V2C_215_100, V2C_269_100, V2C_445_100, V2C_485_100, V2C_569_100, V2C_583_100, V2C_656_100, V2C_702_100, V2C_871_100, V2C_943_100, V2C_979_100, V2C_1009_100, V2C_1084_100, V2C_1148_100, V2C_1251_100, V2C_1252_100, V2C_15_101, V2C_73_101, V2C_108_101, V2C_179_101, V2C_195_101, V2C_261_101, V2C_310_101, V2C_377_101, V2C_456_101, V2C_690_101, V2C_754_101, V2C_808_101, V2C_886_101, V2C_934_101, V2C_977_101, V2C_1029_101, V2C_1078_101, V2C_1126_101, V2C_1252_101, V2C_1253_101, V2C_46_102, V2C_70_102, V2C_110_102, V2C_178_102, V2C_212_102, V2C_243_102, V2C_296_102, V2C_448_102, V2C_545_102, V2C_578_102, V2C_782_102, V2C_858_102, V2C_891_102, V2C_953_102, V2C_988_102, V2C_1055_102, V2C_1071_102, V2C_1121_102, V2C_1253_102, V2C_1254_102, V2C_22_103, V2C_58_103, V2C_126_103, V2C_187_103, V2C_201_103, V2C_244_103, V2C_344_103, V2C_398_103, V2C_495_103, V2C_731_103, V2C_779_103, V2C_827_103, V2C_868_103, V2C_957_103, V2C_991_103, V2C_1030_103, V2C_1104_103, V2C_1115_103, V2C_1254_103, V2C_1255_103, V2C_31_104, V2C_80_104, V2C_136_104, V2C_184_104, V2C_213_104, V2C_282_104, V2C_333_104, V2C_392_104, V2C_481_104, V2C_641_104, V2C_702_104, V2C_822_104, V2C_912_104, V2C_927_104, V2C_1006_104, V2C_1038_104, V2C_1057_104, V2C_1136_104, V2C_1255_104, V2C_1256_104, V2C_26_105, V2C_53_105, V2C_118_105, V2C_152_105, V2C_218_105, V2C_285_105, V2C_382_105, V2C_389_105, V2C_548_105, V2C_605_105, V2C_633_105, V2C_737_105, V2C_868_105, V2C_960_105, V2C_985_105, V2C_1045_105, V2C_1075_105, V2C_1120_105, V2C_1256_105, V2C_1257_105, V2C_45_106, V2C_56_106, V2C_143_106, V2C_151_106, V2C_216_106, V2C_270_106, V2C_446_106, V2C_486_106, V2C_570_106, V2C_584_106, V2C_657_106, V2C_703_106, V2C_872_106, V2C_944_106, V2C_980_106, V2C_1010_106, V2C_1085_106, V2C_1149_106, V2C_1257_106, V2C_1258_106, V2C_16_107, V2C_74_107, V2C_109_107, V2C_180_107, V2C_196_107, V2C_262_107, V2C_311_107, V2C_378_107, V2C_457_107, V2C_691_107, V2C_755_107, V2C_809_107, V2C_887_107, V2C_935_107, V2C_978_107, V2C_1030_107, V2C_1079_107, V2C_1127_107, V2C_1258_107, V2C_1259_107, V2C_47_108, V2C_71_108, V2C_111_108, V2C_179_108, V2C_213_108, V2C_244_108, V2C_297_108, V2C_449_108, V2C_546_108, V2C_579_108, V2C_783_108, V2C_859_108, V2C_892_108, V2C_954_108, V2C_989_108, V2C_1056_108, V2C_1072_108, V2C_1122_108, V2C_1259_108, V2C_1260_108, V2C_23_109, V2C_59_109, V2C_127_109, V2C_188_109, V2C_202_109, V2C_245_109, V2C_345_109, V2C_399_109, V2C_496_109, V2C_732_109, V2C_780_109, V2C_828_109, V2C_869_109, V2C_958_109, V2C_992_109, V2C_1031_109, V2C_1057_109, V2C_1116_109, V2C_1260_109, V2C_1261_109, V2C_32_110, V2C_81_110, V2C_137_110, V2C_185_110, V2C_214_110, V2C_283_110, V2C_334_110, V2C_393_110, V2C_482_110, V2C_642_110, V2C_703_110, V2C_823_110, V2C_865_110, V2C_928_110, V2C_1007_110, V2C_1039_110, V2C_1058_110, V2C_1137_110, V2C_1261_110, V2C_1262_110, V2C_27_111, V2C_54_111, V2C_119_111, V2C_153_111, V2C_219_111, V2C_286_111, V2C_383_111, V2C_390_111, V2C_549_111, V2C_606_111, V2C_634_111, V2C_738_111, V2C_869_111, V2C_913_111, V2C_986_111, V2C_1046_111, V2C_1076_111, V2C_1121_111, V2C_1262_111, V2C_1263_111, V2C_46_112, V2C_57_112, V2C_144_112, V2C_152_112, V2C_217_112, V2C_271_112, V2C_447_112, V2C_487_112, V2C_571_112, V2C_585_112, V2C_658_112, V2C_704_112, V2C_873_112, V2C_945_112, V2C_981_112, V2C_1011_112, V2C_1086_112, V2C_1150_112, V2C_1263_112, V2C_1264_112, V2C_17_113, V2C_75_113, V2C_110_113, V2C_181_113, V2C_197_113, V2C_263_113, V2C_312_113, V2C_379_113, V2C_458_113, V2C_692_113, V2C_756_113, V2C_810_113, V2C_888_113, V2C_936_113, V2C_979_113, V2C_1031_113, V2C_1080_113, V2C_1128_113, V2C_1264_113, V2C_1265_113, V2C_48_114, V2C_72_114, V2C_112_114, V2C_180_114, V2C_214_114, V2C_245_114, V2C_298_114, V2C_450_114, V2C_547_114, V2C_580_114, V2C_784_114, V2C_860_114, V2C_893_114, V2C_955_114, V2C_990_114, V2C_1009_114, V2C_1073_114, V2C_1123_114, V2C_1265_114, V2C_1266_114, V2C_24_115, V2C_60_115, V2C_128_115, V2C_189_115, V2C_203_115, V2C_246_115, V2C_346_115, V2C_400_115, V2C_497_115, V2C_733_115, V2C_781_115, V2C_829_115, V2C_870_115, V2C_959_115, V2C_993_115, V2C_1032_115, V2C_1058_115, V2C_1117_115, V2C_1266_115, V2C_1267_115, V2C_33_116, V2C_82_116, V2C_138_116, V2C_186_116, V2C_215_116, V2C_284_116, V2C_335_116, V2C_394_116, V2C_483_116, V2C_643_116, V2C_704_116, V2C_824_116, V2C_866_116, V2C_929_116, V2C_1008_116, V2C_1040_116, V2C_1059_116, V2C_1138_116, V2C_1267_116, V2C_1268_116, V2C_28_117, V2C_55_117, V2C_120_117, V2C_154_117, V2C_220_117, V2C_287_117, V2C_384_117, V2C_391_117, V2C_550_117, V2C_607_117, V2C_635_117, V2C_739_117, V2C_870_117, V2C_914_117, V2C_987_117, V2C_1047_117, V2C_1077_117, V2C_1122_117, V2C_1268_117, V2C_1269_117, V2C_47_118, V2C_58_118, V2C_97_118, V2C_153_118, V2C_218_118, V2C_272_118, V2C_448_118, V2C_488_118, V2C_572_118, V2C_586_118, V2C_659_118, V2C_705_118, V2C_874_118, V2C_946_118, V2C_982_118, V2C_1012_118, V2C_1087_118, V2C_1151_118, V2C_1269_118, V2C_1270_118, V2C_18_119, V2C_76_119, V2C_111_119, V2C_182_119, V2C_198_119, V2C_264_119, V2C_313_119, V2C_380_119, V2C_459_119, V2C_693_119, V2C_757_119, V2C_811_119, V2C_889_119, V2C_937_119, V2C_980_119, V2C_1032_119, V2C_1081_119, V2C_1129_119, V2C_1270_119, V2C_1271_119, V2C_1_120, V2C_73_120, V2C_113_120, V2C_181_120, V2C_215_120, V2C_246_120, V2C_299_120, V2C_451_120, V2C_548_120, V2C_581_120, V2C_785_120, V2C_861_120, V2C_894_120, V2C_956_120, V2C_991_120, V2C_1010_120, V2C_1074_120, V2C_1124_120, V2C_1271_120, V2C_1272_120, V2C_25_121, V2C_61_121, V2C_129_121, V2C_190_121, V2C_204_121, V2C_247_121, V2C_347_121, V2C_401_121, V2C_498_121, V2C_734_121, V2C_782_121, V2C_830_121, V2C_871_121, V2C_960_121, V2C_994_121, V2C_1033_121, V2C_1059_121, V2C_1118_121, V2C_1272_121, V2C_1273_121, V2C_34_122, V2C_83_122, V2C_139_122, V2C_187_122, V2C_216_122, V2C_285_122, V2C_336_122, V2C_395_122, V2C_484_122, V2C_644_122, V2C_705_122, V2C_825_122, V2C_867_122, V2C_930_122, V2C_961_122, V2C_1041_122, V2C_1060_122, V2C_1139_122, V2C_1273_122, V2C_1274_122, V2C_29_123, V2C_56_123, V2C_121_123, V2C_155_123, V2C_221_123, V2C_288_123, V2C_337_123, V2C_392_123, V2C_551_123, V2C_608_123, V2C_636_123, V2C_740_123, V2C_871_123, V2C_915_123, V2C_988_123, V2C_1048_123, V2C_1078_123, V2C_1123_123, V2C_1274_123, V2C_1275_123, V2C_48_124, V2C_59_124, V2C_98_124, V2C_154_124, V2C_219_124, V2C_273_124, V2C_449_124, V2C_489_124, V2C_573_124, V2C_587_124, V2C_660_124, V2C_706_124, V2C_875_124, V2C_947_124, V2C_983_124, V2C_1013_124, V2C_1088_124, V2C_1152_124, V2C_1275_124, V2C_1276_124, V2C_19_125, V2C_77_125, V2C_112_125, V2C_183_125, V2C_199_125, V2C_265_125, V2C_314_125, V2C_381_125, V2C_460_125, V2C_694_125, V2C_758_125, V2C_812_125, V2C_890_125, V2C_938_125, V2C_981_125, V2C_1033_125, V2C_1082_125, V2C_1130_125, V2C_1276_125, V2C_1277_125, V2C_2_126, V2C_74_126, V2C_114_126, V2C_182_126, V2C_216_126, V2C_247_126, V2C_300_126, V2C_452_126, V2C_549_126, V2C_582_126, V2C_786_126, V2C_862_126, V2C_895_126, V2C_957_126, V2C_992_126, V2C_1011_126, V2C_1075_126, V2C_1125_126, V2C_1277_126, V2C_1278_126, V2C_26_127, V2C_62_127, V2C_130_127, V2C_191_127, V2C_205_127, V2C_248_127, V2C_348_127, V2C_402_127, V2C_499_127, V2C_735_127, V2C_783_127, V2C_831_127, V2C_872_127, V2C_913_127, V2C_995_127, V2C_1034_127, V2C_1060_127, V2C_1119_127, V2C_1278_127, V2C_1279_127, V2C_35_128, V2C_84_128, V2C_140_128, V2C_188_128, V2C_217_128, V2C_286_128, V2C_289_128, V2C_396_128, V2C_485_128, V2C_645_128, V2C_706_128, V2C_826_128, V2C_868_128, V2C_931_128, V2C_962_128, V2C_1042_128, V2C_1061_128, V2C_1140_128, V2C_1279_128, V2C_1280_128, V2C_30_129, V2C_57_129, V2C_122_129, V2C_156_129, V2C_222_129, V2C_241_129, V2C_338_129, V2C_393_129, V2C_552_129, V2C_609_129, V2C_637_129, V2C_741_129, V2C_872_129, V2C_916_129, V2C_989_129, V2C_1049_129, V2C_1079_129, V2C_1124_129, V2C_1280_129, V2C_1281_129, V2C_1_130, V2C_60_130, V2C_99_130, V2C_155_130, V2C_220_130, V2C_274_130, V2C_450_130, V2C_490_130, V2C_574_130, V2C_588_130, V2C_661_130, V2C_707_130, V2C_876_130, V2C_948_130, V2C_984_130, V2C_1014_130, V2C_1089_130, V2C_1105_130, V2C_1281_130, V2C_1282_130, V2C_20_131, V2C_78_131, V2C_113_131, V2C_184_131, V2C_200_131, V2C_266_131, V2C_315_131, V2C_382_131, V2C_461_131, V2C_695_131, V2C_759_131, V2C_813_131, V2C_891_131, V2C_939_131, V2C_982_131, V2C_1034_131, V2C_1083_131, V2C_1131_131, V2C_1282_131, V2C_1283_131, V2C_3_132, V2C_75_132, V2C_115_132, V2C_183_132, V2C_217_132, V2C_248_132, V2C_301_132, V2C_453_132, V2C_550_132, V2C_583_132, V2C_787_132, V2C_863_132, V2C_896_132, V2C_958_132, V2C_993_132, V2C_1012_132, V2C_1076_132, V2C_1126_132, V2C_1283_132, V2C_1284_132, V2C_27_133, V2C_63_133, V2C_131_133, V2C_192_133, V2C_206_133, V2C_249_133, V2C_349_133, V2C_403_133, V2C_500_133, V2C_736_133, V2C_784_133, V2C_832_133, V2C_873_133, V2C_914_133, V2C_996_133, V2C_1035_133, V2C_1061_133, V2C_1120_133, V2C_1284_133, V2C_1285_133, V2C_36_134, V2C_85_134, V2C_141_134, V2C_189_134, V2C_218_134, V2C_287_134, V2C_290_134, V2C_397_134, V2C_486_134, V2C_646_134, V2C_707_134, V2C_827_134, V2C_869_134, V2C_932_134, V2C_963_134, V2C_1043_134, V2C_1062_134, V2C_1141_134, V2C_1285_134, V2C_1286_134, V2C_31_135, V2C_58_135, V2C_123_135, V2C_157_135, V2C_223_135, V2C_242_135, V2C_339_135, V2C_394_135, V2C_553_135, V2C_610_135, V2C_638_135, V2C_742_135, V2C_873_135, V2C_917_135, V2C_990_135, V2C_1050_135, V2C_1080_135, V2C_1125_135, V2C_1286_135, V2C_1287_135, V2C_2_136, V2C_61_136, V2C_100_136, V2C_156_136, V2C_221_136, V2C_275_136, V2C_451_136, V2C_491_136, V2C_575_136, V2C_589_136, V2C_662_136, V2C_708_136, V2C_877_136, V2C_949_136, V2C_985_136, V2C_1015_136, V2C_1090_136, V2C_1106_136, V2C_1287_136, V2C_1288_136, V2C_21_137, V2C_79_137, V2C_114_137, V2C_185_137, V2C_201_137, V2C_267_137, V2C_316_137, V2C_383_137, V2C_462_137, V2C_696_137, V2C_760_137, V2C_814_137, V2C_892_137, V2C_940_137, V2C_983_137, V2C_1035_137, V2C_1084_137, V2C_1132_137, V2C_1288_137, V2C_1289_137, V2C_4_138, V2C_76_138, V2C_116_138, V2C_184_138, V2C_218_138, V2C_249_138, V2C_302_138, V2C_454_138, V2C_551_138, V2C_584_138, V2C_788_138, V2C_864_138, V2C_897_138, V2C_959_138, V2C_994_138, V2C_1013_138, V2C_1077_138, V2C_1127_138, V2C_1289_138, V2C_1290_138, V2C_28_139, V2C_64_139, V2C_132_139, V2C_145_139, V2C_207_139, V2C_250_139, V2C_350_139, V2C_404_139, V2C_501_139, V2C_737_139, V2C_785_139, V2C_833_139, V2C_874_139, V2C_915_139, V2C_997_139, V2C_1036_139, V2C_1062_139, V2C_1121_139, V2C_1290_139, V2C_1291_139, V2C_37_140, V2C_86_140, V2C_142_140, V2C_190_140, V2C_219_140, V2C_288_140, V2C_291_140, V2C_398_140, V2C_487_140, V2C_647_140, V2C_708_140, V2C_828_140, V2C_870_140, V2C_933_140, V2C_964_140, V2C_1044_140, V2C_1063_140, V2C_1142_140, V2C_1291_140, V2C_1292_140, V2C_32_141, V2C_59_141, V2C_124_141, V2C_158_141, V2C_224_141, V2C_243_141, V2C_340_141, V2C_395_141, V2C_554_141, V2C_611_141, V2C_639_141, V2C_743_141, V2C_874_141, V2C_918_141, V2C_991_141, V2C_1051_141, V2C_1081_141, V2C_1126_141, V2C_1292_141, V2C_1293_141, V2C_3_142, V2C_62_142, V2C_101_142, V2C_157_142, V2C_222_142, V2C_276_142, V2C_452_142, V2C_492_142, V2C_576_142, V2C_590_142, V2C_663_142, V2C_709_142, V2C_878_142, V2C_950_142, V2C_986_142, V2C_1016_142, V2C_1091_142, V2C_1107_142, V2C_1293_142, V2C_1294_142, V2C_22_143, V2C_80_143, V2C_115_143, V2C_186_143, V2C_202_143, V2C_268_143, V2C_317_143, V2C_384_143, V2C_463_143, V2C_697_143, V2C_761_143, V2C_815_143, V2C_893_143, V2C_941_143, V2C_984_143, V2C_1036_143, V2C_1085_143, V2C_1133_143, V2C_1294_143, V2C_1295_143, V2C_5_144, V2C_77_144, V2C_117_144, V2C_185_144, V2C_219_144, V2C_250_144, V2C_303_144, V2C_455_144, V2C_552_144, V2C_585_144, V2C_789_144, V2C_817_144, V2C_898_144, V2C_960_144, V2C_995_144, V2C_1014_144, V2C_1078_144, V2C_1128_144, V2C_1295_144, V2C_1296_144, V2C_29_145, V2C_65_145, V2C_133_145, V2C_146_145, V2C_208_145, V2C_251_145, V2C_351_145, V2C_405_145, V2C_502_145, V2C_738_145, V2C_786_145, V2C_834_145, V2C_875_145, V2C_916_145, V2C_998_145, V2C_1037_145, V2C_1063_145, V2C_1122_145, V2C_1296_145, V2C_1297_145, V2C_38_146, V2C_87_146, V2C_143_146, V2C_191_146, V2C_220_146, V2C_241_146, V2C_292_146, V2C_399_146, V2C_488_146, V2C_648_146, V2C_709_146, V2C_829_146, V2C_871_146, V2C_934_146, V2C_965_146, V2C_1045_146, V2C_1064_146, V2C_1143_146, V2C_1297_146, V2C_1298_146, V2C_33_147, V2C_60_147, V2C_125_147, V2C_159_147, V2C_225_147, V2C_244_147, V2C_341_147, V2C_396_147, V2C_555_147, V2C_612_147, V2C_640_147, V2C_744_147, V2C_875_147, V2C_919_147, V2C_992_147, V2C_1052_147, V2C_1082_147, V2C_1127_147, V2C_1298_147, V2C_1299_147, V2C_4_148, V2C_63_148, V2C_102_148, V2C_158_148, V2C_223_148, V2C_277_148, V2C_453_148, V2C_493_148, V2C_529_148, V2C_591_148, V2C_664_148, V2C_710_148, V2C_879_148, V2C_951_148, V2C_987_148, V2C_1017_148, V2C_1092_148, V2C_1108_148, V2C_1299_148, V2C_1300_148, V2C_23_149, V2C_81_149, V2C_116_149, V2C_187_149, V2C_203_149, V2C_269_149, V2C_318_149, V2C_337_149, V2C_464_149, V2C_698_149, V2C_762_149, V2C_816_149, V2C_894_149, V2C_942_149, V2C_985_149, V2C_1037_149, V2C_1086_149, V2C_1134_149, V2C_1300_149, V2C_1301_149, V2C_6_150, V2C_78_150, V2C_118_150, V2C_186_150, V2C_220_150, V2C_251_150, V2C_304_150, V2C_456_150, V2C_553_150, V2C_586_150, V2C_790_150, V2C_818_150, V2C_899_150, V2C_913_150, V2C_996_150, V2C_1015_150, V2C_1079_150, V2C_1129_150, V2C_1301_150, V2C_1302_150, V2C_30_151, V2C_66_151, V2C_134_151, V2C_147_151, V2C_209_151, V2C_252_151, V2C_352_151, V2C_406_151, V2C_503_151, V2C_739_151, V2C_787_151, V2C_835_151, V2C_876_151, V2C_917_151, V2C_999_151, V2C_1038_151, V2C_1064_151, V2C_1123_151, V2C_1302_151, V2C_1303_151, V2C_39_152, V2C_88_152, V2C_144_152, V2C_192_152, V2C_221_152, V2C_242_152, V2C_293_152, V2C_400_152, V2C_489_152, V2C_649_152, V2C_710_152, V2C_830_152, V2C_872_152, V2C_935_152, V2C_966_152, V2C_1046_152, V2C_1065_152, V2C_1144_152, V2C_1303_152, V2C_1304_152, V2C_34_153, V2C_61_153, V2C_126_153, V2C_160_153, V2C_226_153, V2C_245_153, V2C_342_153, V2C_397_153, V2C_556_153, V2C_613_153, V2C_641_153, V2C_745_153, V2C_876_153, V2C_920_153, V2C_993_153, V2C_1053_153, V2C_1083_153, V2C_1128_153, V2C_1304_153, V2C_1305_153, V2C_5_154, V2C_64_154, V2C_103_154, V2C_159_154, V2C_224_154, V2C_278_154, V2C_454_154, V2C_494_154, V2C_530_154, V2C_592_154, V2C_665_154, V2C_711_154, V2C_880_154, V2C_952_154, V2C_988_154, V2C_1018_154, V2C_1093_154, V2C_1109_154, V2C_1305_154, V2C_1306_154, V2C_24_155, V2C_82_155, V2C_117_155, V2C_188_155, V2C_204_155, V2C_270_155, V2C_319_155, V2C_338_155, V2C_465_155, V2C_699_155, V2C_763_155, V2C_769_155, V2C_895_155, V2C_943_155, V2C_986_155, V2C_1038_155, V2C_1087_155, V2C_1135_155, V2C_1306_155, V2C_1307_155, V2C_7_156, V2C_79_156, V2C_119_156, V2C_187_156, V2C_221_156, V2C_252_156, V2C_305_156, V2C_457_156, V2C_554_156, V2C_587_156, V2C_791_156, V2C_819_156, V2C_900_156, V2C_914_156, V2C_997_156, V2C_1016_156, V2C_1080_156, V2C_1130_156, V2C_1307_156, V2C_1308_156, V2C_31_157, V2C_67_157, V2C_135_157, V2C_148_157, V2C_210_157, V2C_253_157, V2C_353_157, V2C_407_157, V2C_504_157, V2C_740_157, V2C_788_157, V2C_836_157, V2C_877_157, V2C_918_157, V2C_1000_157, V2C_1039_157, V2C_1065_157, V2C_1124_157, V2C_1308_157, V2C_1309_157, V2C_40_158, V2C_89_158, V2C_97_158, V2C_145_158, V2C_222_158, V2C_243_158, V2C_294_158, V2C_401_158, V2C_490_158, V2C_650_158, V2C_711_158, V2C_831_158, V2C_873_158, V2C_936_158, V2C_967_158, V2C_1047_158, V2C_1066_158, V2C_1145_158, V2C_1309_158, V2C_1310_158, V2C_35_159, V2C_62_159, V2C_127_159, V2C_161_159, V2C_227_159, V2C_246_159, V2C_343_159, V2C_398_159, V2C_557_159, V2C_614_159, V2C_642_159, V2C_746_159, V2C_877_159, V2C_921_159, V2C_994_159, V2C_1054_159, V2C_1084_159, V2C_1129_159, V2C_1310_159, V2C_1311_159, V2C_6_160, V2C_65_160, V2C_104_160, V2C_160_160, V2C_225_160, V2C_279_160, V2C_455_160, V2C_495_160, V2C_531_160, V2C_593_160, V2C_666_160, V2C_712_160, V2C_881_160, V2C_953_160, V2C_989_160, V2C_1019_160, V2C_1094_160, V2C_1110_160, V2C_1311_160, V2C_1312_160, V2C_25_161, V2C_83_161, V2C_118_161, V2C_189_161, V2C_205_161, V2C_271_161, V2C_320_161, V2C_339_161, V2C_466_161, V2C_700_161, V2C_764_161, V2C_770_161, V2C_896_161, V2C_944_161, V2C_987_161, V2C_1039_161, V2C_1088_161, V2C_1136_161, V2C_1312_161, V2C_1313_161, V2C_8_162, V2C_80_162, V2C_120_162, V2C_188_162, V2C_222_162, V2C_253_162, V2C_306_162, V2C_458_162, V2C_555_162, V2C_588_162, V2C_792_162, V2C_820_162, V2C_901_162, V2C_915_162, V2C_998_162, V2C_1017_162, V2C_1081_162, V2C_1131_162, V2C_1313_162, V2C_1314_162, V2C_32_163, V2C_68_163, V2C_136_163, V2C_149_163, V2C_211_163, V2C_254_163, V2C_354_163, V2C_408_163, V2C_505_163, V2C_741_163, V2C_789_163, V2C_837_163, V2C_878_163, V2C_919_163, V2C_1001_163, V2C_1040_163, V2C_1066_163, V2C_1125_163, V2C_1314_163, V2C_1315_163, V2C_41_164, V2C_90_164, V2C_98_164, V2C_146_164, V2C_223_164, V2C_244_164, V2C_295_164, V2C_402_164, V2C_491_164, V2C_651_164, V2C_712_164, V2C_832_164, V2C_874_164, V2C_937_164, V2C_968_164, V2C_1048_164, V2C_1067_164, V2C_1146_164, V2C_1315_164, V2C_1316_164, V2C_36_165, V2C_63_165, V2C_128_165, V2C_162_165, V2C_228_165, V2C_247_165, V2C_344_165, V2C_399_165, V2C_558_165, V2C_615_165, V2C_643_165, V2C_747_165, V2C_878_165, V2C_922_165, V2C_995_165, V2C_1055_165, V2C_1085_165, V2C_1130_165, V2C_1316_165, V2C_1317_165, V2C_7_166, V2C_66_166, V2C_105_166, V2C_161_166, V2C_226_166, V2C_280_166, V2C_456_166, V2C_496_166, V2C_532_166, V2C_594_166, V2C_667_166, V2C_713_166, V2C_882_166, V2C_954_166, V2C_990_166, V2C_1020_166, V2C_1095_166, V2C_1111_166, V2C_1317_166, V2C_1318_166, V2C_26_167, V2C_84_167, V2C_119_167, V2C_190_167, V2C_206_167, V2C_272_167, V2C_321_167, V2C_340_167, V2C_467_167, V2C_701_167, V2C_765_167, V2C_771_167, V2C_897_167, V2C_945_167, V2C_988_167, V2C_1040_167, V2C_1089_167, V2C_1137_167, V2C_1318_167, V2C_1319_167, V2C_9_168, V2C_81_168, V2C_121_168, V2C_189_168, V2C_223_168, V2C_254_168, V2C_307_168, V2C_459_168, V2C_556_168, V2C_589_168, V2C_793_168, V2C_821_168, V2C_902_168, V2C_916_168, V2C_999_168, V2C_1018_168, V2C_1082_168, V2C_1132_168, V2C_1319_168, V2C_1320_168, V2C_33_169, V2C_69_169, V2C_137_169, V2C_150_169, V2C_212_169, V2C_255_169, V2C_355_169, V2C_409_169, V2C_506_169, V2C_742_169, V2C_790_169, V2C_838_169, V2C_879_169, V2C_920_169, V2C_1002_169, V2C_1041_169, V2C_1067_169, V2C_1126_169, V2C_1320_169, V2C_1321_169, V2C_42_170, V2C_91_170, V2C_99_170, V2C_147_170, V2C_224_170, V2C_245_170, V2C_296_170, V2C_403_170, V2C_492_170, V2C_652_170, V2C_713_170, V2C_833_170, V2C_875_170, V2C_938_170, V2C_969_170, V2C_1049_170, V2C_1068_170, V2C_1147_170, V2C_1321_170, V2C_1322_170, V2C_37_171, V2C_64_171, V2C_129_171, V2C_163_171, V2C_229_171, V2C_248_171, V2C_345_171, V2C_400_171, V2C_559_171, V2C_616_171, V2C_644_171, V2C_748_171, V2C_879_171, V2C_923_171, V2C_996_171, V2C_1056_171, V2C_1086_171, V2C_1131_171, V2C_1322_171, V2C_1323_171, V2C_8_172, V2C_67_172, V2C_106_172, V2C_162_172, V2C_227_172, V2C_281_172, V2C_457_172, V2C_497_172, V2C_533_172, V2C_595_172, V2C_668_172, V2C_714_172, V2C_883_172, V2C_955_172, V2C_991_172, V2C_1021_172, V2C_1096_172, V2C_1112_172, V2C_1323_172, V2C_1324_172, V2C_27_173, V2C_85_173, V2C_120_173, V2C_191_173, V2C_207_173, V2C_273_173, V2C_322_173, V2C_341_173, V2C_468_173, V2C_702_173, V2C_766_173, V2C_772_173, V2C_898_173, V2C_946_173, V2C_989_173, V2C_1041_173, V2C_1090_173, V2C_1138_173, V2C_1324_173, V2C_1325_173, V2C_10_174, V2C_82_174, V2C_122_174, V2C_190_174, V2C_224_174, V2C_255_174, V2C_308_174, V2C_460_174, V2C_557_174, V2C_590_174, V2C_794_174, V2C_822_174, V2C_903_174, V2C_917_174, V2C_1000_174, V2C_1019_174, V2C_1083_174, V2C_1133_174, V2C_1325_174, V2C_1326_174, V2C_34_175, V2C_70_175, V2C_138_175, V2C_151_175, V2C_213_175, V2C_256_175, V2C_356_175, V2C_410_175, V2C_507_175, V2C_743_175, V2C_791_175, V2C_839_175, V2C_880_175, V2C_921_175, V2C_1003_175, V2C_1042_175, V2C_1068_175, V2C_1127_175, V2C_1326_175, V2C_1327_175, V2C_43_176, V2C_92_176, V2C_100_176, V2C_148_176, V2C_225_176, V2C_246_176, V2C_297_176, V2C_404_176, V2C_493_176, V2C_653_176, V2C_714_176, V2C_834_176, V2C_876_176, V2C_939_176, V2C_970_176, V2C_1050_176, V2C_1069_176, V2C_1148_176, V2C_1327_176, V2C_1328_176, V2C_38_177, V2C_65_177, V2C_130_177, V2C_164_177, V2C_230_177, V2C_249_177, V2C_346_177, V2C_401_177, V2C_560_177, V2C_617_177, V2C_645_177, V2C_749_177, V2C_880_177, V2C_924_177, V2C_997_177, V2C_1009_177, V2C_1087_177, V2C_1132_177, V2C_1328_177, V2C_1329_177, V2C_9_178, V2C_68_178, V2C_107_178, V2C_163_178, V2C_228_178, V2C_282_178, V2C_458_178, V2C_498_178, V2C_534_178, V2C_596_178, V2C_669_178, V2C_715_178, V2C_884_178, V2C_956_178, V2C_992_178, V2C_1022_178, V2C_1097_178, V2C_1113_178, V2C_1329_178, V2C_1330_178, V2C_28_179, V2C_86_179, V2C_121_179, V2C_192_179, V2C_208_179, V2C_274_179, V2C_323_179, V2C_342_179, V2C_469_179, V2C_703_179, V2C_767_179, V2C_773_179, V2C_899_179, V2C_947_179, V2C_990_179, V2C_1042_179, V2C_1091_179, V2C_1139_179, V2C_1330_179, V2C_1331_179, V2C_11_180, V2C_83_180, V2C_123_180, V2C_191_180, V2C_225_180, V2C_256_180, V2C_309_180, V2C_461_180, V2C_558_180, V2C_591_180, V2C_795_180, V2C_823_180, V2C_904_180, V2C_918_180, V2C_1001_180, V2C_1020_180, V2C_1084_180, V2C_1134_180, V2C_1331_180, V2C_1332_180, V2C_35_181, V2C_71_181, V2C_139_181, V2C_152_181, V2C_214_181, V2C_257_181, V2C_357_181, V2C_411_181, V2C_508_181, V2C_744_181, V2C_792_181, V2C_840_181, V2C_881_181, V2C_922_181, V2C_1004_181, V2C_1043_181, V2C_1069_181, V2C_1128_181, V2C_1332_181, V2C_1333_181, V2C_44_182, V2C_93_182, V2C_101_182, V2C_149_182, V2C_226_182, V2C_247_182, V2C_298_182, V2C_405_182, V2C_494_182, V2C_654_182, V2C_715_182, V2C_835_182, V2C_877_182, V2C_940_182, V2C_971_182, V2C_1051_182, V2C_1070_182, V2C_1149_182, V2C_1333_182, V2C_1334_182, V2C_39_183, V2C_66_183, V2C_131_183, V2C_165_183, V2C_231_183, V2C_250_183, V2C_347_183, V2C_402_183, V2C_561_183, V2C_618_183, V2C_646_183, V2C_750_183, V2C_881_183, V2C_925_183, V2C_998_183, V2C_1010_183, V2C_1088_183, V2C_1133_183, V2C_1334_183, V2C_1335_183, V2C_10_184, V2C_69_184, V2C_108_184, V2C_164_184, V2C_229_184, V2C_283_184, V2C_459_184, V2C_499_184, V2C_535_184, V2C_597_184, V2C_670_184, V2C_716_184, V2C_885_184, V2C_957_184, V2C_993_184, V2C_1023_184, V2C_1098_184, V2C_1114_184, V2C_1335_184, V2C_1336_184, V2C_29_185, V2C_87_185, V2C_122_185, V2C_145_185, V2C_209_185, V2C_275_185, V2C_324_185, V2C_343_185, V2C_470_185, V2C_704_185, V2C_768_185, V2C_774_185, V2C_900_185, V2C_948_185, V2C_991_185, V2C_1043_185, V2C_1092_185, V2C_1140_185, V2C_1336_185, V2C_1337_185, V2C_12_186, V2C_84_186, V2C_124_186, V2C_192_186, V2C_226_186, V2C_257_186, V2C_310_186, V2C_462_186, V2C_559_186, V2C_592_186, V2C_796_186, V2C_824_186, V2C_905_186, V2C_919_186, V2C_1002_186, V2C_1021_186, V2C_1085_186, V2C_1135_186, V2C_1337_186, V2C_1338_186, V2C_36_187, V2C_72_187, V2C_140_187, V2C_153_187, V2C_215_187, V2C_258_187, V2C_358_187, V2C_412_187, V2C_509_187, V2C_745_187, V2C_793_187, V2C_841_187, V2C_882_187, V2C_923_187, V2C_1005_187, V2C_1044_187, V2C_1070_187, V2C_1129_187, V2C_1338_187, V2C_1339_187, V2C_45_188, V2C_94_188, V2C_102_188, V2C_150_188, V2C_227_188, V2C_248_188, V2C_299_188, V2C_406_188, V2C_495_188, V2C_655_188, V2C_716_188, V2C_836_188, V2C_878_188, V2C_941_188, V2C_972_188, V2C_1052_188, V2C_1071_188, V2C_1150_188, V2C_1339_188, V2C_1340_188, V2C_40_189, V2C_67_189, V2C_132_189, V2C_166_189, V2C_232_189, V2C_251_189, V2C_348_189, V2C_403_189, V2C_562_189, V2C_619_189, V2C_647_189, V2C_751_189, V2C_882_189, V2C_926_189, V2C_999_189, V2C_1011_189, V2C_1089_189, V2C_1134_189, V2C_1340_189, V2C_1341_189, V2C_11_190, V2C_70_190, V2C_109_190, V2C_165_190, V2C_230_190, V2C_284_190, V2C_460_190, V2C_500_190, V2C_536_190, V2C_598_190, V2C_671_190, V2C_717_190, V2C_886_190, V2C_958_190, V2C_994_190, V2C_1024_190, V2C_1099_190, V2C_1115_190, V2C_1341_190, V2C_1342_190, V2C_30_191, V2C_88_191, V2C_123_191, V2C_146_191, V2C_210_191, V2C_276_191, V2C_325_191, V2C_344_191, V2C_471_191, V2C_705_191, V2C_721_191, V2C_775_191, V2C_901_191, V2C_949_191, V2C_992_191, V2C_1044_191, V2C_1093_191, V2C_1141_191, V2C_1342_191, V2C_1343_191, V2C_13_192, V2C_85_192, V2C_125_192, V2C_145_192, V2C_227_192, V2C_258_192, V2C_311_192, V2C_463_192, V2C_560_192, V2C_593_192, V2C_797_192, V2C_825_192, V2C_906_192, V2C_920_192, V2C_1003_192, V2C_1022_192, V2C_1086_192, V2C_1136_192, V2C_1343_192, V2C_1344_192, V2C_37_193, V2C_73_193, V2C_141_193, V2C_154_193, V2C_216_193, V2C_259_193, V2C_359_193, V2C_413_193, V2C_510_193, V2C_746_193, V2C_794_193, V2C_842_193, V2C_883_193, V2C_924_193, V2C_1006_193, V2C_1045_193, V2C_1071_193, V2C_1130_193, V2C_1344_193, V2C_1345_193, V2C_46_194, V2C_95_194, V2C_103_194, V2C_151_194, V2C_228_194, V2C_249_194, V2C_300_194, V2C_407_194, V2C_496_194, V2C_656_194, V2C_717_194, V2C_837_194, V2C_879_194, V2C_942_194, V2C_973_194, V2C_1053_194, V2C_1072_194, V2C_1151_194, V2C_1345_194, V2C_1346_194, V2C_41_195, V2C_68_195, V2C_133_195, V2C_167_195, V2C_233_195, V2C_252_195, V2C_349_195, V2C_404_195, V2C_563_195, V2C_620_195, V2C_648_195, V2C_752_195, V2C_883_195, V2C_927_195, V2C_1000_195, V2C_1012_195, V2C_1090_195, V2C_1135_195, V2C_1346_195, V2C_1347_195, V2C_12_196, V2C_71_196, V2C_110_196, V2C_166_196, V2C_231_196, V2C_285_196, V2C_461_196, V2C_501_196, V2C_537_196, V2C_599_196, V2C_672_196, V2C_718_196, V2C_887_196, V2C_959_196, V2C_995_196, V2C_1025_196, V2C_1100_196, V2C_1116_196, V2C_1347_196, V2C_1348_196, V2C_31_197, V2C_89_197, V2C_124_197, V2C_147_197, V2C_211_197, V2C_277_197, V2C_326_197, V2C_345_197, V2C_472_197, V2C_706_197, V2C_722_197, V2C_776_197, V2C_902_197, V2C_950_197, V2C_993_197, V2C_1045_197, V2C_1094_197, V2C_1142_197, V2C_1348_197, V2C_1349_197, V2C_14_198, V2C_86_198, V2C_126_198, V2C_146_198, V2C_228_198, V2C_259_198, V2C_312_198, V2C_464_198, V2C_561_198, V2C_594_198, V2C_798_198, V2C_826_198, V2C_907_198, V2C_921_198, V2C_1004_198, V2C_1023_198, V2C_1087_198, V2C_1137_198, V2C_1349_198, V2C_1350_198, V2C_38_199, V2C_74_199, V2C_142_199, V2C_155_199, V2C_217_199, V2C_260_199, V2C_360_199, V2C_414_199, V2C_511_199, V2C_747_199, V2C_795_199, V2C_843_199, V2C_884_199, V2C_925_199, V2C_1007_199, V2C_1046_199, V2C_1072_199, V2C_1131_199, V2C_1350_199, V2C_1351_199, V2C_47_200, V2C_96_200, V2C_104_200, V2C_152_200, V2C_229_200, V2C_250_200, V2C_301_200, V2C_408_200, V2C_497_200, V2C_657_200, V2C_718_200, V2C_838_200, V2C_880_200, V2C_943_200, V2C_974_200, V2C_1054_200, V2C_1073_200, V2C_1152_200, V2C_1351_200, V2C_1352_200, V2C_42_201, V2C_69_201, V2C_134_201, V2C_168_201, V2C_234_201, V2C_253_201, V2C_350_201, V2C_405_201, V2C_564_201, V2C_621_201, V2C_649_201, V2C_753_201, V2C_884_201, V2C_928_201, V2C_1001_201, V2C_1013_201, V2C_1091_201, V2C_1136_201, V2C_1352_201, V2C_1353_201, V2C_13_202, V2C_72_202, V2C_111_202, V2C_167_202, V2C_232_202, V2C_286_202, V2C_462_202, V2C_502_202, V2C_538_202, V2C_600_202, V2C_625_202, V2C_719_202, V2C_888_202, V2C_960_202, V2C_996_202, V2C_1026_202, V2C_1101_202, V2C_1117_202, V2C_1353_202, V2C_1354_202, V2C_32_203, V2C_90_203, V2C_125_203, V2C_148_203, V2C_212_203, V2C_278_203, V2C_327_203, V2C_346_203, V2C_473_203, V2C_707_203, V2C_723_203, V2C_777_203, V2C_903_203, V2C_951_203, V2C_994_203, V2C_1046_203, V2C_1095_203, V2C_1143_203, V2C_1354_203, V2C_1355_203, V2C_15_204, V2C_87_204, V2C_127_204, V2C_147_204, V2C_229_204, V2C_260_204, V2C_313_204, V2C_465_204, V2C_562_204, V2C_595_204, V2C_799_204, V2C_827_204, V2C_908_204, V2C_922_204, V2C_1005_204, V2C_1024_204, V2C_1088_204, V2C_1138_204, V2C_1355_204, V2C_1356_204, V2C_39_205, V2C_75_205, V2C_143_205, V2C_156_205, V2C_218_205, V2C_261_205, V2C_361_205, V2C_415_205, V2C_512_205, V2C_748_205, V2C_796_205, V2C_844_205, V2C_885_205, V2C_926_205, V2C_1008_205, V2C_1047_205, V2C_1073_205, V2C_1132_205, V2C_1356_205, V2C_1357_205, V2C_48_206, V2C_49_206, V2C_105_206, V2C_153_206, V2C_230_206, V2C_251_206, V2C_302_206, V2C_409_206, V2C_498_206, V2C_658_206, V2C_719_206, V2C_839_206, V2C_881_206, V2C_944_206, V2C_975_206, V2C_1055_206, V2C_1074_206, V2C_1105_206, V2C_1357_206, V2C_1358_206, V2C_43_207, V2C_70_207, V2C_135_207, V2C_169_207, V2C_235_207, V2C_254_207, V2C_351_207, V2C_406_207, V2C_565_207, V2C_622_207, V2C_650_207, V2C_754_207, V2C_885_207, V2C_929_207, V2C_1002_207, V2C_1014_207, V2C_1092_207, V2C_1137_207, V2C_1358_207, V2C_1359_207, V2C_14_208, V2C_73_208, V2C_112_208, V2C_168_208, V2C_233_208, V2C_287_208, V2C_463_208, V2C_503_208, V2C_539_208, V2C_601_208, V2C_626_208, V2C_720_208, V2C_889_208, V2C_913_208, V2C_997_208, V2C_1027_208, V2C_1102_208, V2C_1118_208, V2C_1359_208, V2C_1360_208, V2C_33_209, V2C_91_209, V2C_126_209, V2C_149_209, V2C_213_209, V2C_279_209, V2C_328_209, V2C_347_209, V2C_474_209, V2C_708_209, V2C_724_209, V2C_778_209, V2C_904_209, V2C_952_209, V2C_995_209, V2C_1047_209, V2C_1096_209, V2C_1144_209, V2C_1360_209, V2C_1361_209, V2C_16_210, V2C_88_210, V2C_128_210, V2C_148_210, V2C_230_210, V2C_261_210, V2C_314_210, V2C_466_210, V2C_563_210, V2C_596_210, V2C_800_210, V2C_828_210, V2C_909_210, V2C_923_210, V2C_1006_210, V2C_1025_210, V2C_1089_210, V2C_1139_210, V2C_1361_210, V2C_1362_210, V2C_40_211, V2C_76_211, V2C_144_211, V2C_157_211, V2C_219_211, V2C_262_211, V2C_362_211, V2C_416_211, V2C_513_211, V2C_749_211, V2C_797_211, V2C_845_211, V2C_886_211, V2C_927_211, V2C_961_211, V2C_1048_211, V2C_1074_211, V2C_1133_211, V2C_1362_211, V2C_1363_211, V2C_1_212, V2C_50_212, V2C_106_212, V2C_154_212, V2C_231_212, V2C_252_212, V2C_303_212, V2C_410_212, V2C_499_212, V2C_659_212, V2C_720_212, V2C_840_212, V2C_882_212, V2C_945_212, V2C_976_212, V2C_1056_212, V2C_1075_212, V2C_1106_212, V2C_1363_212, V2C_1364_212, V2C_44_213, V2C_71_213, V2C_136_213, V2C_170_213, V2C_236_213, V2C_255_213, V2C_352_213, V2C_407_213, V2C_566_213, V2C_623_213, V2C_651_213, V2C_755_213, V2C_886_213, V2C_930_213, V2C_1003_213, V2C_1015_213, V2C_1093_213, V2C_1138_213, V2C_1364_213, V2C_1365_213, V2C_15_214, V2C_74_214, V2C_113_214, V2C_169_214, V2C_234_214, V2C_288_214, V2C_464_214, V2C_504_214, V2C_540_214, V2C_602_214, V2C_627_214, V2C_673_214, V2C_890_214, V2C_914_214, V2C_998_214, V2C_1028_214, V2C_1103_214, V2C_1119_214, V2C_1365_214, V2C_1366_214, V2C_34_215, V2C_92_215, V2C_127_215, V2C_150_215, V2C_214_215, V2C_280_215, V2C_329_215, V2C_348_215, V2C_475_215, V2C_709_215, V2C_725_215, V2C_779_215, V2C_905_215, V2C_953_215, V2C_996_215, V2C_1048_215, V2C_1097_215, V2C_1145_215, V2C_1366_215, V2C_1367_215, V2C_17_216, V2C_89_216, V2C_129_216, V2C_149_216, V2C_231_216, V2C_262_216, V2C_315_216, V2C_467_216, V2C_564_216, V2C_597_216, V2C_801_216, V2C_829_216, V2C_910_216, V2C_924_216, V2C_1007_216, V2C_1026_216, V2C_1090_216, V2C_1140_216, V2C_1367_216, V2C_1368_216, V2C_41_217, V2C_77_217, V2C_97_217, V2C_158_217, V2C_220_217, V2C_263_217, V2C_363_217, V2C_417_217, V2C_514_217, V2C_750_217, V2C_798_217, V2C_846_217, V2C_887_217, V2C_928_217, V2C_962_217, V2C_1049_217, V2C_1075_217, V2C_1134_217, V2C_1368_217, V2C_1369_217, V2C_2_218, V2C_51_218, V2C_107_218, V2C_155_218, V2C_232_218, V2C_253_218, V2C_304_218, V2C_411_218, V2C_500_218, V2C_660_218, V2C_673_218, V2C_841_218, V2C_883_218, V2C_946_218, V2C_977_218, V2C_1009_218, V2C_1076_218, V2C_1107_218, V2C_1369_218, V2C_1370_218, V2C_45_219, V2C_72_219, V2C_137_219, V2C_171_219, V2C_237_219, V2C_256_219, V2C_353_219, V2C_408_219, V2C_567_219, V2C_624_219, V2C_652_219, V2C_756_219, V2C_887_219, V2C_931_219, V2C_1004_219, V2C_1016_219, V2C_1094_219, V2C_1139_219, V2C_1370_219, V2C_1371_219, V2C_16_220, V2C_75_220, V2C_114_220, V2C_170_220, V2C_235_220, V2C_241_220, V2C_465_220, V2C_505_220, V2C_541_220, V2C_603_220, V2C_628_220, V2C_674_220, V2C_891_220, V2C_915_220, V2C_999_220, V2C_1029_220, V2C_1104_220, V2C_1120_220, V2C_1371_220, V2C_1372_220, V2C_35_221, V2C_93_221, V2C_128_221, V2C_151_221, V2C_215_221, V2C_281_221, V2C_330_221, V2C_349_221, V2C_476_221, V2C_710_221, V2C_726_221, V2C_780_221, V2C_906_221, V2C_954_221, V2C_997_221, V2C_1049_221, V2C_1098_221, V2C_1146_221, V2C_1372_221, V2C_1373_221, V2C_18_222, V2C_90_222, V2C_130_222, V2C_150_222, V2C_232_222, V2C_263_222, V2C_316_222, V2C_468_222, V2C_565_222, V2C_598_222, V2C_802_222, V2C_830_222, V2C_911_222, V2C_925_222, V2C_1008_222, V2C_1027_222, V2C_1091_222, V2C_1141_222, V2C_1373_222, V2C_1374_222, V2C_42_223, V2C_78_223, V2C_98_223, V2C_159_223, V2C_221_223, V2C_264_223, V2C_364_223, V2C_418_223, V2C_515_223, V2C_751_223, V2C_799_223, V2C_847_223, V2C_888_223, V2C_929_223, V2C_963_223, V2C_1050_223, V2C_1076_223, V2C_1135_223, V2C_1374_223, V2C_1375_223, V2C_3_224, V2C_52_224, V2C_108_224, V2C_156_224, V2C_233_224, V2C_254_224, V2C_305_224, V2C_412_224, V2C_501_224, V2C_661_224, V2C_674_224, V2C_842_224, V2C_884_224, V2C_947_224, V2C_978_224, V2C_1010_224, V2C_1077_224, V2C_1108_224, V2C_1375_224, V2C_1376_224, V2C_46_225, V2C_73_225, V2C_138_225, V2C_172_225, V2C_238_225, V2C_257_225, V2C_354_225, V2C_409_225, V2C_568_225, V2C_577_225, V2C_653_225, V2C_757_225, V2C_888_225, V2C_932_225, V2C_1005_225, V2C_1017_225, V2C_1095_225, V2C_1140_225, V2C_1376_225, V2C_1377_225, V2C_17_226, V2C_76_226, V2C_115_226, V2C_171_226, V2C_236_226, V2C_242_226, V2C_466_226, V2C_506_226, V2C_542_226, V2C_604_226, V2C_629_226, V2C_675_226, V2C_892_226, V2C_916_226, V2C_1000_226, V2C_1030_226, V2C_1057_226, V2C_1121_226, V2C_1377_226, V2C_1378_226, V2C_36_227, V2C_94_227, V2C_129_227, V2C_152_227, V2C_216_227, V2C_282_227, V2C_331_227, V2C_350_227, V2C_477_227, V2C_711_227, V2C_727_227, V2C_781_227, V2C_907_227, V2C_955_227, V2C_998_227, V2C_1050_227, V2C_1099_227, V2C_1147_227, V2C_1378_227, V2C_1379_227, V2C_19_228, V2C_91_228, V2C_131_228, V2C_151_228, V2C_233_228, V2C_264_228, V2C_317_228, V2C_469_228, V2C_566_228, V2C_599_228, V2C_803_228, V2C_831_228, V2C_912_228, V2C_926_228, V2C_961_228, V2C_1028_228, V2C_1092_228, V2C_1142_228, V2C_1379_228, V2C_1380_228, V2C_43_229, V2C_79_229, V2C_99_229, V2C_160_229, V2C_222_229, V2C_265_229, V2C_365_229, V2C_419_229, V2C_516_229, V2C_752_229, V2C_800_229, V2C_848_229, V2C_889_229, V2C_930_229, V2C_964_229, V2C_1051_229, V2C_1077_229, V2C_1136_229, V2C_1380_229, V2C_1381_229, V2C_4_230, V2C_53_230, V2C_109_230, V2C_157_230, V2C_234_230, V2C_255_230, V2C_306_230, V2C_413_230, V2C_502_230, V2C_662_230, V2C_675_230, V2C_843_230, V2C_885_230, V2C_948_230, V2C_979_230, V2C_1011_230, V2C_1078_230, V2C_1109_230, V2C_1381_230, V2C_1382_230, V2C_47_231, V2C_74_231, V2C_139_231, V2C_173_231, V2C_239_231, V2C_258_231, V2C_355_231, V2C_410_231, V2C_569_231, V2C_578_231, V2C_654_231, V2C_758_231, V2C_889_231, V2C_933_231, V2C_1006_231, V2C_1018_231, V2C_1096_231, V2C_1141_231, V2C_1382_231, V2C_1383_231, V2C_18_232, V2C_77_232, V2C_116_232, V2C_172_232, V2C_237_232, V2C_243_232, V2C_467_232, V2C_507_232, V2C_543_232, V2C_605_232, V2C_630_232, V2C_676_232, V2C_893_232, V2C_917_232, V2C_1001_232, V2C_1031_232, V2C_1058_232, V2C_1122_232, V2C_1383_232, V2C_1384_232, V2C_37_233, V2C_95_233, V2C_130_233, V2C_153_233, V2C_217_233, V2C_283_233, V2C_332_233, V2C_351_233, V2C_478_233, V2C_712_233, V2C_728_233, V2C_782_233, V2C_908_233, V2C_956_233, V2C_999_233, V2C_1051_233, V2C_1100_233, V2C_1148_233, V2C_1384_233, V2C_1385_233, V2C_20_234, V2C_92_234, V2C_132_234, V2C_152_234, V2C_234_234, V2C_265_234, V2C_318_234, V2C_470_234, V2C_567_234, V2C_600_234, V2C_804_234, V2C_832_234, V2C_865_234, V2C_927_234, V2C_962_234, V2C_1029_234, V2C_1093_234, V2C_1143_234, V2C_1385_234, V2C_1386_234, V2C_44_235, V2C_80_235, V2C_100_235, V2C_161_235, V2C_223_235, V2C_266_235, V2C_366_235, V2C_420_235, V2C_517_235, V2C_753_235, V2C_801_235, V2C_849_235, V2C_890_235, V2C_931_235, V2C_965_235, V2C_1052_235, V2C_1078_235, V2C_1137_235, V2C_1386_235, V2C_1387_235, V2C_5_236, V2C_54_236, V2C_110_236, V2C_158_236, V2C_235_236, V2C_256_236, V2C_307_236, V2C_414_236, V2C_503_236, V2C_663_236, V2C_676_236, V2C_844_236, V2C_886_236, V2C_949_236, V2C_980_236, V2C_1012_236, V2C_1079_236, V2C_1110_236, V2C_1387_236, V2C_1388_236, V2C_48_237, V2C_75_237, V2C_140_237, V2C_174_237, V2C_240_237, V2C_259_237, V2C_356_237, V2C_411_237, V2C_570_237, V2C_579_237, V2C_655_237, V2C_759_237, V2C_890_237, V2C_934_237, V2C_1007_237, V2C_1019_237, V2C_1097_237, V2C_1142_237, V2C_1388_237, V2C_1389_237, V2C_19_238, V2C_78_238, V2C_117_238, V2C_173_238, V2C_238_238, V2C_244_238, V2C_468_238, V2C_508_238, V2C_544_238, V2C_606_238, V2C_631_238, V2C_677_238, V2C_894_238, V2C_918_238, V2C_1002_238, V2C_1032_238, V2C_1059_238, V2C_1123_238, V2C_1389_238, V2C_1390_238, V2C_38_239, V2C_96_239, V2C_131_239, V2C_154_239, V2C_218_239, V2C_284_239, V2C_333_239, V2C_352_239, V2C_479_239, V2C_713_239, V2C_729_239, V2C_783_239, V2C_909_239, V2C_957_239, V2C_1000_239, V2C_1052_239, V2C_1101_239, V2C_1149_239, V2C_1390_239, V2C_1391_239, V2C_21_240, V2C_93_240, V2C_133_240, V2C_153_240, V2C_235_240, V2C_266_240, V2C_319_240, V2C_471_240, V2C_568_240, V2C_601_240, V2C_805_240, V2C_833_240, V2C_866_240, V2C_928_240, V2C_963_240, V2C_1030_240, V2C_1094_240, V2C_1144_240, V2C_1391_240, V2C_1392_240, V2C_45_241, V2C_81_241, V2C_101_241, V2C_162_241, V2C_224_241, V2C_267_241, V2C_367_241, V2C_421_241, V2C_518_241, V2C_754_241, V2C_802_241, V2C_850_241, V2C_891_241, V2C_932_241, V2C_966_241, V2C_1053_241, V2C_1079_241, V2C_1138_241, V2C_1392_241, V2C_1393_241, V2C_6_242, V2C_55_242, V2C_111_242, V2C_159_242, V2C_236_242, V2C_257_242, V2C_308_242, V2C_415_242, V2C_504_242, V2C_664_242, V2C_677_242, V2C_845_242, V2C_887_242, V2C_950_242, V2C_981_242, V2C_1013_242, V2C_1080_242, V2C_1111_242, V2C_1393_242, V2C_1394_242, V2C_1_243, V2C_76_243, V2C_141_243, V2C_175_243, V2C_193_243, V2C_260_243, V2C_357_243, V2C_412_243, V2C_571_243, V2C_580_243, V2C_656_243, V2C_760_243, V2C_891_243, V2C_935_243, V2C_1008_243, V2C_1020_243, V2C_1098_243, V2C_1143_243, V2C_1394_243, V2C_1395_243, V2C_20_244, V2C_79_244, V2C_118_244, V2C_174_244, V2C_239_244, V2C_245_244, V2C_469_244, V2C_509_244, V2C_545_244, V2C_607_244, V2C_632_244, V2C_678_244, V2C_895_244, V2C_919_244, V2C_1003_244, V2C_1033_244, V2C_1060_244, V2C_1124_244, V2C_1395_244, V2C_1396_244, V2C_39_245, V2C_49_245, V2C_132_245, V2C_155_245, V2C_219_245, V2C_285_245, V2C_334_245, V2C_353_245, V2C_480_245, V2C_714_245, V2C_730_245, V2C_784_245, V2C_910_245, V2C_958_245, V2C_1001_245, V2C_1053_245, V2C_1102_245, V2C_1150_245, V2C_1396_245, V2C_1397_245, V2C_22_246, V2C_94_246, V2C_134_246, V2C_154_246, V2C_236_246, V2C_267_246, V2C_320_246, V2C_472_246, V2C_569_246, V2C_602_246, V2C_806_246, V2C_834_246, V2C_867_246, V2C_929_246, V2C_964_246, V2C_1031_246, V2C_1095_246, V2C_1145_246, V2C_1397_246, V2C_1398_246, V2C_46_247, V2C_82_247, V2C_102_247, V2C_163_247, V2C_225_247, V2C_268_247, V2C_368_247, V2C_422_247, V2C_519_247, V2C_755_247, V2C_803_247, V2C_851_247, V2C_892_247, V2C_933_247, V2C_967_247, V2C_1054_247, V2C_1080_247, V2C_1139_247, V2C_1398_247, V2C_1399_247, V2C_7_248, V2C_56_248, V2C_112_248, V2C_160_248, V2C_237_248, V2C_258_248, V2C_309_248, V2C_416_248, V2C_505_248, V2C_665_248, V2C_678_248, V2C_846_248, V2C_888_248, V2C_951_248, V2C_982_248, V2C_1014_248, V2C_1081_248, V2C_1112_248, V2C_1399_248, V2C_1400_248, V2C_2_249, V2C_77_249, V2C_142_249, V2C_176_249, V2C_194_249, V2C_261_249, V2C_358_249, V2C_413_249, V2C_572_249, V2C_581_249, V2C_657_249, V2C_761_249, V2C_892_249, V2C_936_249, V2C_961_249, V2C_1021_249, V2C_1099_249, V2C_1144_249, V2C_1400_249, V2C_1401_249, V2C_21_250, V2C_80_250, V2C_119_250, V2C_175_250, V2C_240_250, V2C_246_250, V2C_470_250, V2C_510_250, V2C_546_250, V2C_608_250, V2C_633_250, V2C_679_250, V2C_896_250, V2C_920_250, V2C_1004_250, V2C_1034_250, V2C_1061_250, V2C_1125_250, V2C_1401_250, V2C_1402_250, V2C_40_251, V2C_50_251, V2C_133_251, V2C_156_251, V2C_220_251, V2C_286_251, V2C_335_251, V2C_354_251, V2C_433_251, V2C_715_251, V2C_731_251, V2C_785_251, V2C_911_251, V2C_959_251, V2C_1002_251, V2C_1054_251, V2C_1103_251, V2C_1151_251, V2C_1402_251, V2C_1403_251, V2C_23_252, V2C_95_252, V2C_135_252, V2C_155_252, V2C_237_252, V2C_268_252, V2C_321_252, V2C_473_252, V2C_570_252, V2C_603_252, V2C_807_252, V2C_835_252, V2C_868_252, V2C_930_252, V2C_965_252, V2C_1032_252, V2C_1096_252, V2C_1146_252, V2C_1403_252, V2C_1404_252, V2C_47_253, V2C_83_253, V2C_103_253, V2C_164_253, V2C_226_253, V2C_269_253, V2C_369_253, V2C_423_253, V2C_520_253, V2C_756_253, V2C_804_253, V2C_852_253, V2C_893_253, V2C_934_253, V2C_968_253, V2C_1055_253, V2C_1081_253, V2C_1140_253, V2C_1404_253, V2C_1405_253, V2C_8_254, V2C_57_254, V2C_113_254, V2C_161_254, V2C_238_254, V2C_259_254, V2C_310_254, V2C_417_254, V2C_506_254, V2C_666_254, V2C_679_254, V2C_847_254, V2C_889_254, V2C_952_254, V2C_983_254, V2C_1015_254, V2C_1082_254, V2C_1113_254, V2C_1405_254, V2C_1406_254, V2C_3_255, V2C_78_255, V2C_143_255, V2C_177_255, V2C_195_255, V2C_262_255, V2C_359_255, V2C_414_255, V2C_573_255, V2C_582_255, V2C_658_255, V2C_762_255, V2C_893_255, V2C_937_255, V2C_962_255, V2C_1022_255, V2C_1100_255, V2C_1145_255, V2C_1406_255, V2C_1407_255, V2C_22_256, V2C_81_256, V2C_120_256, V2C_176_256, V2C_193_256, V2C_247_256, V2C_471_256, V2C_511_256, V2C_547_256, V2C_609_256, V2C_634_256, V2C_680_256, V2C_897_256, V2C_921_256, V2C_1005_256, V2C_1035_256, V2C_1062_256, V2C_1126_256, V2C_1407_256, V2C_1408_256, V2C_41_257, V2C_51_257, V2C_134_257, V2C_157_257, V2C_221_257, V2C_287_257, V2C_336_257, V2C_355_257, V2C_434_257, V2C_716_257, V2C_732_257, V2C_786_257, V2C_912_257, V2C_960_257, V2C_1003_257, V2C_1055_257, V2C_1104_257, V2C_1152_257, V2C_1408_257, V2C_1409_257, V2C_24_258, V2C_96_258, V2C_136_258, V2C_156_258, V2C_238_258, V2C_269_258, V2C_322_258, V2C_474_258, V2C_571_258, V2C_604_258, V2C_808_258, V2C_836_258, V2C_869_258, V2C_931_258, V2C_966_258, V2C_1033_258, V2C_1097_258, V2C_1147_258, V2C_1409_258, V2C_1410_258, V2C_48_259, V2C_84_259, V2C_104_259, V2C_165_259, V2C_227_259, V2C_270_259, V2C_370_259, V2C_424_259, V2C_521_259, V2C_757_259, V2C_805_259, V2C_853_259, V2C_894_259, V2C_935_259, V2C_969_259, V2C_1056_259, V2C_1082_259, V2C_1141_259, V2C_1410_259, V2C_1411_259, V2C_9_260, V2C_58_260, V2C_114_260, V2C_162_260, V2C_239_260, V2C_260_260, V2C_311_260, V2C_418_260, V2C_507_260, V2C_667_260, V2C_680_260, V2C_848_260, V2C_890_260, V2C_953_260, V2C_984_260, V2C_1016_260, V2C_1083_260, V2C_1114_260, V2C_1411_260, V2C_1412_260, V2C_4_261, V2C_79_261, V2C_144_261, V2C_178_261, V2C_196_261, V2C_263_261, V2C_360_261, V2C_415_261, V2C_574_261, V2C_583_261, V2C_659_261, V2C_763_261, V2C_894_261, V2C_938_261, V2C_963_261, V2C_1023_261, V2C_1101_261, V2C_1146_261, V2C_1412_261, V2C_1413_261, V2C_23_262, V2C_82_262, V2C_121_262, V2C_177_262, V2C_194_262, V2C_248_262, V2C_472_262, V2C_512_262, V2C_548_262, V2C_610_262, V2C_635_262, V2C_681_262, V2C_898_262, V2C_922_262, V2C_1006_262, V2C_1036_262, V2C_1063_262, V2C_1127_262, V2C_1413_262, V2C_1414_262, V2C_42_263, V2C_52_263, V2C_135_263, V2C_158_263, V2C_222_263, V2C_288_263, V2C_289_263, V2C_356_263, V2C_435_263, V2C_717_263, V2C_733_263, V2C_787_263, V2C_865_263, V2C_913_263, V2C_1004_263, V2C_1056_263, V2C_1057_263, V2C_1105_263, V2C_1414_263, V2C_1415_263, V2C_25_264, V2C_49_264, V2C_137_264, V2C_157_264, V2C_239_264, V2C_270_264, V2C_323_264, V2C_475_264, V2C_572_264, V2C_605_264, V2C_809_264, V2C_837_264, V2C_870_264, V2C_932_264, V2C_967_264, V2C_1034_264, V2C_1098_264, V2C_1148_264, V2C_1415_264, V2C_1416_264, V2C_1_265, V2C_85_265, V2C_105_265, V2C_166_265, V2C_228_265, V2C_271_265, V2C_371_265, V2C_425_265, V2C_522_265, V2C_758_265, V2C_806_265, V2C_854_265, V2C_895_265, V2C_936_265, V2C_970_265, V2C_1009_265, V2C_1083_265, V2C_1142_265, V2C_1416_265, V2C_1417_265, V2C_10_266, V2C_59_266, V2C_115_266, V2C_163_266, V2C_240_266, V2C_261_266, V2C_312_266, V2C_419_266, V2C_508_266, V2C_668_266, V2C_681_266, V2C_849_266, V2C_891_266, V2C_954_266, V2C_985_266, V2C_1017_266, V2C_1084_266, V2C_1115_266, V2C_1417_266, V2C_1418_266, V2C_5_267, V2C_80_267, V2C_97_267, V2C_179_267, V2C_197_267, V2C_264_267, V2C_361_267, V2C_416_267, V2C_575_267, V2C_584_267, V2C_660_267, V2C_764_267, V2C_895_267, V2C_939_267, V2C_964_267, V2C_1024_267, V2C_1102_267, V2C_1147_267, V2C_1418_267, V2C_1419_267, V2C_24_268, V2C_83_268, V2C_122_268, V2C_178_268, V2C_195_268, V2C_249_268, V2C_473_268, V2C_513_268, V2C_549_268, V2C_611_268, V2C_636_268, V2C_682_268, V2C_899_268, V2C_923_268, V2C_1007_268, V2C_1037_268, V2C_1064_268, V2C_1128_268, V2C_1419_268, V2C_1420_268, V2C_43_269, V2C_53_269, V2C_136_269, V2C_159_269, V2C_223_269, V2C_241_269, V2C_290_269, V2C_357_269, V2C_436_269, V2C_718_269, V2C_734_269, V2C_788_269, V2C_866_269, V2C_914_269, V2C_1005_269, V2C_1009_269, V2C_1058_269, V2C_1106_269, V2C_1420_269, V2C_1421_269, V2C_26_270, V2C_50_270, V2C_138_270, V2C_158_270, V2C_240_270, V2C_271_270, V2C_324_270, V2C_476_270, V2C_573_270, V2C_606_270, V2C_810_270, V2C_838_270, V2C_871_270, V2C_933_270, V2C_968_270, V2C_1035_270, V2C_1099_270, V2C_1149_270, V2C_1421_270, V2C_1422_270, V2C_2_271, V2C_86_271, V2C_106_271, V2C_167_271, V2C_229_271, V2C_272_271, V2C_372_271, V2C_426_271, V2C_523_271, V2C_759_271, V2C_807_271, V2C_855_271, V2C_896_271, V2C_937_271, V2C_971_271, V2C_1010_271, V2C_1084_271, V2C_1143_271, V2C_1422_271, V2C_1423_271, V2C_11_272, V2C_60_272, V2C_116_272, V2C_164_272, V2C_193_272, V2C_262_272, V2C_313_272, V2C_420_272, V2C_509_272, V2C_669_272, V2C_682_272, V2C_850_272, V2C_892_272, V2C_955_272, V2C_986_272, V2C_1018_272, V2C_1085_272, V2C_1116_272, V2C_1423_272, V2C_1424_272, V2C_6_273, V2C_81_273, V2C_98_273, V2C_180_273, V2C_198_273, V2C_265_273, V2C_362_273, V2C_417_273, V2C_576_273, V2C_585_273, V2C_661_273, V2C_765_273, V2C_896_273, V2C_940_273, V2C_965_273, V2C_1025_273, V2C_1103_273, V2C_1148_273, V2C_1424_273, V2C_1425_273, V2C_25_274, V2C_84_274, V2C_123_274, V2C_179_274, V2C_196_274, V2C_250_274, V2C_474_274, V2C_514_274, V2C_550_274, V2C_612_274, V2C_637_274, V2C_683_274, V2C_900_274, V2C_924_274, V2C_1008_274, V2C_1038_274, V2C_1065_274, V2C_1129_274, V2C_1425_274, V2C_1426_274, V2C_44_275, V2C_54_275, V2C_137_275, V2C_160_275, V2C_224_275, V2C_242_275, V2C_291_275, V2C_358_275, V2C_437_275, V2C_719_275, V2C_735_275, V2C_789_275, V2C_867_275, V2C_915_275, V2C_1006_275, V2C_1010_275, V2C_1059_275, V2C_1107_275, V2C_1426_275, V2C_1427_275, V2C_27_276, V2C_51_276, V2C_139_276, V2C_159_276, V2C_193_276, V2C_272_276, V2C_325_276, V2C_477_276, V2C_574_276, V2C_607_276, V2C_811_276, V2C_839_276, V2C_872_276, V2C_934_276, V2C_969_276, V2C_1036_276, V2C_1100_276, V2C_1150_276, V2C_1427_276, V2C_1428_276, V2C_3_277, V2C_87_277, V2C_107_277, V2C_168_277, V2C_230_277, V2C_273_277, V2C_373_277, V2C_427_277, V2C_524_277, V2C_760_277, V2C_808_277, V2C_856_277, V2C_897_277, V2C_938_277, V2C_972_277, V2C_1011_277, V2C_1085_277, V2C_1144_277, V2C_1428_277, V2C_1429_277, V2C_12_278, V2C_61_278, V2C_117_278, V2C_165_278, V2C_194_278, V2C_263_278, V2C_314_278, V2C_421_278, V2C_510_278, V2C_670_278, V2C_683_278, V2C_851_278, V2C_893_278, V2C_956_278, V2C_987_278, V2C_1019_278, V2C_1086_278, V2C_1117_278, V2C_1429_278, V2C_1430_278, V2C_7_279, V2C_82_279, V2C_99_279, V2C_181_279, V2C_199_279, V2C_266_279, V2C_363_279, V2C_418_279, V2C_529_279, V2C_586_279, V2C_662_279, V2C_766_279, V2C_897_279, V2C_941_279, V2C_966_279, V2C_1026_279, V2C_1104_279, V2C_1149_279, V2C_1430_279, V2C_1431_279, V2C_26_280, V2C_85_280, V2C_124_280, V2C_180_280, V2C_197_280, V2C_251_280, V2C_475_280, V2C_515_280, V2C_551_280, V2C_613_280, V2C_638_280, V2C_684_280, V2C_901_280, V2C_925_280, V2C_961_280, V2C_1039_280, V2C_1066_280, V2C_1130_280, V2C_1431_280, V2C_1432_280, V2C_45_281, V2C_55_281, V2C_138_281, V2C_161_281, V2C_225_281, V2C_243_281, V2C_292_281, V2C_359_281, V2C_438_281, V2C_720_281, V2C_736_281, V2C_790_281, V2C_868_281, V2C_916_281, V2C_1007_281, V2C_1011_281, V2C_1060_281, V2C_1108_281, V2C_1432_281, V2C_1433_281, V2C_28_282, V2C_52_282, V2C_140_282, V2C_160_282, V2C_194_282, V2C_273_282, V2C_326_282, V2C_478_282, V2C_575_282, V2C_608_282, V2C_812_282, V2C_840_282, V2C_873_282, V2C_935_282, V2C_970_282, V2C_1037_282, V2C_1101_282, V2C_1151_282, V2C_1433_282, V2C_1434_282, V2C_4_283, V2C_88_283, V2C_108_283, V2C_169_283, V2C_231_283, V2C_274_283, V2C_374_283, V2C_428_283, V2C_525_283, V2C_761_283, V2C_809_283, V2C_857_283, V2C_898_283, V2C_939_283, V2C_973_283, V2C_1012_283, V2C_1086_283, V2C_1145_283, V2C_1434_283, V2C_1435_283, V2C_13_284, V2C_62_284, V2C_118_284, V2C_166_284, V2C_195_284, V2C_264_284, V2C_315_284, V2C_422_284, V2C_511_284, V2C_671_284, V2C_684_284, V2C_852_284, V2C_894_284, V2C_957_284, V2C_988_284, V2C_1020_284, V2C_1087_284, V2C_1118_284, V2C_1435_284, V2C_1436_284, V2C_8_285, V2C_83_285, V2C_100_285, V2C_182_285, V2C_200_285, V2C_267_285, V2C_364_285, V2C_419_285, V2C_530_285, V2C_587_285, V2C_663_285, V2C_767_285, V2C_898_285, V2C_942_285, V2C_967_285, V2C_1027_285, V2C_1057_285, V2C_1150_285, V2C_1436_285, V2C_1437_285, V2C_27_286, V2C_86_286, V2C_125_286, V2C_181_286, V2C_198_286, V2C_252_286, V2C_476_286, V2C_516_286, V2C_552_286, V2C_614_286, V2C_639_286, V2C_685_286, V2C_902_286, V2C_926_286, V2C_962_286, V2C_1040_286, V2C_1067_286, V2C_1131_286, V2C_1437_286, V2C_1438_286, V2C_46_287, V2C_56_287, V2C_139_287, V2C_162_287, V2C_226_287, V2C_244_287, V2C_293_287, V2C_360_287, V2C_439_287, V2C_673_287, V2C_737_287, V2C_791_287, V2C_869_287, V2C_917_287, V2C_1008_287, V2C_1012_287, V2C_1061_287, V2C_1109_287, V2C_1438_287, V2C_1439_287, V2C_29_288, V2C_53_288, V2C_141_288, V2C_161_288, V2C_195_288, V2C_274_288, V2C_327_288, V2C_479_288, V2C_576_288, V2C_609_288, V2C_813_288, V2C_841_288, V2C_874_288, V2C_936_288, V2C_971_288, V2C_1038_288, V2C_1102_288, V2C_1152_288, V2C_1439_288, V2C_1440_288, V2C_0_0;
wire [quan_width - 1:0] V_1, V_2, V_3, V_4, V_5, V_6, V_7, V_8, V_9, V_10, V_11, V_12, V_13, V_14, V_15, V_16, V_17, V_18, V_19, V_20, V_21, V_22, V_23, V_24, V_25, V_26, V_27, V_28, V_29, V_30, V_31, V_32, V_33, V_34, V_35, V_36, V_37, V_38, V_39, V_40, V_41, V_42, V_43, V_44, V_45, V_46, V_47, V_48, V_49, V_50, V_51, V_52, V_53, V_54, V_55, V_56, V_57, V_58, V_59, V_60, V_61, V_62, V_63, V_64, V_65, V_66, V_67, V_68, V_69, V_70, V_71, V_72, V_73, V_74, V_75, V_76, V_77, V_78, V_79, V_80, V_81, V_82, V_83, V_84, V_85, V_86, V_87, V_88, V_89, V_90, V_91, V_92, V_93, V_94, V_95, V_96, V_97, V_98, V_99, V_100, V_101, V_102, V_103, V_104, V_105, V_106, V_107, V_108, V_109, V_110, V_111, V_112, V_113, V_114, V_115, V_116, V_117, V_118, V_119, V_120, V_121, V_122, V_123, V_124, V_125, V_126, V_127, V_128, V_129, V_130, V_131, V_132, V_133, V_134, V_135, V_136, V_137, V_138, V_139, V_140, V_141, V_142, V_143, V_144, V_145, V_146, V_147, V_148, V_149, V_150, V_151, V_152, V_153, V_154, V_155, V_156, V_157, V_158, V_159, V_160, V_161, V_162, V_163, V_164, V_165, V_166, V_167, V_168, V_169, V_170, V_171, V_172, V_173, V_174, V_175, V_176, V_177, V_178, V_179, V_180, V_181, V_182, V_183, V_184, V_185, V_186, V_187, V_188, V_189, V_190, V_191, V_192, V_193, V_194, V_195, V_196, V_197, V_198, V_199, V_200, V_201, V_202, V_203, V_204, V_205, V_206, V_207, V_208, V_209, V_210, V_211, V_212, V_213, V_214, V_215, V_216, V_217, V_218, V_219, V_220, V_221, V_222, V_223, V_224, V_225, V_226, V_227, V_228, V_229, V_230, V_231, V_232, V_233, V_234, V_235, V_236, V_237, V_238, V_239, V_240, V_241, V_242, V_243, V_244, V_245, V_246, V_247, V_248, V_249, V_250, V_251, V_252, V_253, V_254, V_255, V_256, V_257, V_258, V_259, V_260, V_261, V_262, V_263, V_264, V_265, V_266, V_267, V_268, V_269, V_270, V_271, V_272, V_273, V_274, V_275, V_276, V_277, V_278, V_279, V_280, V_281, V_282, V_283, V_284, V_285, V_286, V_287, V_288, V_289, V_290, V_291, V_292, V_293, V_294, V_295, V_296, V_297, V_298, V_299, V_300, V_301, V_302, V_303, V_304, V_305, V_306, V_307, V_308, V_309, V_310, V_311, V_312, V_313, V_314, V_315, V_316, V_317, V_318, V_319, V_320, V_321, V_322, V_323, V_324, V_325, V_326, V_327, V_328, V_329, V_330, V_331, V_332, V_333, V_334, V_335, V_336, V_337, V_338, V_339, V_340, V_341, V_342, V_343, V_344, V_345, V_346, V_347, V_348, V_349, V_350, V_351, V_352, V_353, V_354, V_355, V_356, V_357, V_358, V_359, V_360, V_361, V_362, V_363, V_364, V_365, V_366, V_367, V_368, V_369, V_370, V_371, V_372, V_373, V_374, V_375, V_376, V_377, V_378, V_379, V_380, V_381, V_382, V_383, V_384, V_385, V_386, V_387, V_388, V_389, V_390, V_391, V_392, V_393, V_394, V_395, V_396, V_397, V_398, V_399, V_400, V_401, V_402, V_403, V_404, V_405, V_406, V_407, V_408, V_409, V_410, V_411, V_412, V_413, V_414, V_415, V_416, V_417, V_418, V_419, V_420, V_421, V_422, V_423, V_424, V_425, V_426, V_427, V_428, V_429, V_430, V_431, V_432, V_433, V_434, V_435, V_436, V_437, V_438, V_439, V_440, V_441, V_442, V_443, V_444, V_445, V_446, V_447, V_448, V_449, V_450, V_451, V_452, V_453, V_454, V_455, V_456, V_457, V_458, V_459, V_460, V_461, V_462, V_463, V_464, V_465, V_466, V_467, V_468, V_469, V_470, V_471, V_472, V_473, V_474, V_475, V_476, V_477, V_478, V_479, V_480, V_481, V_482, V_483, V_484, V_485, V_486, V_487, V_488, V_489, V_490, V_491, V_492, V_493, V_494, V_495, V_496, V_497, V_498, V_499, V_500, V_501, V_502, V_503, V_504, V_505, V_506, V_507, V_508, V_509, V_510, V_511, V_512, V_513, V_514, V_515, V_516, V_517, V_518, V_519, V_520, V_521, V_522, V_523, V_524, V_525, V_526, V_527, V_528, V_529, V_530, V_531, V_532, V_533, V_534, V_535, V_536, V_537, V_538, V_539, V_540, V_541, V_542, V_543, V_544, V_545, V_546, V_547, V_548, V_549, V_550, V_551, V_552, V_553, V_554, V_555, V_556, V_557, V_558, V_559, V_560, V_561, V_562, V_563, V_564, V_565, V_566, V_567, V_568, V_569, V_570, V_571, V_572, V_573, V_574, V_575, V_576, V_577, V_578, V_579, V_580, V_581, V_582, V_583, V_584, V_585, V_586, V_587, V_588, V_589, V_590, V_591, V_592, V_593, V_594, V_595, V_596, V_597, V_598, V_599, V_600, V_601, V_602, V_603, V_604, V_605, V_606, V_607, V_608, V_609, V_610, V_611, V_612, V_613, V_614, V_615, V_616, V_617, V_618, V_619, V_620, V_621, V_622, V_623, V_624, V_625, V_626, V_627, V_628, V_629, V_630, V_631, V_632, V_633, V_634, V_635, V_636, V_637, V_638, V_639, V_640, V_641, V_642, V_643, V_644, V_645, V_646, V_647, V_648, V_649, V_650, V_651, V_652, V_653, V_654, V_655, V_656, V_657, V_658, V_659, V_660, V_661, V_662, V_663, V_664, V_665, V_666, V_667, V_668, V_669, V_670, V_671, V_672, V_673, V_674, V_675, V_676, V_677, V_678, V_679, V_680, V_681, V_682, V_683, V_684, V_685, V_686, V_687, V_688, V_689, V_690, V_691, V_692, V_693, V_694, V_695, V_696, V_697, V_698, V_699, V_700, V_701, V_702, V_703, V_704, V_705, V_706, V_707, V_708, V_709, V_710, V_711, V_712, V_713, V_714, V_715, V_716, V_717, V_718, V_719, V_720, V_721, V_722, V_723, V_724, V_725, V_726, V_727, V_728, V_729, V_730, V_731, V_732, V_733, V_734, V_735, V_736, V_737, V_738, V_739, V_740, V_741, V_742, V_743, V_744, V_745, V_746, V_747, V_748, V_749, V_750, V_751, V_752, V_753, V_754, V_755, V_756, V_757, V_758, V_759, V_760, V_761, V_762, V_763, V_764, V_765, V_766, V_767, V_768, V_769, V_770, V_771, V_772, V_773, V_774, V_775, V_776, V_777, V_778, V_779, V_780, V_781, V_782, V_783, V_784, V_785, V_786, V_787, V_788, V_789, V_790, V_791, V_792, V_793, V_794, V_795, V_796, V_797, V_798, V_799, V_800, V_801, V_802, V_803, V_804, V_805, V_806, V_807, V_808, V_809, V_810, V_811, V_812, V_813, V_814, V_815, V_816, V_817, V_818, V_819, V_820, V_821, V_822, V_823, V_824, V_825, V_826, V_827, V_828, V_829, V_830, V_831, V_832, V_833, V_834, V_835, V_836, V_837, V_838, V_839, V_840, V_841, V_842, V_843, V_844, V_845, V_846, V_847, V_848, V_849, V_850, V_851, V_852, V_853, V_854, V_855, V_856, V_857, V_858, V_859, V_860, V_861, V_862, V_863, V_864, V_865, V_866, V_867, V_868, V_869, V_870, V_871, V_872, V_873, V_874, V_875, V_876, V_877, V_878, V_879, V_880, V_881, V_882, V_883, V_884, V_885, V_886, V_887, V_888, V_889, V_890, V_891, V_892, V_893, V_894, V_895, V_896, V_897, V_898, V_899, V_900, V_901, V_902, V_903, V_904, V_905, V_906, V_907, V_908, V_909, V_910, V_911, V_912, V_913, V_914, V_915, V_916, V_917, V_918, V_919, V_920, V_921, V_922, V_923, V_924, V_925, V_926, V_927, V_928, V_929, V_930, V_931, V_932, V_933, V_934, V_935, V_936, V_937, V_938, V_939, V_940, V_941, V_942, V_943, V_944, V_945, V_946, V_947, V_948, V_949, V_950, V_951, V_952, V_953, V_954, V_955, V_956, V_957, V_958, V_959, V_960, V_961, V_962, V_963, V_964, V_965, V_966, V_967, V_968, V_969, V_970, V_971, V_972, V_973, V_974, V_975, V_976, V_977, V_978, V_979, V_980, V_981, V_982, V_983, V_984, V_985, V_986, V_987, V_988, V_989, V_990, V_991, V_992, V_993, V_994, V_995, V_996, V_997, V_998, V_999, V_1000, V_1001, V_1002, V_1003, V_1004, V_1005, V_1006, V_1007, V_1008, V_1009, V_1010, V_1011, V_1012, V_1013, V_1014, V_1015, V_1016, V_1017, V_1018, V_1019, V_1020, V_1021, V_1022, V_1023, V_1024, V_1025, V_1026, V_1027, V_1028, V_1029, V_1030, V_1031, V_1032, V_1033, V_1034, V_1035, V_1036, V_1037, V_1038, V_1039, V_1040, V_1041, V_1042, V_1043, V_1044, V_1045, V_1046, V_1047, V_1048, V_1049, V_1050, V_1051, V_1052, V_1053, V_1054, V_1055, V_1056, V_1057, V_1058, V_1059, V_1060, V_1061, V_1062, V_1063, V_1064, V_1065, V_1066, V_1067, V_1068, V_1069, V_1070, V_1071, V_1072, V_1073, V_1074, V_1075, V_1076, V_1077, V_1078, V_1079, V_1080, V_1081, V_1082, V_1083, V_1084, V_1085, V_1086, V_1087, V_1088, V_1089, V_1090, V_1091, V_1092, V_1093, V_1094, V_1095, V_1096, V_1097, V_1098, V_1099, V_1100, V_1101, V_1102, V_1103, V_1104, V_1105, V_1106, V_1107, V_1108, V_1109, V_1110, V_1111, V_1112, V_1113, V_1114, V_1115, V_1116, V_1117, V_1118, V_1119, V_1120, V_1121, V_1122, V_1123, V_1124, V_1125, V_1126, V_1127, V_1128, V_1129, V_1130, V_1131, V_1132, V_1133, V_1134, V_1135, V_1136, V_1137, V_1138, V_1139, V_1140, V_1141, V_1142, V_1143, V_1144, V_1145, V_1146, V_1147, V_1148, V_1149, V_1150, V_1151, V_1152, V_1153, V_1154, V_1155, V_1156, V_1157, V_1158, V_1159, V_1160, V_1161, V_1162, V_1163, V_1164, V_1165, V_1166, V_1167, V_1168, V_1169, V_1170, V_1171, V_1172, V_1173, V_1174, V_1175, V_1176, V_1177, V_1178, V_1179, V_1180, V_1181, V_1182, V_1183, V_1184, V_1185, V_1186, V_1187, V_1188, V_1189, V_1190, V_1191, V_1192, V_1193, V_1194, V_1195, V_1196, V_1197, V_1198, V_1199, V_1200, V_1201, V_1202, V_1203, V_1204, V_1205, V_1206, V_1207, V_1208, V_1209, V_1210, V_1211, V_1212, V_1213, V_1214, V_1215, V_1216, V_1217, V_1218, V_1219, V_1220, V_1221, V_1222, V_1223, V_1224, V_1225, V_1226, V_1227, V_1228, V_1229, V_1230, V_1231, V_1232, V_1233, V_1234, V_1235, V_1236, V_1237, V_1238, V_1239, V_1240, V_1241, V_1242, V_1243, V_1244, V_1245, V_1246, V_1247, V_1248, V_1249, V_1250, V_1251, V_1252, V_1253, V_1254, V_1255, V_1256, V_1257, V_1258, V_1259, V_1260, V_1261, V_1262, V_1263, V_1264, V_1265, V_1266, V_1267, V_1268, V_1269, V_1270, V_1271, V_1272, V_1273, V_1274, V_1275, V_1276, V_1277, V_1278, V_1279, V_1280, V_1281, V_1282, V_1283, V_1284, V_1285, V_1286, V_1287, V_1288, V_1289, V_1290, V_1291, V_1292, V_1293, V_1294, V_1295, V_1296, V_1297, V_1298, V_1299, V_1300, V_1301, V_1302, V_1303, V_1304, V_1305, V_1306, V_1307, V_1308, V_1309, V_1310, V_1311, V_1312, V_1313, V_1314, V_1315, V_1316, V_1317, V_1318, V_1319, V_1320, V_1321, V_1322, V_1323, V_1324, V_1325, V_1326, V_1327, V_1328, V_1329, V_1330, V_1331, V_1332, V_1333, V_1334, V_1335, V_1336, V_1337, V_1338, V_1339, V_1340, V_1341, V_1342, V_1343, V_1344, V_1345, V_1346, V_1347, V_1348, V_1349, V_1350, V_1351, V_1352, V_1353, V_1354, V_1355, V_1356, V_1357, V_1358, V_1359, V_1360, V_1361, V_1362, V_1363, V_1364, V_1365, V_1366, V_1367, V_1368, V_1369, V_1370, V_1371, V_1372, V_1373, V_1374, V_1375, V_1376, V_1377, V_1378, V_1379, V_1380, V_1381, V_1382, V_1383, V_1384, V_1385, V_1386, V_1387, V_1388, V_1389, V_1390, V_1391, V_1392, V_1393, V_1394, V_1395, V_1396, V_1397, V_1398, V_1399, V_1400, V_1401, V_1402, V_1403, V_1404, V_1405, V_1406, V_1407, V_1408, V_1409, V_1410, V_1411, V_1412, V_1413, V_1414, V_1415, V_1416, V_1417, V_1418, V_1419, V_1420, V_1421, V_1422, V_1423, V_1424, V_1425, V_1426, V_1427, V_1428, V_1429, V_1430, V_1431, V_1432, V_1433, V_1434, V_1435, V_1436, V_1437, V_1438, V_1439, V_1440;

always @ (posedge clk) begin
	case ({in_valid, in_index})
		{1'b1, 16'd0}: begin L_1 <= data_in[quan_width-1:0]; L_2 <= data_in[quan_width*2-1:quan_width]; L_3 <= data_in[quan_width*3-1:quan_width*2]; L_4 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd4}: begin L_5 <= data_in[quan_width-1:0]; L_6 <= data_in[quan_width*2-1:quan_width]; L_7 <= data_in[quan_width*3-1:quan_width*2]; L_8 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd8}: begin L_9 <= data_in[quan_width-1:0]; L_10 <= data_in[quan_width*2-1:quan_width]; L_11 <= data_in[quan_width*3-1:quan_width*2]; L_12 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd12}: begin L_13 <= data_in[quan_width-1:0]; L_14 <= data_in[quan_width*2-1:quan_width]; L_15 <= data_in[quan_width*3-1:quan_width*2]; L_16 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd16}: begin L_17 <= data_in[quan_width-1:0]; L_18 <= data_in[quan_width*2-1:quan_width]; L_19 <= data_in[quan_width*3-1:quan_width*2]; L_20 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd20}: begin L_21 <= data_in[quan_width-1:0]; L_22 <= data_in[quan_width*2-1:quan_width]; L_23 <= data_in[quan_width*3-1:quan_width*2]; L_24 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd24}: begin L_25 <= data_in[quan_width-1:0]; L_26 <= data_in[quan_width*2-1:quan_width]; L_27 <= data_in[quan_width*3-1:quan_width*2]; L_28 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd28}: begin L_29 <= data_in[quan_width-1:0]; L_30 <= data_in[quan_width*2-1:quan_width]; L_31 <= data_in[quan_width*3-1:quan_width*2]; L_32 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd32}: begin L_33 <= data_in[quan_width-1:0]; L_34 <= data_in[quan_width*2-1:quan_width]; L_35 <= data_in[quan_width*3-1:quan_width*2]; L_36 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd36}: begin L_37 <= data_in[quan_width-1:0]; L_38 <= data_in[quan_width*2-1:quan_width]; L_39 <= data_in[quan_width*3-1:quan_width*2]; L_40 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd40}: begin L_41 <= data_in[quan_width-1:0]; L_42 <= data_in[quan_width*2-1:quan_width]; L_43 <= data_in[quan_width*3-1:quan_width*2]; L_44 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd44}: begin L_45 <= data_in[quan_width-1:0]; L_46 <= data_in[quan_width*2-1:quan_width]; L_47 <= data_in[quan_width*3-1:quan_width*2]; L_48 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd48}: begin L_49 <= data_in[quan_width-1:0]; L_50 <= data_in[quan_width*2-1:quan_width]; L_51 <= data_in[quan_width*3-1:quan_width*2]; L_52 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd52}: begin L_53 <= data_in[quan_width-1:0]; L_54 <= data_in[quan_width*2-1:quan_width]; L_55 <= data_in[quan_width*3-1:quan_width*2]; L_56 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd56}: begin L_57 <= data_in[quan_width-1:0]; L_58 <= data_in[quan_width*2-1:quan_width]; L_59 <= data_in[quan_width*3-1:quan_width*2]; L_60 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd60}: begin L_61 <= data_in[quan_width-1:0]; L_62 <= data_in[quan_width*2-1:quan_width]; L_63 <= data_in[quan_width*3-1:quan_width*2]; L_64 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd64}: begin L_65 <= data_in[quan_width-1:0]; L_66 <= data_in[quan_width*2-1:quan_width]; L_67 <= data_in[quan_width*3-1:quan_width*2]; L_68 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd68}: begin L_69 <= data_in[quan_width-1:0]; L_70 <= data_in[quan_width*2-1:quan_width]; L_71 <= data_in[quan_width*3-1:quan_width*2]; L_72 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd72}: begin L_73 <= data_in[quan_width-1:0]; L_74 <= data_in[quan_width*2-1:quan_width]; L_75 <= data_in[quan_width*3-1:quan_width*2]; L_76 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd76}: begin L_77 <= data_in[quan_width-1:0]; L_78 <= data_in[quan_width*2-1:quan_width]; L_79 <= data_in[quan_width*3-1:quan_width*2]; L_80 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd80}: begin L_81 <= data_in[quan_width-1:0]; L_82 <= data_in[quan_width*2-1:quan_width]; L_83 <= data_in[quan_width*3-1:quan_width*2]; L_84 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd84}: begin L_85 <= data_in[quan_width-1:0]; L_86 <= data_in[quan_width*2-1:quan_width]; L_87 <= data_in[quan_width*3-1:quan_width*2]; L_88 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd88}: begin L_89 <= data_in[quan_width-1:0]; L_90 <= data_in[quan_width*2-1:quan_width]; L_91 <= data_in[quan_width*3-1:quan_width*2]; L_92 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd92}: begin L_93 <= data_in[quan_width-1:0]; L_94 <= data_in[quan_width*2-1:quan_width]; L_95 <= data_in[quan_width*3-1:quan_width*2]; L_96 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd96}: begin L_97 <= data_in[quan_width-1:0]; L_98 <= data_in[quan_width*2-1:quan_width]; L_99 <= data_in[quan_width*3-1:quan_width*2]; L_100 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd100}: begin L_101 <= data_in[quan_width-1:0]; L_102 <= data_in[quan_width*2-1:quan_width]; L_103 <= data_in[quan_width*3-1:quan_width*2]; L_104 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd104}: begin L_105 <= data_in[quan_width-1:0]; L_106 <= data_in[quan_width*2-1:quan_width]; L_107 <= data_in[quan_width*3-1:quan_width*2]; L_108 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd108}: begin L_109 <= data_in[quan_width-1:0]; L_110 <= data_in[quan_width*2-1:quan_width]; L_111 <= data_in[quan_width*3-1:quan_width*2]; L_112 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd112}: begin L_113 <= data_in[quan_width-1:0]; L_114 <= data_in[quan_width*2-1:quan_width]; L_115 <= data_in[quan_width*3-1:quan_width*2]; L_116 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd116}: begin L_117 <= data_in[quan_width-1:0]; L_118 <= data_in[quan_width*2-1:quan_width]; L_119 <= data_in[quan_width*3-1:quan_width*2]; L_120 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd120}: begin L_121 <= data_in[quan_width-1:0]; L_122 <= data_in[quan_width*2-1:quan_width]; L_123 <= data_in[quan_width*3-1:quan_width*2]; L_124 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd124}: begin L_125 <= data_in[quan_width-1:0]; L_126 <= data_in[quan_width*2-1:quan_width]; L_127 <= data_in[quan_width*3-1:quan_width*2]; L_128 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd128}: begin L_129 <= data_in[quan_width-1:0]; L_130 <= data_in[quan_width*2-1:quan_width]; L_131 <= data_in[quan_width*3-1:quan_width*2]; L_132 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd132}: begin L_133 <= data_in[quan_width-1:0]; L_134 <= data_in[quan_width*2-1:quan_width]; L_135 <= data_in[quan_width*3-1:quan_width*2]; L_136 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd136}: begin L_137 <= data_in[quan_width-1:0]; L_138 <= data_in[quan_width*2-1:quan_width]; L_139 <= data_in[quan_width*3-1:quan_width*2]; L_140 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd140}: begin L_141 <= data_in[quan_width-1:0]; L_142 <= data_in[quan_width*2-1:quan_width]; L_143 <= data_in[quan_width*3-1:quan_width*2]; L_144 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd144}: begin L_145 <= data_in[quan_width-1:0]; L_146 <= data_in[quan_width*2-1:quan_width]; L_147 <= data_in[quan_width*3-1:quan_width*2]; L_148 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd148}: begin L_149 <= data_in[quan_width-1:0]; L_150 <= data_in[quan_width*2-1:quan_width]; L_151 <= data_in[quan_width*3-1:quan_width*2]; L_152 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd152}: begin L_153 <= data_in[quan_width-1:0]; L_154 <= data_in[quan_width*2-1:quan_width]; L_155 <= data_in[quan_width*3-1:quan_width*2]; L_156 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd156}: begin L_157 <= data_in[quan_width-1:0]; L_158 <= data_in[quan_width*2-1:quan_width]; L_159 <= data_in[quan_width*3-1:quan_width*2]; L_160 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd160}: begin L_161 <= data_in[quan_width-1:0]; L_162 <= data_in[quan_width*2-1:quan_width]; L_163 <= data_in[quan_width*3-1:quan_width*2]; L_164 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd164}: begin L_165 <= data_in[quan_width-1:0]; L_166 <= data_in[quan_width*2-1:quan_width]; L_167 <= data_in[quan_width*3-1:quan_width*2]; L_168 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd168}: begin L_169 <= data_in[quan_width-1:0]; L_170 <= data_in[quan_width*2-1:quan_width]; L_171 <= data_in[quan_width*3-1:quan_width*2]; L_172 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd172}: begin L_173 <= data_in[quan_width-1:0]; L_174 <= data_in[quan_width*2-1:quan_width]; L_175 <= data_in[quan_width*3-1:quan_width*2]; L_176 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd176}: begin L_177 <= data_in[quan_width-1:0]; L_178 <= data_in[quan_width*2-1:quan_width]; L_179 <= data_in[quan_width*3-1:quan_width*2]; L_180 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd180}: begin L_181 <= data_in[quan_width-1:0]; L_182 <= data_in[quan_width*2-1:quan_width]; L_183 <= data_in[quan_width*3-1:quan_width*2]; L_184 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd184}: begin L_185 <= data_in[quan_width-1:0]; L_186 <= data_in[quan_width*2-1:quan_width]; L_187 <= data_in[quan_width*3-1:quan_width*2]; L_188 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd188}: begin L_189 <= data_in[quan_width-1:0]; L_190 <= data_in[quan_width*2-1:quan_width]; L_191 <= data_in[quan_width*3-1:quan_width*2]; L_192 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd192}: begin L_193 <= data_in[quan_width-1:0]; L_194 <= data_in[quan_width*2-1:quan_width]; L_195 <= data_in[quan_width*3-1:quan_width*2]; L_196 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd196}: begin L_197 <= data_in[quan_width-1:0]; L_198 <= data_in[quan_width*2-1:quan_width]; L_199 <= data_in[quan_width*3-1:quan_width*2]; L_200 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd200}: begin L_201 <= data_in[quan_width-1:0]; L_202 <= data_in[quan_width*2-1:quan_width]; L_203 <= data_in[quan_width*3-1:quan_width*2]; L_204 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd204}: begin L_205 <= data_in[quan_width-1:0]; L_206 <= data_in[quan_width*2-1:quan_width]; L_207 <= data_in[quan_width*3-1:quan_width*2]; L_208 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd208}: begin L_209 <= data_in[quan_width-1:0]; L_210 <= data_in[quan_width*2-1:quan_width]; L_211 <= data_in[quan_width*3-1:quan_width*2]; L_212 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd212}: begin L_213 <= data_in[quan_width-1:0]; L_214 <= data_in[quan_width*2-1:quan_width]; L_215 <= data_in[quan_width*3-1:quan_width*2]; L_216 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd216}: begin L_217 <= data_in[quan_width-1:0]; L_218 <= data_in[quan_width*2-1:quan_width]; L_219 <= data_in[quan_width*3-1:quan_width*2]; L_220 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd220}: begin L_221 <= data_in[quan_width-1:0]; L_222 <= data_in[quan_width*2-1:quan_width]; L_223 <= data_in[quan_width*3-1:quan_width*2]; L_224 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd224}: begin L_225 <= data_in[quan_width-1:0]; L_226 <= data_in[quan_width*2-1:quan_width]; L_227 <= data_in[quan_width*3-1:quan_width*2]; L_228 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd228}: begin L_229 <= data_in[quan_width-1:0]; L_230 <= data_in[quan_width*2-1:quan_width]; L_231 <= data_in[quan_width*3-1:quan_width*2]; L_232 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd232}: begin L_233 <= data_in[quan_width-1:0]; L_234 <= data_in[quan_width*2-1:quan_width]; L_235 <= data_in[quan_width*3-1:quan_width*2]; L_236 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd236}: begin L_237 <= data_in[quan_width-1:0]; L_238 <= data_in[quan_width*2-1:quan_width]; L_239 <= data_in[quan_width*3-1:quan_width*2]; L_240 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd240}: begin L_241 <= data_in[quan_width-1:0]; L_242 <= data_in[quan_width*2-1:quan_width]; L_243 <= data_in[quan_width*3-1:quan_width*2]; L_244 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd244}: begin L_245 <= data_in[quan_width-1:0]; L_246 <= data_in[quan_width*2-1:quan_width]; L_247 <= data_in[quan_width*3-1:quan_width*2]; L_248 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd248}: begin L_249 <= data_in[quan_width-1:0]; L_250 <= data_in[quan_width*2-1:quan_width]; L_251 <= data_in[quan_width*3-1:quan_width*2]; L_252 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd252}: begin L_253 <= data_in[quan_width-1:0]; L_254 <= data_in[quan_width*2-1:quan_width]; L_255 <= data_in[quan_width*3-1:quan_width*2]; L_256 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd256}: begin L_257 <= data_in[quan_width-1:0]; L_258 <= data_in[quan_width*2-1:quan_width]; L_259 <= data_in[quan_width*3-1:quan_width*2]; L_260 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd260}: begin L_261 <= data_in[quan_width-1:0]; L_262 <= data_in[quan_width*2-1:quan_width]; L_263 <= data_in[quan_width*3-1:quan_width*2]; L_264 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd264}: begin L_265 <= data_in[quan_width-1:0]; L_266 <= data_in[quan_width*2-1:quan_width]; L_267 <= data_in[quan_width*3-1:quan_width*2]; L_268 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd268}: begin L_269 <= data_in[quan_width-1:0]; L_270 <= data_in[quan_width*2-1:quan_width]; L_271 <= data_in[quan_width*3-1:quan_width*2]; L_272 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd272}: begin L_273 <= data_in[quan_width-1:0]; L_274 <= data_in[quan_width*2-1:quan_width]; L_275 <= data_in[quan_width*3-1:quan_width*2]; L_276 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd276}: begin L_277 <= data_in[quan_width-1:0]; L_278 <= data_in[quan_width*2-1:quan_width]; L_279 <= data_in[quan_width*3-1:quan_width*2]; L_280 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd280}: begin L_281 <= data_in[quan_width-1:0]; L_282 <= data_in[quan_width*2-1:quan_width]; L_283 <= data_in[quan_width*3-1:quan_width*2]; L_284 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd284}: begin L_285 <= data_in[quan_width-1:0]; L_286 <= data_in[quan_width*2-1:quan_width]; L_287 <= data_in[quan_width*3-1:quan_width*2]; L_288 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd288}: begin L_289 <= data_in[quan_width-1:0]; L_290 <= data_in[quan_width*2-1:quan_width]; L_291 <= data_in[quan_width*3-1:quan_width*2]; L_292 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd292}: begin L_293 <= data_in[quan_width-1:0]; L_294 <= data_in[quan_width*2-1:quan_width]; L_295 <= data_in[quan_width*3-1:quan_width*2]; L_296 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd296}: begin L_297 <= data_in[quan_width-1:0]; L_298 <= data_in[quan_width*2-1:quan_width]; L_299 <= data_in[quan_width*3-1:quan_width*2]; L_300 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd300}: begin L_301 <= data_in[quan_width-1:0]; L_302 <= data_in[quan_width*2-1:quan_width]; L_303 <= data_in[quan_width*3-1:quan_width*2]; L_304 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd304}: begin L_305 <= data_in[quan_width-1:0]; L_306 <= data_in[quan_width*2-1:quan_width]; L_307 <= data_in[quan_width*3-1:quan_width*2]; L_308 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd308}: begin L_309 <= data_in[quan_width-1:0]; L_310 <= data_in[quan_width*2-1:quan_width]; L_311 <= data_in[quan_width*3-1:quan_width*2]; L_312 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd312}: begin L_313 <= data_in[quan_width-1:0]; L_314 <= data_in[quan_width*2-1:quan_width]; L_315 <= data_in[quan_width*3-1:quan_width*2]; L_316 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd316}: begin L_317 <= data_in[quan_width-1:0]; L_318 <= data_in[quan_width*2-1:quan_width]; L_319 <= data_in[quan_width*3-1:quan_width*2]; L_320 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd320}: begin L_321 <= data_in[quan_width-1:0]; L_322 <= data_in[quan_width*2-1:quan_width]; L_323 <= data_in[quan_width*3-1:quan_width*2]; L_324 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd324}: begin L_325 <= data_in[quan_width-1:0]; L_326 <= data_in[quan_width*2-1:quan_width]; L_327 <= data_in[quan_width*3-1:quan_width*2]; L_328 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd328}: begin L_329 <= data_in[quan_width-1:0]; L_330 <= data_in[quan_width*2-1:quan_width]; L_331 <= data_in[quan_width*3-1:quan_width*2]; L_332 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd332}: begin L_333 <= data_in[quan_width-1:0]; L_334 <= data_in[quan_width*2-1:quan_width]; L_335 <= data_in[quan_width*3-1:quan_width*2]; L_336 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd336}: begin L_337 <= data_in[quan_width-1:0]; L_338 <= data_in[quan_width*2-1:quan_width]; L_339 <= data_in[quan_width*3-1:quan_width*2]; L_340 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd340}: begin L_341 <= data_in[quan_width-1:0]; L_342 <= data_in[quan_width*2-1:quan_width]; L_343 <= data_in[quan_width*3-1:quan_width*2]; L_344 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd344}: begin L_345 <= data_in[quan_width-1:0]; L_346 <= data_in[quan_width*2-1:quan_width]; L_347 <= data_in[quan_width*3-1:quan_width*2]; L_348 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd348}: begin L_349 <= data_in[quan_width-1:0]; L_350 <= data_in[quan_width*2-1:quan_width]; L_351 <= data_in[quan_width*3-1:quan_width*2]; L_352 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd352}: begin L_353 <= data_in[quan_width-1:0]; L_354 <= data_in[quan_width*2-1:quan_width]; L_355 <= data_in[quan_width*3-1:quan_width*2]; L_356 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd356}: begin L_357 <= data_in[quan_width-1:0]; L_358 <= data_in[quan_width*2-1:quan_width]; L_359 <= data_in[quan_width*3-1:quan_width*2]; L_360 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd360}: begin L_361 <= data_in[quan_width-1:0]; L_362 <= data_in[quan_width*2-1:quan_width]; L_363 <= data_in[quan_width*3-1:quan_width*2]; L_364 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd364}: begin L_365 <= data_in[quan_width-1:0]; L_366 <= data_in[quan_width*2-1:quan_width]; L_367 <= data_in[quan_width*3-1:quan_width*2]; L_368 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd368}: begin L_369 <= data_in[quan_width-1:0]; L_370 <= data_in[quan_width*2-1:quan_width]; L_371 <= data_in[quan_width*3-1:quan_width*2]; L_372 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd372}: begin L_373 <= data_in[quan_width-1:0]; L_374 <= data_in[quan_width*2-1:quan_width]; L_375 <= data_in[quan_width*3-1:quan_width*2]; L_376 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd376}: begin L_377 <= data_in[quan_width-1:0]; L_378 <= data_in[quan_width*2-1:quan_width]; L_379 <= data_in[quan_width*3-1:quan_width*2]; L_380 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd380}: begin L_381 <= data_in[quan_width-1:0]; L_382 <= data_in[quan_width*2-1:quan_width]; L_383 <= data_in[quan_width*3-1:quan_width*2]; L_384 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd384}: begin L_385 <= data_in[quan_width-1:0]; L_386 <= data_in[quan_width*2-1:quan_width]; L_387 <= data_in[quan_width*3-1:quan_width*2]; L_388 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd388}: begin L_389 <= data_in[quan_width-1:0]; L_390 <= data_in[quan_width*2-1:quan_width]; L_391 <= data_in[quan_width*3-1:quan_width*2]; L_392 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd392}: begin L_393 <= data_in[quan_width-1:0]; L_394 <= data_in[quan_width*2-1:quan_width]; L_395 <= data_in[quan_width*3-1:quan_width*2]; L_396 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd396}: begin L_397 <= data_in[quan_width-1:0]; L_398 <= data_in[quan_width*2-1:quan_width]; L_399 <= data_in[quan_width*3-1:quan_width*2]; L_400 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd400}: begin L_401 <= data_in[quan_width-1:0]; L_402 <= data_in[quan_width*2-1:quan_width]; L_403 <= data_in[quan_width*3-1:quan_width*2]; L_404 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd404}: begin L_405 <= data_in[quan_width-1:0]; L_406 <= data_in[quan_width*2-1:quan_width]; L_407 <= data_in[quan_width*3-1:quan_width*2]; L_408 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd408}: begin L_409 <= data_in[quan_width-1:0]; L_410 <= data_in[quan_width*2-1:quan_width]; L_411 <= data_in[quan_width*3-1:quan_width*2]; L_412 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd412}: begin L_413 <= data_in[quan_width-1:0]; L_414 <= data_in[quan_width*2-1:quan_width]; L_415 <= data_in[quan_width*3-1:quan_width*2]; L_416 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd416}: begin L_417 <= data_in[quan_width-1:0]; L_418 <= data_in[quan_width*2-1:quan_width]; L_419 <= data_in[quan_width*3-1:quan_width*2]; L_420 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd420}: begin L_421 <= data_in[quan_width-1:0]; L_422 <= data_in[quan_width*2-1:quan_width]; L_423 <= data_in[quan_width*3-1:quan_width*2]; L_424 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd424}: begin L_425 <= data_in[quan_width-1:0]; L_426 <= data_in[quan_width*2-1:quan_width]; L_427 <= data_in[quan_width*3-1:quan_width*2]; L_428 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd428}: begin L_429 <= data_in[quan_width-1:0]; L_430 <= data_in[quan_width*2-1:quan_width]; L_431 <= data_in[quan_width*3-1:quan_width*2]; L_432 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd432}: begin L_433 <= data_in[quan_width-1:0]; L_434 <= data_in[quan_width*2-1:quan_width]; L_435 <= data_in[quan_width*3-1:quan_width*2]; L_436 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd436}: begin L_437 <= data_in[quan_width-1:0]; L_438 <= data_in[quan_width*2-1:quan_width]; L_439 <= data_in[quan_width*3-1:quan_width*2]; L_440 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd440}: begin L_441 <= data_in[quan_width-1:0]; L_442 <= data_in[quan_width*2-1:quan_width]; L_443 <= data_in[quan_width*3-1:quan_width*2]; L_444 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd444}: begin L_445 <= data_in[quan_width-1:0]; L_446 <= data_in[quan_width*2-1:quan_width]; L_447 <= data_in[quan_width*3-1:quan_width*2]; L_448 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd448}: begin L_449 <= data_in[quan_width-1:0]; L_450 <= data_in[quan_width*2-1:quan_width]; L_451 <= data_in[quan_width*3-1:quan_width*2]; L_452 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd452}: begin L_453 <= data_in[quan_width-1:0]; L_454 <= data_in[quan_width*2-1:quan_width]; L_455 <= data_in[quan_width*3-1:quan_width*2]; L_456 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd456}: begin L_457 <= data_in[quan_width-1:0]; L_458 <= data_in[quan_width*2-1:quan_width]; L_459 <= data_in[quan_width*3-1:quan_width*2]; L_460 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd460}: begin L_461 <= data_in[quan_width-1:0]; L_462 <= data_in[quan_width*2-1:quan_width]; L_463 <= data_in[quan_width*3-1:quan_width*2]; L_464 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd464}: begin L_465 <= data_in[quan_width-1:0]; L_466 <= data_in[quan_width*2-1:quan_width]; L_467 <= data_in[quan_width*3-1:quan_width*2]; L_468 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd468}: begin L_469 <= data_in[quan_width-1:0]; L_470 <= data_in[quan_width*2-1:quan_width]; L_471 <= data_in[quan_width*3-1:quan_width*2]; L_472 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd472}: begin L_473 <= data_in[quan_width-1:0]; L_474 <= data_in[quan_width*2-1:quan_width]; L_475 <= data_in[quan_width*3-1:quan_width*2]; L_476 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd476}: begin L_477 <= data_in[quan_width-1:0]; L_478 <= data_in[quan_width*2-1:quan_width]; L_479 <= data_in[quan_width*3-1:quan_width*2]; L_480 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd480}: begin L_481 <= data_in[quan_width-1:0]; L_482 <= data_in[quan_width*2-1:quan_width]; L_483 <= data_in[quan_width*3-1:quan_width*2]; L_484 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd484}: begin L_485 <= data_in[quan_width-1:0]; L_486 <= data_in[quan_width*2-1:quan_width]; L_487 <= data_in[quan_width*3-1:quan_width*2]; L_488 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd488}: begin L_489 <= data_in[quan_width-1:0]; L_490 <= data_in[quan_width*2-1:quan_width]; L_491 <= data_in[quan_width*3-1:quan_width*2]; L_492 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd492}: begin L_493 <= data_in[quan_width-1:0]; L_494 <= data_in[quan_width*2-1:quan_width]; L_495 <= data_in[quan_width*3-1:quan_width*2]; L_496 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd496}: begin L_497 <= data_in[quan_width-1:0]; L_498 <= data_in[quan_width*2-1:quan_width]; L_499 <= data_in[quan_width*3-1:quan_width*2]; L_500 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd500}: begin L_501 <= data_in[quan_width-1:0]; L_502 <= data_in[quan_width*2-1:quan_width]; L_503 <= data_in[quan_width*3-1:quan_width*2]; L_504 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd504}: begin L_505 <= data_in[quan_width-1:0]; L_506 <= data_in[quan_width*2-1:quan_width]; L_507 <= data_in[quan_width*3-1:quan_width*2]; L_508 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd508}: begin L_509 <= data_in[quan_width-1:0]; L_510 <= data_in[quan_width*2-1:quan_width]; L_511 <= data_in[quan_width*3-1:quan_width*2]; L_512 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd512}: begin L_513 <= data_in[quan_width-1:0]; L_514 <= data_in[quan_width*2-1:quan_width]; L_515 <= data_in[quan_width*3-1:quan_width*2]; L_516 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd516}: begin L_517 <= data_in[quan_width-1:0]; L_518 <= data_in[quan_width*2-1:quan_width]; L_519 <= data_in[quan_width*3-1:quan_width*2]; L_520 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd520}: begin L_521 <= data_in[quan_width-1:0]; L_522 <= data_in[quan_width*2-1:quan_width]; L_523 <= data_in[quan_width*3-1:quan_width*2]; L_524 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd524}: begin L_525 <= data_in[quan_width-1:0]; L_526 <= data_in[quan_width*2-1:quan_width]; L_527 <= data_in[quan_width*3-1:quan_width*2]; L_528 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd528}: begin L_529 <= data_in[quan_width-1:0]; L_530 <= data_in[quan_width*2-1:quan_width]; L_531 <= data_in[quan_width*3-1:quan_width*2]; L_532 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd532}: begin L_533 <= data_in[quan_width-1:0]; L_534 <= data_in[quan_width*2-1:quan_width]; L_535 <= data_in[quan_width*3-1:quan_width*2]; L_536 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd536}: begin L_537 <= data_in[quan_width-1:0]; L_538 <= data_in[quan_width*2-1:quan_width]; L_539 <= data_in[quan_width*3-1:quan_width*2]; L_540 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd540}: begin L_541 <= data_in[quan_width-1:0]; L_542 <= data_in[quan_width*2-1:quan_width]; L_543 <= data_in[quan_width*3-1:quan_width*2]; L_544 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd544}: begin L_545 <= data_in[quan_width-1:0]; L_546 <= data_in[quan_width*2-1:quan_width]; L_547 <= data_in[quan_width*3-1:quan_width*2]; L_548 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd548}: begin L_549 <= data_in[quan_width-1:0]; L_550 <= data_in[quan_width*2-1:quan_width]; L_551 <= data_in[quan_width*3-1:quan_width*2]; L_552 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd552}: begin L_553 <= data_in[quan_width-1:0]; L_554 <= data_in[quan_width*2-1:quan_width]; L_555 <= data_in[quan_width*3-1:quan_width*2]; L_556 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd556}: begin L_557 <= data_in[quan_width-1:0]; L_558 <= data_in[quan_width*2-1:quan_width]; L_559 <= data_in[quan_width*3-1:quan_width*2]; L_560 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd560}: begin L_561 <= data_in[quan_width-1:0]; L_562 <= data_in[quan_width*2-1:quan_width]; L_563 <= data_in[quan_width*3-1:quan_width*2]; L_564 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd564}: begin L_565 <= data_in[quan_width-1:0]; L_566 <= data_in[quan_width*2-1:quan_width]; L_567 <= data_in[quan_width*3-1:quan_width*2]; L_568 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd568}: begin L_569 <= data_in[quan_width-1:0]; L_570 <= data_in[quan_width*2-1:quan_width]; L_571 <= data_in[quan_width*3-1:quan_width*2]; L_572 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd572}: begin L_573 <= data_in[quan_width-1:0]; L_574 <= data_in[quan_width*2-1:quan_width]; L_575 <= data_in[quan_width*3-1:quan_width*2]; L_576 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd576}: begin L_577 <= data_in[quan_width-1:0]; L_578 <= data_in[quan_width*2-1:quan_width]; L_579 <= data_in[quan_width*3-1:quan_width*2]; L_580 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd580}: begin L_581 <= data_in[quan_width-1:0]; L_582 <= data_in[quan_width*2-1:quan_width]; L_583 <= data_in[quan_width*3-1:quan_width*2]; L_584 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd584}: begin L_585 <= data_in[quan_width-1:0]; L_586 <= data_in[quan_width*2-1:quan_width]; L_587 <= data_in[quan_width*3-1:quan_width*2]; L_588 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd588}: begin L_589 <= data_in[quan_width-1:0]; L_590 <= data_in[quan_width*2-1:quan_width]; L_591 <= data_in[quan_width*3-1:quan_width*2]; L_592 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd592}: begin L_593 <= data_in[quan_width-1:0]; L_594 <= data_in[quan_width*2-1:quan_width]; L_595 <= data_in[quan_width*3-1:quan_width*2]; L_596 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd596}: begin L_597 <= data_in[quan_width-1:0]; L_598 <= data_in[quan_width*2-1:quan_width]; L_599 <= data_in[quan_width*3-1:quan_width*2]; L_600 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd600}: begin L_601 <= data_in[quan_width-1:0]; L_602 <= data_in[quan_width*2-1:quan_width]; L_603 <= data_in[quan_width*3-1:quan_width*2]; L_604 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd604}: begin L_605 <= data_in[quan_width-1:0]; L_606 <= data_in[quan_width*2-1:quan_width]; L_607 <= data_in[quan_width*3-1:quan_width*2]; L_608 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd608}: begin L_609 <= data_in[quan_width-1:0]; L_610 <= data_in[quan_width*2-1:quan_width]; L_611 <= data_in[quan_width*3-1:quan_width*2]; L_612 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd612}: begin L_613 <= data_in[quan_width-1:0]; L_614 <= data_in[quan_width*2-1:quan_width]; L_615 <= data_in[quan_width*3-1:quan_width*2]; L_616 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd616}: begin L_617 <= data_in[quan_width-1:0]; L_618 <= data_in[quan_width*2-1:quan_width]; L_619 <= data_in[quan_width*3-1:quan_width*2]; L_620 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd620}: begin L_621 <= data_in[quan_width-1:0]; L_622 <= data_in[quan_width*2-1:quan_width]; L_623 <= data_in[quan_width*3-1:quan_width*2]; L_624 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd624}: begin L_625 <= data_in[quan_width-1:0]; L_626 <= data_in[quan_width*2-1:quan_width]; L_627 <= data_in[quan_width*3-1:quan_width*2]; L_628 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd628}: begin L_629 <= data_in[quan_width-1:0]; L_630 <= data_in[quan_width*2-1:quan_width]; L_631 <= data_in[quan_width*3-1:quan_width*2]; L_632 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd632}: begin L_633 <= data_in[quan_width-1:0]; L_634 <= data_in[quan_width*2-1:quan_width]; L_635 <= data_in[quan_width*3-1:quan_width*2]; L_636 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd636}: begin L_637 <= data_in[quan_width-1:0]; L_638 <= data_in[quan_width*2-1:quan_width]; L_639 <= data_in[quan_width*3-1:quan_width*2]; L_640 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd640}: begin L_641 <= data_in[quan_width-1:0]; L_642 <= data_in[quan_width*2-1:quan_width]; L_643 <= data_in[quan_width*3-1:quan_width*2]; L_644 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd644}: begin L_645 <= data_in[quan_width-1:0]; L_646 <= data_in[quan_width*2-1:quan_width]; L_647 <= data_in[quan_width*3-1:quan_width*2]; L_648 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd648}: begin L_649 <= data_in[quan_width-1:0]; L_650 <= data_in[quan_width*2-1:quan_width]; L_651 <= data_in[quan_width*3-1:quan_width*2]; L_652 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd652}: begin L_653 <= data_in[quan_width-1:0]; L_654 <= data_in[quan_width*2-1:quan_width]; L_655 <= data_in[quan_width*3-1:quan_width*2]; L_656 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd656}: begin L_657 <= data_in[quan_width-1:0]; L_658 <= data_in[quan_width*2-1:quan_width]; L_659 <= data_in[quan_width*3-1:quan_width*2]; L_660 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd660}: begin L_661 <= data_in[quan_width-1:0]; L_662 <= data_in[quan_width*2-1:quan_width]; L_663 <= data_in[quan_width*3-1:quan_width*2]; L_664 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd664}: begin L_665 <= data_in[quan_width-1:0]; L_666 <= data_in[quan_width*2-1:quan_width]; L_667 <= data_in[quan_width*3-1:quan_width*2]; L_668 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd668}: begin L_669 <= data_in[quan_width-1:0]; L_670 <= data_in[quan_width*2-1:quan_width]; L_671 <= data_in[quan_width*3-1:quan_width*2]; L_672 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd672}: begin L_673 <= data_in[quan_width-1:0]; L_674 <= data_in[quan_width*2-1:quan_width]; L_675 <= data_in[quan_width*3-1:quan_width*2]; L_676 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd676}: begin L_677 <= data_in[quan_width-1:0]; L_678 <= data_in[quan_width*2-1:quan_width]; L_679 <= data_in[quan_width*3-1:quan_width*2]; L_680 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd680}: begin L_681 <= data_in[quan_width-1:0]; L_682 <= data_in[quan_width*2-1:quan_width]; L_683 <= data_in[quan_width*3-1:quan_width*2]; L_684 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd684}: begin L_685 <= data_in[quan_width-1:0]; L_686 <= data_in[quan_width*2-1:quan_width]; L_687 <= data_in[quan_width*3-1:quan_width*2]; L_688 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd688}: begin L_689 <= data_in[quan_width-1:0]; L_690 <= data_in[quan_width*2-1:quan_width]; L_691 <= data_in[quan_width*3-1:quan_width*2]; L_692 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd692}: begin L_693 <= data_in[quan_width-1:0]; L_694 <= data_in[quan_width*2-1:quan_width]; L_695 <= data_in[quan_width*3-1:quan_width*2]; L_696 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd696}: begin L_697 <= data_in[quan_width-1:0]; L_698 <= data_in[quan_width*2-1:quan_width]; L_699 <= data_in[quan_width*3-1:quan_width*2]; L_700 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd700}: begin L_701 <= data_in[quan_width-1:0]; L_702 <= data_in[quan_width*2-1:quan_width]; L_703 <= data_in[quan_width*3-1:quan_width*2]; L_704 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd704}: begin L_705 <= data_in[quan_width-1:0]; L_706 <= data_in[quan_width*2-1:quan_width]; L_707 <= data_in[quan_width*3-1:quan_width*2]; L_708 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd708}: begin L_709 <= data_in[quan_width-1:0]; L_710 <= data_in[quan_width*2-1:quan_width]; L_711 <= data_in[quan_width*3-1:quan_width*2]; L_712 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd712}: begin L_713 <= data_in[quan_width-1:0]; L_714 <= data_in[quan_width*2-1:quan_width]; L_715 <= data_in[quan_width*3-1:quan_width*2]; L_716 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd716}: begin L_717 <= data_in[quan_width-1:0]; L_718 <= data_in[quan_width*2-1:quan_width]; L_719 <= data_in[quan_width*3-1:quan_width*2]; L_720 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd720}: begin L_721 <= data_in[quan_width-1:0]; L_722 <= data_in[quan_width*2-1:quan_width]; L_723 <= data_in[quan_width*3-1:quan_width*2]; L_724 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd724}: begin L_725 <= data_in[quan_width-1:0]; L_726 <= data_in[quan_width*2-1:quan_width]; L_727 <= data_in[quan_width*3-1:quan_width*2]; L_728 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd728}: begin L_729 <= data_in[quan_width-1:0]; L_730 <= data_in[quan_width*2-1:quan_width]; L_731 <= data_in[quan_width*3-1:quan_width*2]; L_732 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd732}: begin L_733 <= data_in[quan_width-1:0]; L_734 <= data_in[quan_width*2-1:quan_width]; L_735 <= data_in[quan_width*3-1:quan_width*2]; L_736 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd736}: begin L_737 <= data_in[quan_width-1:0]; L_738 <= data_in[quan_width*2-1:quan_width]; L_739 <= data_in[quan_width*3-1:quan_width*2]; L_740 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd740}: begin L_741 <= data_in[quan_width-1:0]; L_742 <= data_in[quan_width*2-1:quan_width]; L_743 <= data_in[quan_width*3-1:quan_width*2]; L_744 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd744}: begin L_745 <= data_in[quan_width-1:0]; L_746 <= data_in[quan_width*2-1:quan_width]; L_747 <= data_in[quan_width*3-1:quan_width*2]; L_748 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd748}: begin L_749 <= data_in[quan_width-1:0]; L_750 <= data_in[quan_width*2-1:quan_width]; L_751 <= data_in[quan_width*3-1:quan_width*2]; L_752 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd752}: begin L_753 <= data_in[quan_width-1:0]; L_754 <= data_in[quan_width*2-1:quan_width]; L_755 <= data_in[quan_width*3-1:quan_width*2]; L_756 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd756}: begin L_757 <= data_in[quan_width-1:0]; L_758 <= data_in[quan_width*2-1:quan_width]; L_759 <= data_in[quan_width*3-1:quan_width*2]; L_760 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd760}: begin L_761 <= data_in[quan_width-1:0]; L_762 <= data_in[quan_width*2-1:quan_width]; L_763 <= data_in[quan_width*3-1:quan_width*2]; L_764 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd764}: begin L_765 <= data_in[quan_width-1:0]; L_766 <= data_in[quan_width*2-1:quan_width]; L_767 <= data_in[quan_width*3-1:quan_width*2]; L_768 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd768}: begin L_769 <= data_in[quan_width-1:0]; L_770 <= data_in[quan_width*2-1:quan_width]; L_771 <= data_in[quan_width*3-1:quan_width*2]; L_772 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd772}: begin L_773 <= data_in[quan_width-1:0]; L_774 <= data_in[quan_width*2-1:quan_width]; L_775 <= data_in[quan_width*3-1:quan_width*2]; L_776 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd776}: begin L_777 <= data_in[quan_width-1:0]; L_778 <= data_in[quan_width*2-1:quan_width]; L_779 <= data_in[quan_width*3-1:quan_width*2]; L_780 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd780}: begin L_781 <= data_in[quan_width-1:0]; L_782 <= data_in[quan_width*2-1:quan_width]; L_783 <= data_in[quan_width*3-1:quan_width*2]; L_784 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd784}: begin L_785 <= data_in[quan_width-1:0]; L_786 <= data_in[quan_width*2-1:quan_width]; L_787 <= data_in[quan_width*3-1:quan_width*2]; L_788 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd788}: begin L_789 <= data_in[quan_width-1:0]; L_790 <= data_in[quan_width*2-1:quan_width]; L_791 <= data_in[quan_width*3-1:quan_width*2]; L_792 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd792}: begin L_793 <= data_in[quan_width-1:0]; L_794 <= data_in[quan_width*2-1:quan_width]; L_795 <= data_in[quan_width*3-1:quan_width*2]; L_796 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd796}: begin L_797 <= data_in[quan_width-1:0]; L_798 <= data_in[quan_width*2-1:quan_width]; L_799 <= data_in[quan_width*3-1:quan_width*2]; L_800 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd800}: begin L_801 <= data_in[quan_width-1:0]; L_802 <= data_in[quan_width*2-1:quan_width]; L_803 <= data_in[quan_width*3-1:quan_width*2]; L_804 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd804}: begin L_805 <= data_in[quan_width-1:0]; L_806 <= data_in[quan_width*2-1:quan_width]; L_807 <= data_in[quan_width*3-1:quan_width*2]; L_808 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd808}: begin L_809 <= data_in[quan_width-1:0]; L_810 <= data_in[quan_width*2-1:quan_width]; L_811 <= data_in[quan_width*3-1:quan_width*2]; L_812 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd812}: begin L_813 <= data_in[quan_width-1:0]; L_814 <= data_in[quan_width*2-1:quan_width]; L_815 <= data_in[quan_width*3-1:quan_width*2]; L_816 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd816}: begin L_817 <= data_in[quan_width-1:0]; L_818 <= data_in[quan_width*2-1:quan_width]; L_819 <= data_in[quan_width*3-1:quan_width*2]; L_820 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd820}: begin L_821 <= data_in[quan_width-1:0]; L_822 <= data_in[quan_width*2-1:quan_width]; L_823 <= data_in[quan_width*3-1:quan_width*2]; L_824 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd824}: begin L_825 <= data_in[quan_width-1:0]; L_826 <= data_in[quan_width*2-1:quan_width]; L_827 <= data_in[quan_width*3-1:quan_width*2]; L_828 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd828}: begin L_829 <= data_in[quan_width-1:0]; L_830 <= data_in[quan_width*2-1:quan_width]; L_831 <= data_in[quan_width*3-1:quan_width*2]; L_832 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd832}: begin L_833 <= data_in[quan_width-1:0]; L_834 <= data_in[quan_width*2-1:quan_width]; L_835 <= data_in[quan_width*3-1:quan_width*2]; L_836 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd836}: begin L_837 <= data_in[quan_width-1:0]; L_838 <= data_in[quan_width*2-1:quan_width]; L_839 <= data_in[quan_width*3-1:quan_width*2]; L_840 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd840}: begin L_841 <= data_in[quan_width-1:0]; L_842 <= data_in[quan_width*2-1:quan_width]; L_843 <= data_in[quan_width*3-1:quan_width*2]; L_844 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd844}: begin L_845 <= data_in[quan_width-1:0]; L_846 <= data_in[quan_width*2-1:quan_width]; L_847 <= data_in[quan_width*3-1:quan_width*2]; L_848 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd848}: begin L_849 <= data_in[quan_width-1:0]; L_850 <= data_in[quan_width*2-1:quan_width]; L_851 <= data_in[quan_width*3-1:quan_width*2]; L_852 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd852}: begin L_853 <= data_in[quan_width-1:0]; L_854 <= data_in[quan_width*2-1:quan_width]; L_855 <= data_in[quan_width*3-1:quan_width*2]; L_856 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd856}: begin L_857 <= data_in[quan_width-1:0]; L_858 <= data_in[quan_width*2-1:quan_width]; L_859 <= data_in[quan_width*3-1:quan_width*2]; L_860 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd860}: begin L_861 <= data_in[quan_width-1:0]; L_862 <= data_in[quan_width*2-1:quan_width]; L_863 <= data_in[quan_width*3-1:quan_width*2]; L_864 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd864}: begin L_865 <= data_in[quan_width-1:0]; L_866 <= data_in[quan_width*2-1:quan_width]; L_867 <= data_in[quan_width*3-1:quan_width*2]; L_868 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd868}: begin L_869 <= data_in[quan_width-1:0]; L_870 <= data_in[quan_width*2-1:quan_width]; L_871 <= data_in[quan_width*3-1:quan_width*2]; L_872 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd872}: begin L_873 <= data_in[quan_width-1:0]; L_874 <= data_in[quan_width*2-1:quan_width]; L_875 <= data_in[quan_width*3-1:quan_width*2]; L_876 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd876}: begin L_877 <= data_in[quan_width-1:0]; L_878 <= data_in[quan_width*2-1:quan_width]; L_879 <= data_in[quan_width*3-1:quan_width*2]; L_880 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd880}: begin L_881 <= data_in[quan_width-1:0]; L_882 <= data_in[quan_width*2-1:quan_width]; L_883 <= data_in[quan_width*3-1:quan_width*2]; L_884 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd884}: begin L_885 <= data_in[quan_width-1:0]; L_886 <= data_in[quan_width*2-1:quan_width]; L_887 <= data_in[quan_width*3-1:quan_width*2]; L_888 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd888}: begin L_889 <= data_in[quan_width-1:0]; L_890 <= data_in[quan_width*2-1:quan_width]; L_891 <= data_in[quan_width*3-1:quan_width*2]; L_892 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd892}: begin L_893 <= data_in[quan_width-1:0]; L_894 <= data_in[quan_width*2-1:quan_width]; L_895 <= data_in[quan_width*3-1:quan_width*2]; L_896 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd896}: begin L_897 <= data_in[quan_width-1:0]; L_898 <= data_in[quan_width*2-1:quan_width]; L_899 <= data_in[quan_width*3-1:quan_width*2]; L_900 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd900}: begin L_901 <= data_in[quan_width-1:0]; L_902 <= data_in[quan_width*2-1:quan_width]; L_903 <= data_in[quan_width*3-1:quan_width*2]; L_904 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd904}: begin L_905 <= data_in[quan_width-1:0]; L_906 <= data_in[quan_width*2-1:quan_width]; L_907 <= data_in[quan_width*3-1:quan_width*2]; L_908 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd908}: begin L_909 <= data_in[quan_width-1:0]; L_910 <= data_in[quan_width*2-1:quan_width]; L_911 <= data_in[quan_width*3-1:quan_width*2]; L_912 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd912}: begin L_913 <= data_in[quan_width-1:0]; L_914 <= data_in[quan_width*2-1:quan_width]; L_915 <= data_in[quan_width*3-1:quan_width*2]; L_916 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd916}: begin L_917 <= data_in[quan_width-1:0]; L_918 <= data_in[quan_width*2-1:quan_width]; L_919 <= data_in[quan_width*3-1:quan_width*2]; L_920 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd920}: begin L_921 <= data_in[quan_width-1:0]; L_922 <= data_in[quan_width*2-1:quan_width]; L_923 <= data_in[quan_width*3-1:quan_width*2]; L_924 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd924}: begin L_925 <= data_in[quan_width-1:0]; L_926 <= data_in[quan_width*2-1:quan_width]; L_927 <= data_in[quan_width*3-1:quan_width*2]; L_928 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd928}: begin L_929 <= data_in[quan_width-1:0]; L_930 <= data_in[quan_width*2-1:quan_width]; L_931 <= data_in[quan_width*3-1:quan_width*2]; L_932 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd932}: begin L_933 <= data_in[quan_width-1:0]; L_934 <= data_in[quan_width*2-1:quan_width]; L_935 <= data_in[quan_width*3-1:quan_width*2]; L_936 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd936}: begin L_937 <= data_in[quan_width-1:0]; L_938 <= data_in[quan_width*2-1:quan_width]; L_939 <= data_in[quan_width*3-1:quan_width*2]; L_940 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd940}: begin L_941 <= data_in[quan_width-1:0]; L_942 <= data_in[quan_width*2-1:quan_width]; L_943 <= data_in[quan_width*3-1:quan_width*2]; L_944 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd944}: begin L_945 <= data_in[quan_width-1:0]; L_946 <= data_in[quan_width*2-1:quan_width]; L_947 <= data_in[quan_width*3-1:quan_width*2]; L_948 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd948}: begin L_949 <= data_in[quan_width-1:0]; L_950 <= data_in[quan_width*2-1:quan_width]; L_951 <= data_in[quan_width*3-1:quan_width*2]; L_952 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd952}: begin L_953 <= data_in[quan_width-1:0]; L_954 <= data_in[quan_width*2-1:quan_width]; L_955 <= data_in[quan_width*3-1:quan_width*2]; L_956 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd956}: begin L_957 <= data_in[quan_width-1:0]; L_958 <= data_in[quan_width*2-1:quan_width]; L_959 <= data_in[quan_width*3-1:quan_width*2]; L_960 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd960}: begin L_961 <= data_in[quan_width-1:0]; L_962 <= data_in[quan_width*2-1:quan_width]; L_963 <= data_in[quan_width*3-1:quan_width*2]; L_964 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd964}: begin L_965 <= data_in[quan_width-1:0]; L_966 <= data_in[quan_width*2-1:quan_width]; L_967 <= data_in[quan_width*3-1:quan_width*2]; L_968 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd968}: begin L_969 <= data_in[quan_width-1:0]; L_970 <= data_in[quan_width*2-1:quan_width]; L_971 <= data_in[quan_width*3-1:quan_width*2]; L_972 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd972}: begin L_973 <= data_in[quan_width-1:0]; L_974 <= data_in[quan_width*2-1:quan_width]; L_975 <= data_in[quan_width*3-1:quan_width*2]; L_976 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd976}: begin L_977 <= data_in[quan_width-1:0]; L_978 <= data_in[quan_width*2-1:quan_width]; L_979 <= data_in[quan_width*3-1:quan_width*2]; L_980 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd980}: begin L_981 <= data_in[quan_width-1:0]; L_982 <= data_in[quan_width*2-1:quan_width]; L_983 <= data_in[quan_width*3-1:quan_width*2]; L_984 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd984}: begin L_985 <= data_in[quan_width-1:0]; L_986 <= data_in[quan_width*2-1:quan_width]; L_987 <= data_in[quan_width*3-1:quan_width*2]; L_988 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd988}: begin L_989 <= data_in[quan_width-1:0]; L_990 <= data_in[quan_width*2-1:quan_width]; L_991 <= data_in[quan_width*3-1:quan_width*2]; L_992 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd992}: begin L_993 <= data_in[quan_width-1:0]; L_994 <= data_in[quan_width*2-1:quan_width]; L_995 <= data_in[quan_width*3-1:quan_width*2]; L_996 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd996}: begin L_997 <= data_in[quan_width-1:0]; L_998 <= data_in[quan_width*2-1:quan_width]; L_999 <= data_in[quan_width*3-1:quan_width*2]; L_1000 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1000}: begin L_1001 <= data_in[quan_width-1:0]; L_1002 <= data_in[quan_width*2-1:quan_width]; L_1003 <= data_in[quan_width*3-1:quan_width*2]; L_1004 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1004}: begin L_1005 <= data_in[quan_width-1:0]; L_1006 <= data_in[quan_width*2-1:quan_width]; L_1007 <= data_in[quan_width*3-1:quan_width*2]; L_1008 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1008}: begin L_1009 <= data_in[quan_width-1:0]; L_1010 <= data_in[quan_width*2-1:quan_width]; L_1011 <= data_in[quan_width*3-1:quan_width*2]; L_1012 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1012}: begin L_1013 <= data_in[quan_width-1:0]; L_1014 <= data_in[quan_width*2-1:quan_width]; L_1015 <= data_in[quan_width*3-1:quan_width*2]; L_1016 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1016}: begin L_1017 <= data_in[quan_width-1:0]; L_1018 <= data_in[quan_width*2-1:quan_width]; L_1019 <= data_in[quan_width*3-1:quan_width*2]; L_1020 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1020}: begin L_1021 <= data_in[quan_width-1:0]; L_1022 <= data_in[quan_width*2-1:quan_width]; L_1023 <= data_in[quan_width*3-1:quan_width*2]; L_1024 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1024}: begin L_1025 <= data_in[quan_width-1:0]; L_1026 <= data_in[quan_width*2-1:quan_width]; L_1027 <= data_in[quan_width*3-1:quan_width*2]; L_1028 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1028}: begin L_1029 <= data_in[quan_width-1:0]; L_1030 <= data_in[quan_width*2-1:quan_width]; L_1031 <= data_in[quan_width*3-1:quan_width*2]; L_1032 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1032}: begin L_1033 <= data_in[quan_width-1:0]; L_1034 <= data_in[quan_width*2-1:quan_width]; L_1035 <= data_in[quan_width*3-1:quan_width*2]; L_1036 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1036}: begin L_1037 <= data_in[quan_width-1:0]; L_1038 <= data_in[quan_width*2-1:quan_width]; L_1039 <= data_in[quan_width*3-1:quan_width*2]; L_1040 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1040}: begin L_1041 <= data_in[quan_width-1:0]; L_1042 <= data_in[quan_width*2-1:quan_width]; L_1043 <= data_in[quan_width*3-1:quan_width*2]; L_1044 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1044}: begin L_1045 <= data_in[quan_width-1:0]; L_1046 <= data_in[quan_width*2-1:quan_width]; L_1047 <= data_in[quan_width*3-1:quan_width*2]; L_1048 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1048}: begin L_1049 <= data_in[quan_width-1:0]; L_1050 <= data_in[quan_width*2-1:quan_width]; L_1051 <= data_in[quan_width*3-1:quan_width*2]; L_1052 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1052}: begin L_1053 <= data_in[quan_width-1:0]; L_1054 <= data_in[quan_width*2-1:quan_width]; L_1055 <= data_in[quan_width*3-1:quan_width*2]; L_1056 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1056}: begin L_1057 <= data_in[quan_width-1:0]; L_1058 <= data_in[quan_width*2-1:quan_width]; L_1059 <= data_in[quan_width*3-1:quan_width*2]; L_1060 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1060}: begin L_1061 <= data_in[quan_width-1:0]; L_1062 <= data_in[quan_width*2-1:quan_width]; L_1063 <= data_in[quan_width*3-1:quan_width*2]; L_1064 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1064}: begin L_1065 <= data_in[quan_width-1:0]; L_1066 <= data_in[quan_width*2-1:quan_width]; L_1067 <= data_in[quan_width*3-1:quan_width*2]; L_1068 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1068}: begin L_1069 <= data_in[quan_width-1:0]; L_1070 <= data_in[quan_width*2-1:quan_width]; L_1071 <= data_in[quan_width*3-1:quan_width*2]; L_1072 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1072}: begin L_1073 <= data_in[quan_width-1:0]; L_1074 <= data_in[quan_width*2-1:quan_width]; L_1075 <= data_in[quan_width*3-1:quan_width*2]; L_1076 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1076}: begin L_1077 <= data_in[quan_width-1:0]; L_1078 <= data_in[quan_width*2-1:quan_width]; L_1079 <= data_in[quan_width*3-1:quan_width*2]; L_1080 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1080}: begin L_1081 <= data_in[quan_width-1:0]; L_1082 <= data_in[quan_width*2-1:quan_width]; L_1083 <= data_in[quan_width*3-1:quan_width*2]; L_1084 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1084}: begin L_1085 <= data_in[quan_width-1:0]; L_1086 <= data_in[quan_width*2-1:quan_width]; L_1087 <= data_in[quan_width*3-1:quan_width*2]; L_1088 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1088}: begin L_1089 <= data_in[quan_width-1:0]; L_1090 <= data_in[quan_width*2-1:quan_width]; L_1091 <= data_in[quan_width*3-1:quan_width*2]; L_1092 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1092}: begin L_1093 <= data_in[quan_width-1:0]; L_1094 <= data_in[quan_width*2-1:quan_width]; L_1095 <= data_in[quan_width*3-1:quan_width*2]; L_1096 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1096}: begin L_1097 <= data_in[quan_width-1:0]; L_1098 <= data_in[quan_width*2-1:quan_width]; L_1099 <= data_in[quan_width*3-1:quan_width*2]; L_1100 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1100}: begin L_1101 <= data_in[quan_width-1:0]; L_1102 <= data_in[quan_width*2-1:quan_width]; L_1103 <= data_in[quan_width*3-1:quan_width*2]; L_1104 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1104}: begin L_1105 <= data_in[quan_width-1:0]; L_1106 <= data_in[quan_width*2-1:quan_width]; L_1107 <= data_in[quan_width*3-1:quan_width*2]; L_1108 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1108}: begin L_1109 <= data_in[quan_width-1:0]; L_1110 <= data_in[quan_width*2-1:quan_width]; L_1111 <= data_in[quan_width*3-1:quan_width*2]; L_1112 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1112}: begin L_1113 <= data_in[quan_width-1:0]; L_1114 <= data_in[quan_width*2-1:quan_width]; L_1115 <= data_in[quan_width*3-1:quan_width*2]; L_1116 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1116}: begin L_1117 <= data_in[quan_width-1:0]; L_1118 <= data_in[quan_width*2-1:quan_width]; L_1119 <= data_in[quan_width*3-1:quan_width*2]; L_1120 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1120}: begin L_1121 <= data_in[quan_width-1:0]; L_1122 <= data_in[quan_width*2-1:quan_width]; L_1123 <= data_in[quan_width*3-1:quan_width*2]; L_1124 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1124}: begin L_1125 <= data_in[quan_width-1:0]; L_1126 <= data_in[quan_width*2-1:quan_width]; L_1127 <= data_in[quan_width*3-1:quan_width*2]; L_1128 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1128}: begin L_1129 <= data_in[quan_width-1:0]; L_1130 <= data_in[quan_width*2-1:quan_width]; L_1131 <= data_in[quan_width*3-1:quan_width*2]; L_1132 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1132}: begin L_1133 <= data_in[quan_width-1:0]; L_1134 <= data_in[quan_width*2-1:quan_width]; L_1135 <= data_in[quan_width*3-1:quan_width*2]; L_1136 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1136}: begin L_1137 <= data_in[quan_width-1:0]; L_1138 <= data_in[quan_width*2-1:quan_width]; L_1139 <= data_in[quan_width*3-1:quan_width*2]; L_1140 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1140}: begin L_1141 <= data_in[quan_width-1:0]; L_1142 <= data_in[quan_width*2-1:quan_width]; L_1143 <= data_in[quan_width*3-1:quan_width*2]; L_1144 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1144}: begin L_1145 <= data_in[quan_width-1:0]; L_1146 <= data_in[quan_width*2-1:quan_width]; L_1147 <= data_in[quan_width*3-1:quan_width*2]; L_1148 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1148}: begin L_1149 <= data_in[quan_width-1:0]; L_1150 <= data_in[quan_width*2-1:quan_width]; L_1151 <= data_in[quan_width*3-1:quan_width*2]; L_1152 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1152}: begin L_1153 <= data_in[quan_width-1:0]; L_1154 <= data_in[quan_width*2-1:quan_width]; L_1155 <= data_in[quan_width*3-1:quan_width*2]; L_1156 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1156}: begin L_1157 <= data_in[quan_width-1:0]; L_1158 <= data_in[quan_width*2-1:quan_width]; L_1159 <= data_in[quan_width*3-1:quan_width*2]; L_1160 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1160}: begin L_1161 <= data_in[quan_width-1:0]; L_1162 <= data_in[quan_width*2-1:quan_width]; L_1163 <= data_in[quan_width*3-1:quan_width*2]; L_1164 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1164}: begin L_1165 <= data_in[quan_width-1:0]; L_1166 <= data_in[quan_width*2-1:quan_width]; L_1167 <= data_in[quan_width*3-1:quan_width*2]; L_1168 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1168}: begin L_1169 <= data_in[quan_width-1:0]; L_1170 <= data_in[quan_width*2-1:quan_width]; L_1171 <= data_in[quan_width*3-1:quan_width*2]; L_1172 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1172}: begin L_1173 <= data_in[quan_width-1:0]; L_1174 <= data_in[quan_width*2-1:quan_width]; L_1175 <= data_in[quan_width*3-1:quan_width*2]; L_1176 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1176}: begin L_1177 <= data_in[quan_width-1:0]; L_1178 <= data_in[quan_width*2-1:quan_width]; L_1179 <= data_in[quan_width*3-1:quan_width*2]; L_1180 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1180}: begin L_1181 <= data_in[quan_width-1:0]; L_1182 <= data_in[quan_width*2-1:quan_width]; L_1183 <= data_in[quan_width*3-1:quan_width*2]; L_1184 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1184}: begin L_1185 <= data_in[quan_width-1:0]; L_1186 <= data_in[quan_width*2-1:quan_width]; L_1187 <= data_in[quan_width*3-1:quan_width*2]; L_1188 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1188}: begin L_1189 <= data_in[quan_width-1:0]; L_1190 <= data_in[quan_width*2-1:quan_width]; L_1191 <= data_in[quan_width*3-1:quan_width*2]; L_1192 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1192}: begin L_1193 <= data_in[quan_width-1:0]; L_1194 <= data_in[quan_width*2-1:quan_width]; L_1195 <= data_in[quan_width*3-1:quan_width*2]; L_1196 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1196}: begin L_1197 <= data_in[quan_width-1:0]; L_1198 <= data_in[quan_width*2-1:quan_width]; L_1199 <= data_in[quan_width*3-1:quan_width*2]; L_1200 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1200}: begin L_1201 <= data_in[quan_width-1:0]; L_1202 <= data_in[quan_width*2-1:quan_width]; L_1203 <= data_in[quan_width*3-1:quan_width*2]; L_1204 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1204}: begin L_1205 <= data_in[quan_width-1:0]; L_1206 <= data_in[quan_width*2-1:quan_width]; L_1207 <= data_in[quan_width*3-1:quan_width*2]; L_1208 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1208}: begin L_1209 <= data_in[quan_width-1:0]; L_1210 <= data_in[quan_width*2-1:quan_width]; L_1211 <= data_in[quan_width*3-1:quan_width*2]; L_1212 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1212}: begin L_1213 <= data_in[quan_width-1:0]; L_1214 <= data_in[quan_width*2-1:quan_width]; L_1215 <= data_in[quan_width*3-1:quan_width*2]; L_1216 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1216}: begin L_1217 <= data_in[quan_width-1:0]; L_1218 <= data_in[quan_width*2-1:quan_width]; L_1219 <= data_in[quan_width*3-1:quan_width*2]; L_1220 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1220}: begin L_1221 <= data_in[quan_width-1:0]; L_1222 <= data_in[quan_width*2-1:quan_width]; L_1223 <= data_in[quan_width*3-1:quan_width*2]; L_1224 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1224}: begin L_1225 <= data_in[quan_width-1:0]; L_1226 <= data_in[quan_width*2-1:quan_width]; L_1227 <= data_in[quan_width*3-1:quan_width*2]; L_1228 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1228}: begin L_1229 <= data_in[quan_width-1:0]; L_1230 <= data_in[quan_width*2-1:quan_width]; L_1231 <= data_in[quan_width*3-1:quan_width*2]; L_1232 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1232}: begin L_1233 <= data_in[quan_width-1:0]; L_1234 <= data_in[quan_width*2-1:quan_width]; L_1235 <= data_in[quan_width*3-1:quan_width*2]; L_1236 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1236}: begin L_1237 <= data_in[quan_width-1:0]; L_1238 <= data_in[quan_width*2-1:quan_width]; L_1239 <= data_in[quan_width*3-1:quan_width*2]; L_1240 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1240}: begin L_1241 <= data_in[quan_width-1:0]; L_1242 <= data_in[quan_width*2-1:quan_width]; L_1243 <= data_in[quan_width*3-1:quan_width*2]; L_1244 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1244}: begin L_1245 <= data_in[quan_width-1:0]; L_1246 <= data_in[quan_width*2-1:quan_width]; L_1247 <= data_in[quan_width*3-1:quan_width*2]; L_1248 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1248}: begin L_1249 <= data_in[quan_width-1:0]; L_1250 <= data_in[quan_width*2-1:quan_width]; L_1251 <= data_in[quan_width*3-1:quan_width*2]; L_1252 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1252}: begin L_1253 <= data_in[quan_width-1:0]; L_1254 <= data_in[quan_width*2-1:quan_width]; L_1255 <= data_in[quan_width*3-1:quan_width*2]; L_1256 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1256}: begin L_1257 <= data_in[quan_width-1:0]; L_1258 <= data_in[quan_width*2-1:quan_width]; L_1259 <= data_in[quan_width*3-1:quan_width*2]; L_1260 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1260}: begin L_1261 <= data_in[quan_width-1:0]; L_1262 <= data_in[quan_width*2-1:quan_width]; L_1263 <= data_in[quan_width*3-1:quan_width*2]; L_1264 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1264}: begin L_1265 <= data_in[quan_width-1:0]; L_1266 <= data_in[quan_width*2-1:quan_width]; L_1267 <= data_in[quan_width*3-1:quan_width*2]; L_1268 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1268}: begin L_1269 <= data_in[quan_width-1:0]; L_1270 <= data_in[quan_width*2-1:quan_width]; L_1271 <= data_in[quan_width*3-1:quan_width*2]; L_1272 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1272}: begin L_1273 <= data_in[quan_width-1:0]; L_1274 <= data_in[quan_width*2-1:quan_width]; L_1275 <= data_in[quan_width*3-1:quan_width*2]; L_1276 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1276}: begin L_1277 <= data_in[quan_width-1:0]; L_1278 <= data_in[quan_width*2-1:quan_width]; L_1279 <= data_in[quan_width*3-1:quan_width*2]; L_1280 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1280}: begin L_1281 <= data_in[quan_width-1:0]; L_1282 <= data_in[quan_width*2-1:quan_width]; L_1283 <= data_in[quan_width*3-1:quan_width*2]; L_1284 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1284}: begin L_1285 <= data_in[quan_width-1:0]; L_1286 <= data_in[quan_width*2-1:quan_width]; L_1287 <= data_in[quan_width*3-1:quan_width*2]; L_1288 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1288}: begin L_1289 <= data_in[quan_width-1:0]; L_1290 <= data_in[quan_width*2-1:quan_width]; L_1291 <= data_in[quan_width*3-1:quan_width*2]; L_1292 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1292}: begin L_1293 <= data_in[quan_width-1:0]; L_1294 <= data_in[quan_width*2-1:quan_width]; L_1295 <= data_in[quan_width*3-1:quan_width*2]; L_1296 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1296}: begin L_1297 <= data_in[quan_width-1:0]; L_1298 <= data_in[quan_width*2-1:quan_width]; L_1299 <= data_in[quan_width*3-1:quan_width*2]; L_1300 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1300}: begin L_1301 <= data_in[quan_width-1:0]; L_1302 <= data_in[quan_width*2-1:quan_width]; L_1303 <= data_in[quan_width*3-1:quan_width*2]; L_1304 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1304}: begin L_1305 <= data_in[quan_width-1:0]; L_1306 <= data_in[quan_width*2-1:quan_width]; L_1307 <= data_in[quan_width*3-1:quan_width*2]; L_1308 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1308}: begin L_1309 <= data_in[quan_width-1:0]; L_1310 <= data_in[quan_width*2-1:quan_width]; L_1311 <= data_in[quan_width*3-1:quan_width*2]; L_1312 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1312}: begin L_1313 <= data_in[quan_width-1:0]; L_1314 <= data_in[quan_width*2-1:quan_width]; L_1315 <= data_in[quan_width*3-1:quan_width*2]; L_1316 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1316}: begin L_1317 <= data_in[quan_width-1:0]; L_1318 <= data_in[quan_width*2-1:quan_width]; L_1319 <= data_in[quan_width*3-1:quan_width*2]; L_1320 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1320}: begin L_1321 <= data_in[quan_width-1:0]; L_1322 <= data_in[quan_width*2-1:quan_width]; L_1323 <= data_in[quan_width*3-1:quan_width*2]; L_1324 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1324}: begin L_1325 <= data_in[quan_width-1:0]; L_1326 <= data_in[quan_width*2-1:quan_width]; L_1327 <= data_in[quan_width*3-1:quan_width*2]; L_1328 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1328}: begin L_1329 <= data_in[quan_width-1:0]; L_1330 <= data_in[quan_width*2-1:quan_width]; L_1331 <= data_in[quan_width*3-1:quan_width*2]; L_1332 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1332}: begin L_1333 <= data_in[quan_width-1:0]; L_1334 <= data_in[quan_width*2-1:quan_width]; L_1335 <= data_in[quan_width*3-1:quan_width*2]; L_1336 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1336}: begin L_1337 <= data_in[quan_width-1:0]; L_1338 <= data_in[quan_width*2-1:quan_width]; L_1339 <= data_in[quan_width*3-1:quan_width*2]; L_1340 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1340}: begin L_1341 <= data_in[quan_width-1:0]; L_1342 <= data_in[quan_width*2-1:quan_width]; L_1343 <= data_in[quan_width*3-1:quan_width*2]; L_1344 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1344}: begin L_1345 <= data_in[quan_width-1:0]; L_1346 <= data_in[quan_width*2-1:quan_width]; L_1347 <= data_in[quan_width*3-1:quan_width*2]; L_1348 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1348}: begin L_1349 <= data_in[quan_width-1:0]; L_1350 <= data_in[quan_width*2-1:quan_width]; L_1351 <= data_in[quan_width*3-1:quan_width*2]; L_1352 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1352}: begin L_1353 <= data_in[quan_width-1:0]; L_1354 <= data_in[quan_width*2-1:quan_width]; L_1355 <= data_in[quan_width*3-1:quan_width*2]; L_1356 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1356}: begin L_1357 <= data_in[quan_width-1:0]; L_1358 <= data_in[quan_width*2-1:quan_width]; L_1359 <= data_in[quan_width*3-1:quan_width*2]; L_1360 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1360}: begin L_1361 <= data_in[quan_width-1:0]; L_1362 <= data_in[quan_width*2-1:quan_width]; L_1363 <= data_in[quan_width*3-1:quan_width*2]; L_1364 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1364}: begin L_1365 <= data_in[quan_width-1:0]; L_1366 <= data_in[quan_width*2-1:quan_width]; L_1367 <= data_in[quan_width*3-1:quan_width*2]; L_1368 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1368}: begin L_1369 <= data_in[quan_width-1:0]; L_1370 <= data_in[quan_width*2-1:quan_width]; L_1371 <= data_in[quan_width*3-1:quan_width*2]; L_1372 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1372}: begin L_1373 <= data_in[quan_width-1:0]; L_1374 <= data_in[quan_width*2-1:quan_width]; L_1375 <= data_in[quan_width*3-1:quan_width*2]; L_1376 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1376}: begin L_1377 <= data_in[quan_width-1:0]; L_1378 <= data_in[quan_width*2-1:quan_width]; L_1379 <= data_in[quan_width*3-1:quan_width*2]; L_1380 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1380}: begin L_1381 <= data_in[quan_width-1:0]; L_1382 <= data_in[quan_width*2-1:quan_width]; L_1383 <= data_in[quan_width*3-1:quan_width*2]; L_1384 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1384}: begin L_1385 <= data_in[quan_width-1:0]; L_1386 <= data_in[quan_width*2-1:quan_width]; L_1387 <= data_in[quan_width*3-1:quan_width*2]; L_1388 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1388}: begin L_1389 <= data_in[quan_width-1:0]; L_1390 <= data_in[quan_width*2-1:quan_width]; L_1391 <= data_in[quan_width*3-1:quan_width*2]; L_1392 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1392}: begin L_1393 <= data_in[quan_width-1:0]; L_1394 <= data_in[quan_width*2-1:quan_width]; L_1395 <= data_in[quan_width*3-1:quan_width*2]; L_1396 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1396}: begin L_1397 <= data_in[quan_width-1:0]; L_1398 <= data_in[quan_width*2-1:quan_width]; L_1399 <= data_in[quan_width*3-1:quan_width*2]; L_1400 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1400}: begin L_1401 <= data_in[quan_width-1:0]; L_1402 <= data_in[quan_width*2-1:quan_width]; L_1403 <= data_in[quan_width*3-1:quan_width*2]; L_1404 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1404}: begin L_1405 <= data_in[quan_width-1:0]; L_1406 <= data_in[quan_width*2-1:quan_width]; L_1407 <= data_in[quan_width*3-1:quan_width*2]; L_1408 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1408}: begin L_1409 <= data_in[quan_width-1:0]; L_1410 <= data_in[quan_width*2-1:quan_width]; L_1411 <= data_in[quan_width*3-1:quan_width*2]; L_1412 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1412}: begin L_1413 <= data_in[quan_width-1:0]; L_1414 <= data_in[quan_width*2-1:quan_width]; L_1415 <= data_in[quan_width*3-1:quan_width*2]; L_1416 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1416}: begin L_1417 <= data_in[quan_width-1:0]; L_1418 <= data_in[quan_width*2-1:quan_width]; L_1419 <= data_in[quan_width*3-1:quan_width*2]; L_1420 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1420}: begin L_1421 <= data_in[quan_width-1:0]; L_1422 <= data_in[quan_width*2-1:quan_width]; L_1423 <= data_in[quan_width*3-1:quan_width*2]; L_1424 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1424}: begin L_1425 <= data_in[quan_width-1:0]; L_1426 <= data_in[quan_width*2-1:quan_width]; L_1427 <= data_in[quan_width*3-1:quan_width*2]; L_1428 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1428}: begin L_1429 <= data_in[quan_width-1:0]; L_1430 <= data_in[quan_width*2-1:quan_width]; L_1431 <= data_in[quan_width*3-1:quan_width*2]; L_1432 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1432}: begin L_1433 <= data_in[quan_width-1:0]; L_1434 <= data_in[quan_width*2-1:quan_width]; L_1435 <= data_in[quan_width*3-1:quan_width*2]; L_1436 <= data_in[quan_width*4-1:quan_width*3]; end
		{1'b1, 16'd1436}: begin L_1437 <= data_in[quan_width-1:0]; L_1438 <= data_in[quan_width*2-1:quan_width]; L_1439 <= data_in[quan_width*3-1:quan_width*2]; L_1440 <= data_in[quan_width*4-1:quan_width*3]; end
	endcase
end

always @ (posedge clk) begin
if (in_valid == 0 && cnt == 0)
cnt <= 1;
end

always @ (posedge clk) begin
	case ({out_valid, out_index})
		{1'b1, 16'd0}: begin data_out[0] <= Bit_1; data_out[1] <= Bit_2;data_out[2] <= Bit_3; data_out[3] <= Bit_4; end
		{1'b1, 16'd4}: begin data_out[0] <= Bit_5; data_out[1] <= Bit_6;data_out[2] <= Bit_7; data_out[3] <= Bit_8; end
		{1'b1, 16'd8}: begin data_out[0] <= Bit_9; data_out[1] <= Bit_10;data_out[2] <= Bit_11; data_out[3] <= Bit_12; end
		{1'b1, 16'd12}: begin data_out[0] <= Bit_13; data_out[1] <= Bit_14;data_out[2] <= Bit_15; data_out[3] <= Bit_16; end
		{1'b1, 16'd16}: begin data_out[0] <= Bit_17; data_out[1] <= Bit_18;data_out[2] <= Bit_19; data_out[3] <= Bit_20; end
		{1'b1, 16'd20}: begin data_out[0] <= Bit_21; data_out[1] <= Bit_22;data_out[2] <= Bit_23; data_out[3] <= Bit_24; end
		{1'b1, 16'd24}: begin data_out[0] <= Bit_25; data_out[1] <= Bit_26;data_out[2] <= Bit_27; data_out[3] <= Bit_28; end
		{1'b1, 16'd28}: begin data_out[0] <= Bit_29; data_out[1] <= Bit_30;data_out[2] <= Bit_31; data_out[3] <= Bit_32; end
		{1'b1, 16'd32}: begin data_out[0] <= Bit_33; data_out[1] <= Bit_34;data_out[2] <= Bit_35; data_out[3] <= Bit_36; end
		{1'b1, 16'd36}: begin data_out[0] <= Bit_37; data_out[1] <= Bit_38;data_out[2] <= Bit_39; data_out[3] <= Bit_40; end
		{1'b1, 16'd40}: begin data_out[0] <= Bit_41; data_out[1] <= Bit_42;data_out[2] <= Bit_43; data_out[3] <= Bit_44; end
		{1'b1, 16'd44}: begin data_out[0] <= Bit_45; data_out[1] <= Bit_46;data_out[2] <= Bit_47; data_out[3] <= Bit_48; end
		{1'b1, 16'd48}: begin data_out[0] <= Bit_49; data_out[1] <= Bit_50;data_out[2] <= Bit_51; data_out[3] <= Bit_52; end
		{1'b1, 16'd52}: begin data_out[0] <= Bit_53; data_out[1] <= Bit_54;data_out[2] <= Bit_55; data_out[3] <= Bit_56; end
		{1'b1, 16'd56}: begin data_out[0] <= Bit_57; data_out[1] <= Bit_58;data_out[2] <= Bit_59; data_out[3] <= Bit_60; end
		{1'b1, 16'd60}: begin data_out[0] <= Bit_61; data_out[1] <= Bit_62;data_out[2] <= Bit_63; data_out[3] <= Bit_64; end
		{1'b1, 16'd64}: begin data_out[0] <= Bit_65; data_out[1] <= Bit_66;data_out[2] <= Bit_67; data_out[3] <= Bit_68; end
		{1'b1, 16'd68}: begin data_out[0] <= Bit_69; data_out[1] <= Bit_70;data_out[2] <= Bit_71; data_out[3] <= Bit_72; end
		{1'b1, 16'd72}: begin data_out[0] <= Bit_73; data_out[1] <= Bit_74;data_out[2] <= Bit_75; data_out[3] <= Bit_76; end
		{1'b1, 16'd76}: begin data_out[0] <= Bit_77; data_out[1] <= Bit_78;data_out[2] <= Bit_79; data_out[3] <= Bit_80; end
		{1'b1, 16'd80}: begin data_out[0] <= Bit_81; data_out[1] <= Bit_82;data_out[2] <= Bit_83; data_out[3] <= Bit_84; end
		{1'b1, 16'd84}: begin data_out[0] <= Bit_85; data_out[1] <= Bit_86;data_out[2] <= Bit_87; data_out[3] <= Bit_88; end
		{1'b1, 16'd88}: begin data_out[0] <= Bit_89; data_out[1] <= Bit_90;data_out[2] <= Bit_91; data_out[3] <= Bit_92; end
		{1'b1, 16'd92}: begin data_out[0] <= Bit_93; data_out[1] <= Bit_94;data_out[2] <= Bit_95; data_out[3] <= Bit_96; end
		{1'b1, 16'd96}: begin data_out[0] <= Bit_97; data_out[1] <= Bit_98;data_out[2] <= Bit_99; data_out[3] <= Bit_100; end
		{1'b1, 16'd100}: begin data_out[0] <= Bit_101; data_out[1] <= Bit_102;data_out[2] <= Bit_103; data_out[3] <= Bit_104; end
		{1'b1, 16'd104}: begin data_out[0] <= Bit_105; data_out[1] <= Bit_106;data_out[2] <= Bit_107; data_out[3] <= Bit_108; end
		{1'b1, 16'd108}: begin data_out[0] <= Bit_109; data_out[1] <= Bit_110;data_out[2] <= Bit_111; data_out[3] <= Bit_112; end
		{1'b1, 16'd112}: begin data_out[0] <= Bit_113; data_out[1] <= Bit_114;data_out[2] <= Bit_115; data_out[3] <= Bit_116; end
		{1'b1, 16'd116}: begin data_out[0] <= Bit_117; data_out[1] <= Bit_118;data_out[2] <= Bit_119; data_out[3] <= Bit_120; end
		{1'b1, 16'd120}: begin data_out[0] <= Bit_121; data_out[1] <= Bit_122;data_out[2] <= Bit_123; data_out[3] <= Bit_124; end
		{1'b1, 16'd124}: begin data_out[0] <= Bit_125; data_out[1] <= Bit_126;data_out[2] <= Bit_127; data_out[3] <= Bit_128; end
		{1'b1, 16'd128}: begin data_out[0] <= Bit_129; data_out[1] <= Bit_130;data_out[2] <= Bit_131; data_out[3] <= Bit_132; end
		{1'b1, 16'd132}: begin data_out[0] <= Bit_133; data_out[1] <= Bit_134;data_out[2] <= Bit_135; data_out[3] <= Bit_136; end
		{1'b1, 16'd136}: begin data_out[0] <= Bit_137; data_out[1] <= Bit_138;data_out[2] <= Bit_139; data_out[3] <= Bit_140; end
		{1'b1, 16'd140}: begin data_out[0] <= Bit_141; data_out[1] <= Bit_142;data_out[2] <= Bit_143; data_out[3] <= Bit_144; end
		{1'b1, 16'd144}: begin data_out[0] <= Bit_145; data_out[1] <= Bit_146;data_out[2] <= Bit_147; data_out[3] <= Bit_148; end
		{1'b1, 16'd148}: begin data_out[0] <= Bit_149; data_out[1] <= Bit_150;data_out[2] <= Bit_151; data_out[3] <= Bit_152; end
		{1'b1, 16'd152}: begin data_out[0] <= Bit_153; data_out[1] <= Bit_154;data_out[2] <= Bit_155; data_out[3] <= Bit_156; end
		{1'b1, 16'd156}: begin data_out[0] <= Bit_157; data_out[1] <= Bit_158;data_out[2] <= Bit_159; data_out[3] <= Bit_160; end
		{1'b1, 16'd160}: begin data_out[0] <= Bit_161; data_out[1] <= Bit_162;data_out[2] <= Bit_163; data_out[3] <= Bit_164; end
		{1'b1, 16'd164}: begin data_out[0] <= Bit_165; data_out[1] <= Bit_166;data_out[2] <= Bit_167; data_out[3] <= Bit_168; end
		{1'b1, 16'd168}: begin data_out[0] <= Bit_169; data_out[1] <= Bit_170;data_out[2] <= Bit_171; data_out[3] <= Bit_172; end
		{1'b1, 16'd172}: begin data_out[0] <= Bit_173; data_out[1] <= Bit_174;data_out[2] <= Bit_175; data_out[3] <= Bit_176; end
		{1'b1, 16'd176}: begin data_out[0] <= Bit_177; data_out[1] <= Bit_178;data_out[2] <= Bit_179; data_out[3] <= Bit_180; end
		{1'b1, 16'd180}: begin data_out[0] <= Bit_181; data_out[1] <= Bit_182;data_out[2] <= Bit_183; data_out[3] <= Bit_184; end
		{1'b1, 16'd184}: begin data_out[0] <= Bit_185; data_out[1] <= Bit_186;data_out[2] <= Bit_187; data_out[3] <= Bit_188; end
		{1'b1, 16'd188}: begin data_out[0] <= Bit_189; data_out[1] <= Bit_190;data_out[2] <= Bit_191; data_out[3] <= Bit_192; end
		{1'b1, 16'd192}: begin data_out[0] <= Bit_193; data_out[1] <= Bit_194;data_out[2] <= Bit_195; data_out[3] <= Bit_196; end
		{1'b1, 16'd196}: begin data_out[0] <= Bit_197; data_out[1] <= Bit_198;data_out[2] <= Bit_199; data_out[3] <= Bit_200; end
		{1'b1, 16'd200}: begin data_out[0] <= Bit_201; data_out[1] <= Bit_202;data_out[2] <= Bit_203; data_out[3] <= Bit_204; end
		{1'b1, 16'd204}: begin data_out[0] <= Bit_205; data_out[1] <= Bit_206;data_out[2] <= Bit_207; data_out[3] <= Bit_208; end
		{1'b1, 16'd208}: begin data_out[0] <= Bit_209; data_out[1] <= Bit_210;data_out[2] <= Bit_211; data_out[3] <= Bit_212; end
		{1'b1, 16'd212}: begin data_out[0] <= Bit_213; data_out[1] <= Bit_214;data_out[2] <= Bit_215; data_out[3] <= Bit_216; end
		{1'b1, 16'd216}: begin data_out[0] <= Bit_217; data_out[1] <= Bit_218;data_out[2] <= Bit_219; data_out[3] <= Bit_220; end
		{1'b1, 16'd220}: begin data_out[0] <= Bit_221; data_out[1] <= Bit_222;data_out[2] <= Bit_223; data_out[3] <= Bit_224; end
		{1'b1, 16'd224}: begin data_out[0] <= Bit_225; data_out[1] <= Bit_226;data_out[2] <= Bit_227; data_out[3] <= Bit_228; end
		{1'b1, 16'd228}: begin data_out[0] <= Bit_229; data_out[1] <= Bit_230;data_out[2] <= Bit_231; data_out[3] <= Bit_232; end
		{1'b1, 16'd232}: begin data_out[0] <= Bit_233; data_out[1] <= Bit_234;data_out[2] <= Bit_235; data_out[3] <= Bit_236; end
		{1'b1, 16'd236}: begin data_out[0] <= Bit_237; data_out[1] <= Bit_238;data_out[2] <= Bit_239; data_out[3] <= Bit_240; end
		{1'b1, 16'd240}: begin data_out[0] <= Bit_241; data_out[1] <= Bit_242;data_out[2] <= Bit_243; data_out[3] <= Bit_244; end
		{1'b1, 16'd244}: begin data_out[0] <= Bit_245; data_out[1] <= Bit_246;data_out[2] <= Bit_247; data_out[3] <= Bit_248; end
		{1'b1, 16'd248}: begin data_out[0] <= Bit_249; data_out[1] <= Bit_250;data_out[2] <= Bit_251; data_out[3] <= Bit_252; end
		{1'b1, 16'd252}: begin data_out[0] <= Bit_253; data_out[1] <= Bit_254;data_out[2] <= Bit_255; data_out[3] <= Bit_256; end
		{1'b1, 16'd256}: begin data_out[0] <= Bit_257; data_out[1] <= Bit_258;data_out[2] <= Bit_259; data_out[3] <= Bit_260; end
		{1'b1, 16'd260}: begin data_out[0] <= Bit_261; data_out[1] <= Bit_262;data_out[2] <= Bit_263; data_out[3] <= Bit_264; end
		{1'b1, 16'd264}: begin data_out[0] <= Bit_265; data_out[1] <= Bit_266;data_out[2] <= Bit_267; data_out[3] <= Bit_268; end
		{1'b1, 16'd268}: begin data_out[0] <= Bit_269; data_out[1] <= Bit_270;data_out[2] <= Bit_271; data_out[3] <= Bit_272; end
		{1'b1, 16'd272}: begin data_out[0] <= Bit_273; data_out[1] <= Bit_274;data_out[2] <= Bit_275; data_out[3] <= Bit_276; end
		{1'b1, 16'd276}: begin data_out[0] <= Bit_277; data_out[1] <= Bit_278;data_out[2] <= Bit_279; data_out[3] <= Bit_280; end
		{1'b1, 16'd280}: begin data_out[0] <= Bit_281; data_out[1] <= Bit_282;data_out[2] <= Bit_283; data_out[3] <= Bit_284; end
		{1'b1, 16'd284}: begin data_out[0] <= Bit_285; data_out[1] <= Bit_286;data_out[2] <= Bit_287; data_out[3] <= Bit_288; end
		{1'b1, 16'd288}: begin data_out[0] <= Bit_289; data_out[1] <= Bit_290;data_out[2] <= Bit_291; data_out[3] <= Bit_292; end
		{1'b1, 16'd292}: begin data_out[0] <= Bit_293; data_out[1] <= Bit_294;data_out[2] <= Bit_295; data_out[3] <= Bit_296; end
		{1'b1, 16'd296}: begin data_out[0] <= Bit_297; data_out[1] <= Bit_298;data_out[2] <= Bit_299; data_out[3] <= Bit_300; end
		{1'b1, 16'd300}: begin data_out[0] <= Bit_301; data_out[1] <= Bit_302;data_out[2] <= Bit_303; data_out[3] <= Bit_304; end
		{1'b1, 16'd304}: begin data_out[0] <= Bit_305; data_out[1] <= Bit_306;data_out[2] <= Bit_307; data_out[3] <= Bit_308; end
		{1'b1, 16'd308}: begin data_out[0] <= Bit_309; data_out[1] <= Bit_310;data_out[2] <= Bit_311; data_out[3] <= Bit_312; end
		{1'b1, 16'd312}: begin data_out[0] <= Bit_313; data_out[1] <= Bit_314;data_out[2] <= Bit_315; data_out[3] <= Bit_316; end
		{1'b1, 16'd316}: begin data_out[0] <= Bit_317; data_out[1] <= Bit_318;data_out[2] <= Bit_319; data_out[3] <= Bit_320; end
		{1'b1, 16'd320}: begin data_out[0] <= Bit_321; data_out[1] <= Bit_322;data_out[2] <= Bit_323; data_out[3] <= Bit_324; end
		{1'b1, 16'd324}: begin data_out[0] <= Bit_325; data_out[1] <= Bit_326;data_out[2] <= Bit_327; data_out[3] <= Bit_328; end
		{1'b1, 16'd328}: begin data_out[0] <= Bit_329; data_out[1] <= Bit_330;data_out[2] <= Bit_331; data_out[3] <= Bit_332; end
		{1'b1, 16'd332}: begin data_out[0] <= Bit_333; data_out[1] <= Bit_334;data_out[2] <= Bit_335; data_out[3] <= Bit_336; end
		{1'b1, 16'd336}: begin data_out[0] <= Bit_337; data_out[1] <= Bit_338;data_out[2] <= Bit_339; data_out[3] <= Bit_340; end
		{1'b1, 16'd340}: begin data_out[0] <= Bit_341; data_out[1] <= Bit_342;data_out[2] <= Bit_343; data_out[3] <= Bit_344; end
		{1'b1, 16'd344}: begin data_out[0] <= Bit_345; data_out[1] <= Bit_346;data_out[2] <= Bit_347; data_out[3] <= Bit_348; end
		{1'b1, 16'd348}: begin data_out[0] <= Bit_349; data_out[1] <= Bit_350;data_out[2] <= Bit_351; data_out[3] <= Bit_352; end
		{1'b1, 16'd352}: begin data_out[0] <= Bit_353; data_out[1] <= Bit_354;data_out[2] <= Bit_355; data_out[3] <= Bit_356; end
		{1'b1, 16'd356}: begin data_out[0] <= Bit_357; data_out[1] <= Bit_358;data_out[2] <= Bit_359; data_out[3] <= Bit_360; end
		{1'b1, 16'd360}: begin data_out[0] <= Bit_361; data_out[1] <= Bit_362;data_out[2] <= Bit_363; data_out[3] <= Bit_364; end
		{1'b1, 16'd364}: begin data_out[0] <= Bit_365; data_out[1] <= Bit_366;data_out[2] <= Bit_367; data_out[3] <= Bit_368; end
		{1'b1, 16'd368}: begin data_out[0] <= Bit_369; data_out[1] <= Bit_370;data_out[2] <= Bit_371; data_out[3] <= Bit_372; end
		{1'b1, 16'd372}: begin data_out[0] <= Bit_373; data_out[1] <= Bit_374;data_out[2] <= Bit_375; data_out[3] <= Bit_376; end
		{1'b1, 16'd376}: begin data_out[0] <= Bit_377; data_out[1] <= Bit_378;data_out[2] <= Bit_379; data_out[3] <= Bit_380; end
		{1'b1, 16'd380}: begin data_out[0] <= Bit_381; data_out[1] <= Bit_382;data_out[2] <= Bit_383; data_out[3] <= Bit_384; end
		{1'b1, 16'd384}: begin data_out[0] <= Bit_385; data_out[1] <= Bit_386;data_out[2] <= Bit_387; data_out[3] <= Bit_388; end
		{1'b1, 16'd388}: begin data_out[0] <= Bit_389; data_out[1] <= Bit_390;data_out[2] <= Bit_391; data_out[3] <= Bit_392; end
		{1'b1, 16'd392}: begin data_out[0] <= Bit_393; data_out[1] <= Bit_394;data_out[2] <= Bit_395; data_out[3] <= Bit_396; end
		{1'b1, 16'd396}: begin data_out[0] <= Bit_397; data_out[1] <= Bit_398;data_out[2] <= Bit_399; data_out[3] <= Bit_400; end
		{1'b1, 16'd400}: begin data_out[0] <= Bit_401; data_out[1] <= Bit_402;data_out[2] <= Bit_403; data_out[3] <= Bit_404; end
		{1'b1, 16'd404}: begin data_out[0] <= Bit_405; data_out[1] <= Bit_406;data_out[2] <= Bit_407; data_out[3] <= Bit_408; end
		{1'b1, 16'd408}: begin data_out[0] <= Bit_409; data_out[1] <= Bit_410;data_out[2] <= Bit_411; data_out[3] <= Bit_412; end
		{1'b1, 16'd412}: begin data_out[0] <= Bit_413; data_out[1] <= Bit_414;data_out[2] <= Bit_415; data_out[3] <= Bit_416; end
		{1'b1, 16'd416}: begin data_out[0] <= Bit_417; data_out[1] <= Bit_418;data_out[2] <= Bit_419; data_out[3] <= Bit_420; end
		{1'b1, 16'd420}: begin data_out[0] <= Bit_421; data_out[1] <= Bit_422;data_out[2] <= Bit_423; data_out[3] <= Bit_424; end
		{1'b1, 16'd424}: begin data_out[0] <= Bit_425; data_out[1] <= Bit_426;data_out[2] <= Bit_427; data_out[3] <= Bit_428; end
		{1'b1, 16'd428}: begin data_out[0] <= Bit_429; data_out[1] <= Bit_430;data_out[2] <= Bit_431; data_out[3] <= Bit_432; end
		{1'b1, 16'd432}: begin data_out[0] <= Bit_433; data_out[1] <= Bit_434;data_out[2] <= Bit_435; data_out[3] <= Bit_436; end
		{1'b1, 16'd436}: begin data_out[0] <= Bit_437; data_out[1] <= Bit_438;data_out[2] <= Bit_439; data_out[3] <= Bit_440; end
		{1'b1, 16'd440}: begin data_out[0] <= Bit_441; data_out[1] <= Bit_442;data_out[2] <= Bit_443; data_out[3] <= Bit_444; end
		{1'b1, 16'd444}: begin data_out[0] <= Bit_445; data_out[1] <= Bit_446;data_out[2] <= Bit_447; data_out[3] <= Bit_448; end
		{1'b1, 16'd448}: begin data_out[0] <= Bit_449; data_out[1] <= Bit_450;data_out[2] <= Bit_451; data_out[3] <= Bit_452; end
		{1'b1, 16'd452}: begin data_out[0] <= Bit_453; data_out[1] <= Bit_454;data_out[2] <= Bit_455; data_out[3] <= Bit_456; end
		{1'b1, 16'd456}: begin data_out[0] <= Bit_457; data_out[1] <= Bit_458;data_out[2] <= Bit_459; data_out[3] <= Bit_460; end
		{1'b1, 16'd460}: begin data_out[0] <= Bit_461; data_out[1] <= Bit_462;data_out[2] <= Bit_463; data_out[3] <= Bit_464; end
		{1'b1, 16'd464}: begin data_out[0] <= Bit_465; data_out[1] <= Bit_466;data_out[2] <= Bit_467; data_out[3] <= Bit_468; end
		{1'b1, 16'd468}: begin data_out[0] <= Bit_469; data_out[1] <= Bit_470;data_out[2] <= Bit_471; data_out[3] <= Bit_472; end
		{1'b1, 16'd472}: begin data_out[0] <= Bit_473; data_out[1] <= Bit_474;data_out[2] <= Bit_475; data_out[3] <= Bit_476; end
		{1'b1, 16'd476}: begin data_out[0] <= Bit_477; data_out[1] <= Bit_478;data_out[2] <= Bit_479; data_out[3] <= Bit_480; end
		{1'b1, 16'd480}: begin data_out[0] <= Bit_481; data_out[1] <= Bit_482;data_out[2] <= Bit_483; data_out[3] <= Bit_484; end
		{1'b1, 16'd484}: begin data_out[0] <= Bit_485; data_out[1] <= Bit_486;data_out[2] <= Bit_487; data_out[3] <= Bit_488; end
		{1'b1, 16'd488}: begin data_out[0] <= Bit_489; data_out[1] <= Bit_490;data_out[2] <= Bit_491; data_out[3] <= Bit_492; end
		{1'b1, 16'd492}: begin data_out[0] <= Bit_493; data_out[1] <= Bit_494;data_out[2] <= Bit_495; data_out[3] <= Bit_496; end
		{1'b1, 16'd496}: begin data_out[0] <= Bit_497; data_out[1] <= Bit_498;data_out[2] <= Bit_499; data_out[3] <= Bit_500; end
		{1'b1, 16'd500}: begin data_out[0] <= Bit_501; data_out[1] <= Bit_502;data_out[2] <= Bit_503; data_out[3] <= Bit_504; end
		{1'b1, 16'd504}: begin data_out[0] <= Bit_505; data_out[1] <= Bit_506;data_out[2] <= Bit_507; data_out[3] <= Bit_508; end
		{1'b1, 16'd508}: begin data_out[0] <= Bit_509; data_out[1] <= Bit_510;data_out[2] <= Bit_511; data_out[3] <= Bit_512; end
		{1'b1, 16'd512}: begin data_out[0] <= Bit_513; data_out[1] <= Bit_514;data_out[2] <= Bit_515; data_out[3] <= Bit_516; end
		{1'b1, 16'd516}: begin data_out[0] <= Bit_517; data_out[1] <= Bit_518;data_out[2] <= Bit_519; data_out[3] <= Bit_520; end
		{1'b1, 16'd520}: begin data_out[0] <= Bit_521; data_out[1] <= Bit_522;data_out[2] <= Bit_523; data_out[3] <= Bit_524; end
		{1'b1, 16'd524}: begin data_out[0] <= Bit_525; data_out[1] <= Bit_526;data_out[2] <= Bit_527; data_out[3] <= Bit_528; end
		{1'b1, 16'd528}: begin data_out[0] <= Bit_529; data_out[1] <= Bit_530;data_out[2] <= Bit_531; data_out[3] <= Bit_532; end
		{1'b1, 16'd532}: begin data_out[0] <= Bit_533; data_out[1] <= Bit_534;data_out[2] <= Bit_535; data_out[3] <= Bit_536; end
		{1'b1, 16'd536}: begin data_out[0] <= Bit_537; data_out[1] <= Bit_538;data_out[2] <= Bit_539; data_out[3] <= Bit_540; end
		{1'b1, 16'd540}: begin data_out[0] <= Bit_541; data_out[1] <= Bit_542;data_out[2] <= Bit_543; data_out[3] <= Bit_544; end
		{1'b1, 16'd544}: begin data_out[0] <= Bit_545; data_out[1] <= Bit_546;data_out[2] <= Bit_547; data_out[3] <= Bit_548; end
		{1'b1, 16'd548}: begin data_out[0] <= Bit_549; data_out[1] <= Bit_550;data_out[2] <= Bit_551; data_out[3] <= Bit_552; end
		{1'b1, 16'd552}: begin data_out[0] <= Bit_553; data_out[1] <= Bit_554;data_out[2] <= Bit_555; data_out[3] <= Bit_556; end
		{1'b1, 16'd556}: begin data_out[0] <= Bit_557; data_out[1] <= Bit_558;data_out[2] <= Bit_559; data_out[3] <= Bit_560; end
		{1'b1, 16'd560}: begin data_out[0] <= Bit_561; data_out[1] <= Bit_562;data_out[2] <= Bit_563; data_out[3] <= Bit_564; end
		{1'b1, 16'd564}: begin data_out[0] <= Bit_565; data_out[1] <= Bit_566;data_out[2] <= Bit_567; data_out[3] <= Bit_568; end
		{1'b1, 16'd568}: begin data_out[0] <= Bit_569; data_out[1] <= Bit_570;data_out[2] <= Bit_571; data_out[3] <= Bit_572; end
		{1'b1, 16'd572}: begin data_out[0] <= Bit_573; data_out[1] <= Bit_574;data_out[2] <= Bit_575; data_out[3] <= Bit_576; end
		{1'b1, 16'd576}: begin data_out[0] <= Bit_577; data_out[1] <= Bit_578;data_out[2] <= Bit_579; data_out[3] <= Bit_580; end
		{1'b1, 16'd580}: begin data_out[0] <= Bit_581; data_out[1] <= Bit_582;data_out[2] <= Bit_583; data_out[3] <= Bit_584; end
		{1'b1, 16'd584}: begin data_out[0] <= Bit_585; data_out[1] <= Bit_586;data_out[2] <= Bit_587; data_out[3] <= Bit_588; end
		{1'b1, 16'd588}: begin data_out[0] <= Bit_589; data_out[1] <= Bit_590;data_out[2] <= Bit_591; data_out[3] <= Bit_592; end
		{1'b1, 16'd592}: begin data_out[0] <= Bit_593; data_out[1] <= Bit_594;data_out[2] <= Bit_595; data_out[3] <= Bit_596; end
		{1'b1, 16'd596}: begin data_out[0] <= Bit_597; data_out[1] <= Bit_598;data_out[2] <= Bit_599; data_out[3] <= Bit_600; end
		{1'b1, 16'd600}: begin data_out[0] <= Bit_601; data_out[1] <= Bit_602;data_out[2] <= Bit_603; data_out[3] <= Bit_604; end
		{1'b1, 16'd604}: begin data_out[0] <= Bit_605; data_out[1] <= Bit_606;data_out[2] <= Bit_607; data_out[3] <= Bit_608; end
		{1'b1, 16'd608}: begin data_out[0] <= Bit_609; data_out[1] <= Bit_610;data_out[2] <= Bit_611; data_out[3] <= Bit_612; end
		{1'b1, 16'd612}: begin data_out[0] <= Bit_613; data_out[1] <= Bit_614;data_out[2] <= Bit_615; data_out[3] <= Bit_616; end
		{1'b1, 16'd616}: begin data_out[0] <= Bit_617; data_out[1] <= Bit_618;data_out[2] <= Bit_619; data_out[3] <= Bit_620; end
		{1'b1, 16'd620}: begin data_out[0] <= Bit_621; data_out[1] <= Bit_622;data_out[2] <= Bit_623; data_out[3] <= Bit_624; end
		{1'b1, 16'd624}: begin data_out[0] <= Bit_625; data_out[1] <= Bit_626;data_out[2] <= Bit_627; data_out[3] <= Bit_628; end
		{1'b1, 16'd628}: begin data_out[0] <= Bit_629; data_out[1] <= Bit_630;data_out[2] <= Bit_631; data_out[3] <= Bit_632; end
		{1'b1, 16'd632}: begin data_out[0] <= Bit_633; data_out[1] <= Bit_634;data_out[2] <= Bit_635; data_out[3] <= Bit_636; end
		{1'b1, 16'd636}: begin data_out[0] <= Bit_637; data_out[1] <= Bit_638;data_out[2] <= Bit_639; data_out[3] <= Bit_640; end
		{1'b1, 16'd640}: begin data_out[0] <= Bit_641; data_out[1] <= Bit_642;data_out[2] <= Bit_643; data_out[3] <= Bit_644; end
		{1'b1, 16'd644}: begin data_out[0] <= Bit_645; data_out[1] <= Bit_646;data_out[2] <= Bit_647; data_out[3] <= Bit_648; end
		{1'b1, 16'd648}: begin data_out[0] <= Bit_649; data_out[1] <= Bit_650;data_out[2] <= Bit_651; data_out[3] <= Bit_652; end
		{1'b1, 16'd652}: begin data_out[0] <= Bit_653; data_out[1] <= Bit_654;data_out[2] <= Bit_655; data_out[3] <= Bit_656; end
		{1'b1, 16'd656}: begin data_out[0] <= Bit_657; data_out[1] <= Bit_658;data_out[2] <= Bit_659; data_out[3] <= Bit_660; end
		{1'b1, 16'd660}: begin data_out[0] <= Bit_661; data_out[1] <= Bit_662;data_out[2] <= Bit_663; data_out[3] <= Bit_664; end
		{1'b1, 16'd664}: begin data_out[0] <= Bit_665; data_out[1] <= Bit_666;data_out[2] <= Bit_667; data_out[3] <= Bit_668; end
		{1'b1, 16'd668}: begin data_out[0] <= Bit_669; data_out[1] <= Bit_670;data_out[2] <= Bit_671; data_out[3] <= Bit_672; end
		{1'b1, 16'd672}: begin data_out[0] <= Bit_673; data_out[1] <= Bit_674;data_out[2] <= Bit_675; data_out[3] <= Bit_676; end
		{1'b1, 16'd676}: begin data_out[0] <= Bit_677; data_out[1] <= Bit_678;data_out[2] <= Bit_679; data_out[3] <= Bit_680; end
		{1'b1, 16'd680}: begin data_out[0] <= Bit_681; data_out[1] <= Bit_682;data_out[2] <= Bit_683; data_out[3] <= Bit_684; end
		{1'b1, 16'd684}: begin data_out[0] <= Bit_685; data_out[1] <= Bit_686;data_out[2] <= Bit_687; data_out[3] <= Bit_688; end
		{1'b1, 16'd688}: begin data_out[0] <= Bit_689; data_out[1] <= Bit_690;data_out[2] <= Bit_691; data_out[3] <= Bit_692; end
		{1'b1, 16'd692}: begin data_out[0] <= Bit_693; data_out[1] <= Bit_694;data_out[2] <= Bit_695; data_out[3] <= Bit_696; end
		{1'b1, 16'd696}: begin data_out[0] <= Bit_697; data_out[1] <= Bit_698;data_out[2] <= Bit_699; data_out[3] <= Bit_700; end
		{1'b1, 16'd700}: begin data_out[0] <= Bit_701; data_out[1] <= Bit_702;data_out[2] <= Bit_703; data_out[3] <= Bit_704; end
		{1'b1, 16'd704}: begin data_out[0] <= Bit_705; data_out[1] <= Bit_706;data_out[2] <= Bit_707; data_out[3] <= Bit_708; end
		{1'b1, 16'd708}: begin data_out[0] <= Bit_709; data_out[1] <= Bit_710;data_out[2] <= Bit_711; data_out[3] <= Bit_712; end
		{1'b1, 16'd712}: begin data_out[0] <= Bit_713; data_out[1] <= Bit_714;data_out[2] <= Bit_715; data_out[3] <= Bit_716; end
		{1'b1, 16'd716}: begin data_out[0] <= Bit_717; data_out[1] <= Bit_718;data_out[2] <= Bit_719; data_out[3] <= Bit_720; end
		{1'b1, 16'd720}: begin data_out[0] <= Bit_721; data_out[1] <= Bit_722;data_out[2] <= Bit_723; data_out[3] <= Bit_724; end
		{1'b1, 16'd724}: begin data_out[0] <= Bit_725; data_out[1] <= Bit_726;data_out[2] <= Bit_727; data_out[3] <= Bit_728; end
		{1'b1, 16'd728}: begin data_out[0] <= Bit_729; data_out[1] <= Bit_730;data_out[2] <= Bit_731; data_out[3] <= Bit_732; end
		{1'b1, 16'd732}: begin data_out[0] <= Bit_733; data_out[1] <= Bit_734;data_out[2] <= Bit_735; data_out[3] <= Bit_736; end
		{1'b1, 16'd736}: begin data_out[0] <= Bit_737; data_out[1] <= Bit_738;data_out[2] <= Bit_739; data_out[3] <= Bit_740; end
		{1'b1, 16'd740}: begin data_out[0] <= Bit_741; data_out[1] <= Bit_742;data_out[2] <= Bit_743; data_out[3] <= Bit_744; end
		{1'b1, 16'd744}: begin data_out[0] <= Bit_745; data_out[1] <= Bit_746;data_out[2] <= Bit_747; data_out[3] <= Bit_748; end
		{1'b1, 16'd748}: begin data_out[0] <= Bit_749; data_out[1] <= Bit_750;data_out[2] <= Bit_751; data_out[3] <= Bit_752; end
		{1'b1, 16'd752}: begin data_out[0] <= Bit_753; data_out[1] <= Bit_754;data_out[2] <= Bit_755; data_out[3] <= Bit_756; end
		{1'b1, 16'd756}: begin data_out[0] <= Bit_757; data_out[1] <= Bit_758;data_out[2] <= Bit_759; data_out[3] <= Bit_760; end
		{1'b1, 16'd760}: begin data_out[0] <= Bit_761; data_out[1] <= Bit_762;data_out[2] <= Bit_763; data_out[3] <= Bit_764; end
		{1'b1, 16'd764}: begin data_out[0] <= Bit_765; data_out[1] <= Bit_766;data_out[2] <= Bit_767; data_out[3] <= Bit_768; end
		{1'b1, 16'd768}: begin data_out[0] <= Bit_769; data_out[1] <= Bit_770;data_out[2] <= Bit_771; data_out[3] <= Bit_772; end
		{1'b1, 16'd772}: begin data_out[0] <= Bit_773; data_out[1] <= Bit_774;data_out[2] <= Bit_775; data_out[3] <= Bit_776; end
		{1'b1, 16'd776}: begin data_out[0] <= Bit_777; data_out[1] <= Bit_778;data_out[2] <= Bit_779; data_out[3] <= Bit_780; end
		{1'b1, 16'd780}: begin data_out[0] <= Bit_781; data_out[1] <= Bit_782;data_out[2] <= Bit_783; data_out[3] <= Bit_784; end
		{1'b1, 16'd784}: begin data_out[0] <= Bit_785; data_out[1] <= Bit_786;data_out[2] <= Bit_787; data_out[3] <= Bit_788; end
		{1'b1, 16'd788}: begin data_out[0] <= Bit_789; data_out[1] <= Bit_790;data_out[2] <= Bit_791; data_out[3] <= Bit_792; end
		{1'b1, 16'd792}: begin data_out[0] <= Bit_793; data_out[1] <= Bit_794;data_out[2] <= Bit_795; data_out[3] <= Bit_796; end
		{1'b1, 16'd796}: begin data_out[0] <= Bit_797; data_out[1] <= Bit_798;data_out[2] <= Bit_799; data_out[3] <= Bit_800; end
		{1'b1, 16'd800}: begin data_out[0] <= Bit_801; data_out[1] <= Bit_802;data_out[2] <= Bit_803; data_out[3] <= Bit_804; end
		{1'b1, 16'd804}: begin data_out[0] <= Bit_805; data_out[1] <= Bit_806;data_out[2] <= Bit_807; data_out[3] <= Bit_808; end
		{1'b1, 16'd808}: begin data_out[0] <= Bit_809; data_out[1] <= Bit_810;data_out[2] <= Bit_811; data_out[3] <= Bit_812; end
		{1'b1, 16'd812}: begin data_out[0] <= Bit_813; data_out[1] <= Bit_814;data_out[2] <= Bit_815; data_out[3] <= Bit_816; end
		{1'b1, 16'd816}: begin data_out[0] <= Bit_817; data_out[1] <= Bit_818;data_out[2] <= Bit_819; data_out[3] <= Bit_820; end
		{1'b1, 16'd820}: begin data_out[0] <= Bit_821; data_out[1] <= Bit_822;data_out[2] <= Bit_823; data_out[3] <= Bit_824; end
		{1'b1, 16'd824}: begin data_out[0] <= Bit_825; data_out[1] <= Bit_826;data_out[2] <= Bit_827; data_out[3] <= Bit_828; end
		{1'b1, 16'd828}: begin data_out[0] <= Bit_829; data_out[1] <= Bit_830;data_out[2] <= Bit_831; data_out[3] <= Bit_832; end
		{1'b1, 16'd832}: begin data_out[0] <= Bit_833; data_out[1] <= Bit_834;data_out[2] <= Bit_835; data_out[3] <= Bit_836; end
		{1'b1, 16'd836}: begin data_out[0] <= Bit_837; data_out[1] <= Bit_838;data_out[2] <= Bit_839; data_out[3] <= Bit_840; end
		{1'b1, 16'd840}: begin data_out[0] <= Bit_841; data_out[1] <= Bit_842;data_out[2] <= Bit_843; data_out[3] <= Bit_844; end
		{1'b1, 16'd844}: begin data_out[0] <= Bit_845; data_out[1] <= Bit_846;data_out[2] <= Bit_847; data_out[3] <= Bit_848; end
		{1'b1, 16'd848}: begin data_out[0] <= Bit_849; data_out[1] <= Bit_850;data_out[2] <= Bit_851; data_out[3] <= Bit_852; end
		{1'b1, 16'd852}: begin data_out[0] <= Bit_853; data_out[1] <= Bit_854;data_out[2] <= Bit_855; data_out[3] <= Bit_856; end
		{1'b1, 16'd856}: begin data_out[0] <= Bit_857; data_out[1] <= Bit_858;data_out[2] <= Bit_859; data_out[3] <= Bit_860; end
		{1'b1, 16'd860}: begin data_out[0] <= Bit_861; data_out[1] <= Bit_862;data_out[2] <= Bit_863; data_out[3] <= Bit_864; end
		{1'b1, 16'd864}: begin data_out[0] <= Bit_865; data_out[1] <= Bit_866;data_out[2] <= Bit_867; data_out[3] <= Bit_868; end
		{1'b1, 16'd868}: begin data_out[0] <= Bit_869; data_out[1] <= Bit_870;data_out[2] <= Bit_871; data_out[3] <= Bit_872; end
		{1'b1, 16'd872}: begin data_out[0] <= Bit_873; data_out[1] <= Bit_874;data_out[2] <= Bit_875; data_out[3] <= Bit_876; end
		{1'b1, 16'd876}: begin data_out[0] <= Bit_877; data_out[1] <= Bit_878;data_out[2] <= Bit_879; data_out[3] <= Bit_880; end
		{1'b1, 16'd880}: begin data_out[0] <= Bit_881; data_out[1] <= Bit_882;data_out[2] <= Bit_883; data_out[3] <= Bit_884; end
		{1'b1, 16'd884}: begin data_out[0] <= Bit_885; data_out[1] <= Bit_886;data_out[2] <= Bit_887; data_out[3] <= Bit_888; end
		{1'b1, 16'd888}: begin data_out[0] <= Bit_889; data_out[1] <= Bit_890;data_out[2] <= Bit_891; data_out[3] <= Bit_892; end
		{1'b1, 16'd892}: begin data_out[0] <= Bit_893; data_out[1] <= Bit_894;data_out[2] <= Bit_895; data_out[3] <= Bit_896; end
		{1'b1, 16'd896}: begin data_out[0] <= Bit_897; data_out[1] <= Bit_898;data_out[2] <= Bit_899; data_out[3] <= Bit_900; end
		{1'b1, 16'd900}: begin data_out[0] <= Bit_901; data_out[1] <= Bit_902;data_out[2] <= Bit_903; data_out[3] <= Bit_904; end
		{1'b1, 16'd904}: begin data_out[0] <= Bit_905; data_out[1] <= Bit_906;data_out[2] <= Bit_907; data_out[3] <= Bit_908; end
		{1'b1, 16'd908}: begin data_out[0] <= Bit_909; data_out[1] <= Bit_910;data_out[2] <= Bit_911; data_out[3] <= Bit_912; end
		{1'b1, 16'd912}: begin data_out[0] <= Bit_913; data_out[1] <= Bit_914;data_out[2] <= Bit_915; data_out[3] <= Bit_916; end
		{1'b1, 16'd916}: begin data_out[0] <= Bit_917; data_out[1] <= Bit_918;data_out[2] <= Bit_919; data_out[3] <= Bit_920; end
		{1'b1, 16'd920}: begin data_out[0] <= Bit_921; data_out[1] <= Bit_922;data_out[2] <= Bit_923; data_out[3] <= Bit_924; end
		{1'b1, 16'd924}: begin data_out[0] <= Bit_925; data_out[1] <= Bit_926;data_out[2] <= Bit_927; data_out[3] <= Bit_928; end
		{1'b1, 16'd928}: begin data_out[0] <= Bit_929; data_out[1] <= Bit_930;data_out[2] <= Bit_931; data_out[3] <= Bit_932; end
		{1'b1, 16'd932}: begin data_out[0] <= Bit_933; data_out[1] <= Bit_934;data_out[2] <= Bit_935; data_out[3] <= Bit_936; end
		{1'b1, 16'd936}: begin data_out[0] <= Bit_937; data_out[1] <= Bit_938;data_out[2] <= Bit_939; data_out[3] <= Bit_940; end
		{1'b1, 16'd940}: begin data_out[0] <= Bit_941; data_out[1] <= Bit_942;data_out[2] <= Bit_943; data_out[3] <= Bit_944; end
		{1'b1, 16'd944}: begin data_out[0] <= Bit_945; data_out[1] <= Bit_946;data_out[2] <= Bit_947; data_out[3] <= Bit_948; end
		{1'b1, 16'd948}: begin data_out[0] <= Bit_949; data_out[1] <= Bit_950;data_out[2] <= Bit_951; data_out[3] <= Bit_952; end
		{1'b1, 16'd952}: begin data_out[0] <= Bit_953; data_out[1] <= Bit_954;data_out[2] <= Bit_955; data_out[3] <= Bit_956; end
		{1'b1, 16'd956}: begin data_out[0] <= Bit_957; data_out[1] <= Bit_958;data_out[2] <= Bit_959; data_out[3] <= Bit_960; end
		{1'b1, 16'd960}: begin data_out[0] <= Bit_961; data_out[1] <= Bit_962;data_out[2] <= Bit_963; data_out[3] <= Bit_964; end
		{1'b1, 16'd964}: begin data_out[0] <= Bit_965; data_out[1] <= Bit_966;data_out[2] <= Bit_967; data_out[3] <= Bit_968; end
		{1'b1, 16'd968}: begin data_out[0] <= Bit_969; data_out[1] <= Bit_970;data_out[2] <= Bit_971; data_out[3] <= Bit_972; end
		{1'b1, 16'd972}: begin data_out[0] <= Bit_973; data_out[1] <= Bit_974;data_out[2] <= Bit_975; data_out[3] <= Bit_976; end
		{1'b1, 16'd976}: begin data_out[0] <= Bit_977; data_out[1] <= Bit_978;data_out[2] <= Bit_979; data_out[3] <= Bit_980; end
		{1'b1, 16'd980}: begin data_out[0] <= Bit_981; data_out[1] <= Bit_982;data_out[2] <= Bit_983; data_out[3] <= Bit_984; end
		{1'b1, 16'd984}: begin data_out[0] <= Bit_985; data_out[1] <= Bit_986;data_out[2] <= Bit_987; data_out[3] <= Bit_988; end
		{1'b1, 16'd988}: begin data_out[0] <= Bit_989; data_out[1] <= Bit_990;data_out[2] <= Bit_991; data_out[3] <= Bit_992; end
		{1'b1, 16'd992}: begin data_out[0] <= Bit_993; data_out[1] <= Bit_994;data_out[2] <= Bit_995; data_out[3] <= Bit_996; end
		{1'b1, 16'd996}: begin data_out[0] <= Bit_997; data_out[1] <= Bit_998;data_out[2] <= Bit_999; data_out[3] <= Bit_1000; end
		{1'b1, 16'd1000}: begin data_out[0] <= Bit_1001; data_out[1] <= Bit_1002;data_out[2] <= Bit_1003; data_out[3] <= Bit_1004; end
		{1'b1, 16'd1004}: begin data_out[0] <= Bit_1005; data_out[1] <= Bit_1006;data_out[2] <= Bit_1007; data_out[3] <= Bit_1008; end
		{1'b1, 16'd1008}: begin data_out[0] <= Bit_1009; data_out[1] <= Bit_1010;data_out[2] <= Bit_1011; data_out[3] <= Bit_1012; end
		{1'b1, 16'd1012}: begin data_out[0] <= Bit_1013; data_out[1] <= Bit_1014;data_out[2] <= Bit_1015; data_out[3] <= Bit_1016; end
		{1'b1, 16'd1016}: begin data_out[0] <= Bit_1017; data_out[1] <= Bit_1018;data_out[2] <= Bit_1019; data_out[3] <= Bit_1020; end
		{1'b1, 16'd1020}: begin data_out[0] <= Bit_1021; data_out[1] <= Bit_1022;data_out[2] <= Bit_1023; data_out[3] <= Bit_1024; end
		{1'b1, 16'd1024}: begin data_out[0] <= Bit_1025; data_out[1] <= Bit_1026;data_out[2] <= Bit_1027; data_out[3] <= Bit_1028; end
		{1'b1, 16'd1028}: begin data_out[0] <= Bit_1029; data_out[1] <= Bit_1030;data_out[2] <= Bit_1031; data_out[3] <= Bit_1032; end
		{1'b1, 16'd1032}: begin data_out[0] <= Bit_1033; data_out[1] <= Bit_1034;data_out[2] <= Bit_1035; data_out[3] <= Bit_1036; end
		{1'b1, 16'd1036}: begin data_out[0] <= Bit_1037; data_out[1] <= Bit_1038;data_out[2] <= Bit_1039; data_out[3] <= Bit_1040; end
		{1'b1, 16'd1040}: begin data_out[0] <= Bit_1041; data_out[1] <= Bit_1042;data_out[2] <= Bit_1043; data_out[3] <= Bit_1044; end
		{1'b1, 16'd1044}: begin data_out[0] <= Bit_1045; data_out[1] <= Bit_1046;data_out[2] <= Bit_1047; data_out[3] <= Bit_1048; end
		{1'b1, 16'd1048}: begin data_out[0] <= Bit_1049; data_out[1] <= Bit_1050;data_out[2] <= Bit_1051; data_out[3] <= Bit_1052; end
		{1'b1, 16'd1052}: begin data_out[0] <= Bit_1053; data_out[1] <= Bit_1054;data_out[2] <= Bit_1055; data_out[3] <= Bit_1056; end
		{1'b1, 16'd1056}: begin data_out[0] <= Bit_1057; data_out[1] <= Bit_1058;data_out[2] <= Bit_1059; data_out[3] <= Bit_1060; end
		{1'b1, 16'd1060}: begin data_out[0] <= Bit_1061; data_out[1] <= Bit_1062;data_out[2] <= Bit_1063; data_out[3] <= Bit_1064; end
		{1'b1, 16'd1064}: begin data_out[0] <= Bit_1065; data_out[1] <= Bit_1066;data_out[2] <= Bit_1067; data_out[3] <= Bit_1068; end
		{1'b1, 16'd1068}: begin data_out[0] <= Bit_1069; data_out[1] <= Bit_1070;data_out[2] <= Bit_1071; data_out[3] <= Bit_1072; end
		{1'b1, 16'd1072}: begin data_out[0] <= Bit_1073; data_out[1] <= Bit_1074;data_out[2] <= Bit_1075; data_out[3] <= Bit_1076; end
		{1'b1, 16'd1076}: begin data_out[0] <= Bit_1077; data_out[1] <= Bit_1078;data_out[2] <= Bit_1079; data_out[3] <= Bit_1080; end
		{1'b1, 16'd1080}: begin data_out[0] <= Bit_1081; data_out[1] <= Bit_1082;data_out[2] <= Bit_1083; data_out[3] <= Bit_1084; end
		{1'b1, 16'd1084}: begin data_out[0] <= Bit_1085; data_out[1] <= Bit_1086;data_out[2] <= Bit_1087; data_out[3] <= Bit_1088; end
		{1'b1, 16'd1088}: begin data_out[0] <= Bit_1089; data_out[1] <= Bit_1090;data_out[2] <= Bit_1091; data_out[3] <= Bit_1092; end
		{1'b1, 16'd1092}: begin data_out[0] <= Bit_1093; data_out[1] <= Bit_1094;data_out[2] <= Bit_1095; data_out[3] <= Bit_1096; end
		{1'b1, 16'd1096}: begin data_out[0] <= Bit_1097; data_out[1] <= Bit_1098;data_out[2] <= Bit_1099; data_out[3] <= Bit_1100; end
		{1'b1, 16'd1100}: begin data_out[0] <= Bit_1101; data_out[1] <= Bit_1102;data_out[2] <= Bit_1103; data_out[3] <= Bit_1104; end
		{1'b1, 16'd1104}: begin data_out[0] <= Bit_1105; data_out[1] <= Bit_1106;data_out[2] <= Bit_1107; data_out[3] <= Bit_1108; end
		{1'b1, 16'd1108}: begin data_out[0] <= Bit_1109; data_out[1] <= Bit_1110;data_out[2] <= Bit_1111; data_out[3] <= Bit_1112; end
		{1'b1, 16'd1112}: begin data_out[0] <= Bit_1113; data_out[1] <= Bit_1114;data_out[2] <= Bit_1115; data_out[3] <= Bit_1116; end
		{1'b1, 16'd1116}: begin data_out[0] <= Bit_1117; data_out[1] <= Bit_1118;data_out[2] <= Bit_1119; data_out[3] <= Bit_1120; end
		{1'b1, 16'd1120}: begin data_out[0] <= Bit_1121; data_out[1] <= Bit_1122;data_out[2] <= Bit_1123; data_out[3] <= Bit_1124; end
		{1'b1, 16'd1124}: begin data_out[0] <= Bit_1125; data_out[1] <= Bit_1126;data_out[2] <= Bit_1127; data_out[3] <= Bit_1128; end
		{1'b1, 16'd1128}: begin data_out[0] <= Bit_1129; data_out[1] <= Bit_1130;data_out[2] <= Bit_1131; data_out[3] <= Bit_1132; end
		{1'b1, 16'd1132}: begin data_out[0] <= Bit_1133; data_out[1] <= Bit_1134;data_out[2] <= Bit_1135; data_out[3] <= Bit_1136; end
		{1'b1, 16'd1136}: begin data_out[0] <= Bit_1137; data_out[1] <= Bit_1138;data_out[2] <= Bit_1139; data_out[3] <= Bit_1140; end
		{1'b1, 16'd1140}: begin data_out[0] <= Bit_1141; data_out[1] <= Bit_1142;data_out[2] <= Bit_1143; data_out[3] <= Bit_1144; end
		{1'b1, 16'd1144}: begin data_out[0] <= Bit_1145; data_out[1] <= Bit_1146;data_out[2] <= Bit_1147; data_out[3] <= Bit_1148; end
		{1'b1, 16'd1148}: begin data_out[0] <= Bit_1149; data_out[1] <= Bit_1150;data_out[2] <= Bit_1151; data_out[3] <= Bit_1152; end
		{1'b1, 16'd1152}: begin data_out[0] <= Bit_1153; data_out[1] <= Bit_1154;data_out[2] <= Bit_1155; data_out[3] <= Bit_1156; end
		{1'b1, 16'd1156}: begin data_out[0] <= Bit_1157; data_out[1] <= Bit_1158;data_out[2] <= Bit_1159; data_out[3] <= Bit_1160; end
		{1'b1, 16'd1160}: begin data_out[0] <= Bit_1161; data_out[1] <= Bit_1162;data_out[2] <= Bit_1163; data_out[3] <= Bit_1164; end
		{1'b1, 16'd1164}: begin data_out[0] <= Bit_1165; data_out[1] <= Bit_1166;data_out[2] <= Bit_1167; data_out[3] <= Bit_1168; end
		{1'b1, 16'd1168}: begin data_out[0] <= Bit_1169; data_out[1] <= Bit_1170;data_out[2] <= Bit_1171; data_out[3] <= Bit_1172; end
		{1'b1, 16'd1172}: begin data_out[0] <= Bit_1173; data_out[1] <= Bit_1174;data_out[2] <= Bit_1175; data_out[3] <= Bit_1176; end
		{1'b1, 16'd1176}: begin data_out[0] <= Bit_1177; data_out[1] <= Bit_1178;data_out[2] <= Bit_1179; data_out[3] <= Bit_1180; end
		{1'b1, 16'd1180}: begin data_out[0] <= Bit_1181; data_out[1] <= Bit_1182;data_out[2] <= Bit_1183; data_out[3] <= Bit_1184; end
		{1'b1, 16'd1184}: begin data_out[0] <= Bit_1185; data_out[1] <= Bit_1186;data_out[2] <= Bit_1187; data_out[3] <= Bit_1188; end
		{1'b1, 16'd1188}: begin data_out[0] <= Bit_1189; data_out[1] <= Bit_1190;data_out[2] <= Bit_1191; data_out[3] <= Bit_1192; end
		{1'b1, 16'd1192}: begin data_out[0] <= Bit_1193; data_out[1] <= Bit_1194;data_out[2] <= Bit_1195; data_out[3] <= Bit_1196; end
		{1'b1, 16'd1196}: begin data_out[0] <= Bit_1197; data_out[1] <= Bit_1198;data_out[2] <= Bit_1199; data_out[3] <= Bit_1200; end
		{1'b1, 16'd1200}: begin data_out[0] <= Bit_1201; data_out[1] <= Bit_1202;data_out[2] <= Bit_1203; data_out[3] <= Bit_1204; end
		{1'b1, 16'd1204}: begin data_out[0] <= Bit_1205; data_out[1] <= Bit_1206;data_out[2] <= Bit_1207; data_out[3] <= Bit_1208; end
		{1'b1, 16'd1208}: begin data_out[0] <= Bit_1209; data_out[1] <= Bit_1210;data_out[2] <= Bit_1211; data_out[3] <= Bit_1212; end
		{1'b1, 16'd1212}: begin data_out[0] <= Bit_1213; data_out[1] <= Bit_1214;data_out[2] <= Bit_1215; data_out[3] <= Bit_1216; end
		{1'b1, 16'd1216}: begin data_out[0] <= Bit_1217; data_out[1] <= Bit_1218;data_out[2] <= Bit_1219; data_out[3] <= Bit_1220; end
		{1'b1, 16'd1220}: begin data_out[0] <= Bit_1221; data_out[1] <= Bit_1222;data_out[2] <= Bit_1223; data_out[3] <= Bit_1224; end
		{1'b1, 16'd1224}: begin data_out[0] <= Bit_1225; data_out[1] <= Bit_1226;data_out[2] <= Bit_1227; data_out[3] <= Bit_1228; end
		{1'b1, 16'd1228}: begin data_out[0] <= Bit_1229; data_out[1] <= Bit_1230;data_out[2] <= Bit_1231; data_out[3] <= Bit_1232; end
		{1'b1, 16'd1232}: begin data_out[0] <= Bit_1233; data_out[1] <= Bit_1234;data_out[2] <= Bit_1235; data_out[3] <= Bit_1236; end
		{1'b1, 16'd1236}: begin data_out[0] <= Bit_1237; data_out[1] <= Bit_1238;data_out[2] <= Bit_1239; data_out[3] <= Bit_1240; end
		{1'b1, 16'd1240}: begin data_out[0] <= Bit_1241; data_out[1] <= Bit_1242;data_out[2] <= Bit_1243; data_out[3] <= Bit_1244; end
		{1'b1, 16'd1244}: begin data_out[0] <= Bit_1245; data_out[1] <= Bit_1246;data_out[2] <= Bit_1247; data_out[3] <= Bit_1248; end
		{1'b1, 16'd1248}: begin data_out[0] <= Bit_1249; data_out[1] <= Bit_1250;data_out[2] <= Bit_1251; data_out[3] <= Bit_1252; end
		{1'b1, 16'd1252}: begin data_out[0] <= Bit_1253; data_out[1] <= Bit_1254;data_out[2] <= Bit_1255; data_out[3] <= Bit_1256; end
		{1'b1, 16'd1256}: begin data_out[0] <= Bit_1257; data_out[1] <= Bit_1258;data_out[2] <= Bit_1259; data_out[3] <= Bit_1260; end
		{1'b1, 16'd1260}: begin data_out[0] <= Bit_1261; data_out[1] <= Bit_1262;data_out[2] <= Bit_1263; data_out[3] <= Bit_1264; end
		{1'b1, 16'd1264}: begin data_out[0] <= Bit_1265; data_out[1] <= Bit_1266;data_out[2] <= Bit_1267; data_out[3] <= Bit_1268; end
		{1'b1, 16'd1268}: begin data_out[0] <= Bit_1269; data_out[1] <= Bit_1270;data_out[2] <= Bit_1271; data_out[3] <= Bit_1272; end
		{1'b1, 16'd1272}: begin data_out[0] <= Bit_1273; data_out[1] <= Bit_1274;data_out[2] <= Bit_1275; data_out[3] <= Bit_1276; end
		{1'b1, 16'd1276}: begin data_out[0] <= Bit_1277; data_out[1] <= Bit_1278;data_out[2] <= Bit_1279; data_out[3] <= Bit_1280; end
		{1'b1, 16'd1280}: begin data_out[0] <= Bit_1281; data_out[1] <= Bit_1282;data_out[2] <= Bit_1283; data_out[3] <= Bit_1284; end
		{1'b1, 16'd1284}: begin data_out[0] <= Bit_1285; data_out[1] <= Bit_1286;data_out[2] <= Bit_1287; data_out[3] <= Bit_1288; end
		{1'b1, 16'd1288}: begin data_out[0] <= Bit_1289; data_out[1] <= Bit_1290;data_out[2] <= Bit_1291; data_out[3] <= Bit_1292; end
		{1'b1, 16'd1292}: begin data_out[0] <= Bit_1293; data_out[1] <= Bit_1294;data_out[2] <= Bit_1295; data_out[3] <= Bit_1296; end
		{1'b1, 16'd1296}: begin data_out[0] <= Bit_1297; data_out[1] <= Bit_1298;data_out[2] <= Bit_1299; data_out[3] <= Bit_1300; end
		{1'b1, 16'd1300}: begin data_out[0] <= Bit_1301; data_out[1] <= Bit_1302;data_out[2] <= Bit_1303; data_out[3] <= Bit_1304; end
		{1'b1, 16'd1304}: begin data_out[0] <= Bit_1305; data_out[1] <= Bit_1306;data_out[2] <= Bit_1307; data_out[3] <= Bit_1308; end
		{1'b1, 16'd1308}: begin data_out[0] <= Bit_1309; data_out[1] <= Bit_1310;data_out[2] <= Bit_1311; data_out[3] <= Bit_1312; end
		{1'b1, 16'd1312}: begin data_out[0] <= Bit_1313; data_out[1] <= Bit_1314;data_out[2] <= Bit_1315; data_out[3] <= Bit_1316; end
		{1'b1, 16'd1316}: begin data_out[0] <= Bit_1317; data_out[1] <= Bit_1318;data_out[2] <= Bit_1319; data_out[3] <= Bit_1320; end
		{1'b1, 16'd1320}: begin data_out[0] <= Bit_1321; data_out[1] <= Bit_1322;data_out[2] <= Bit_1323; data_out[3] <= Bit_1324; end
		{1'b1, 16'd1324}: begin data_out[0] <= Bit_1325; data_out[1] <= Bit_1326;data_out[2] <= Bit_1327; data_out[3] <= Bit_1328; end
		{1'b1, 16'd1328}: begin data_out[0] <= Bit_1329; data_out[1] <= Bit_1330;data_out[2] <= Bit_1331; data_out[3] <= Bit_1332; end
		{1'b1, 16'd1332}: begin data_out[0] <= Bit_1333; data_out[1] <= Bit_1334;data_out[2] <= Bit_1335; data_out[3] <= Bit_1336; end
		{1'b1, 16'd1336}: begin data_out[0] <= Bit_1337; data_out[1] <= Bit_1338;data_out[2] <= Bit_1339; data_out[3] <= Bit_1340; end
		{1'b1, 16'd1340}: begin data_out[0] <= Bit_1341; data_out[1] <= Bit_1342;data_out[2] <= Bit_1343; data_out[3] <= Bit_1344; end
		{1'b1, 16'd1344}: begin data_out[0] <= Bit_1345; data_out[1] <= Bit_1346;data_out[2] <= Bit_1347; data_out[3] <= Bit_1348; end
		{1'b1, 16'd1348}: begin data_out[0] <= Bit_1349; data_out[1] <= Bit_1350;data_out[2] <= Bit_1351; data_out[3] <= Bit_1352; end
		{1'b1, 16'd1352}: begin data_out[0] <= Bit_1353; data_out[1] <= Bit_1354;data_out[2] <= Bit_1355; data_out[3] <= Bit_1356; end
		{1'b1, 16'd1356}: begin data_out[0] <= Bit_1357; data_out[1] <= Bit_1358;data_out[2] <= Bit_1359; data_out[3] <= Bit_1360; end
		{1'b1, 16'd1360}: begin data_out[0] <= Bit_1361; data_out[1] <= Bit_1362;data_out[2] <= Bit_1363; data_out[3] <= Bit_1364; end
		{1'b1, 16'd1364}: begin data_out[0] <= Bit_1365; data_out[1] <= Bit_1366;data_out[2] <= Bit_1367; data_out[3] <= Bit_1368; end
		{1'b1, 16'd1368}: begin data_out[0] <= Bit_1369; data_out[1] <= Bit_1370;data_out[2] <= Bit_1371; data_out[3] <= Bit_1372; end
		{1'b1, 16'd1372}: begin data_out[0] <= Bit_1373; data_out[1] <= Bit_1374;data_out[2] <= Bit_1375; data_out[3] <= Bit_1376; end
		{1'b1, 16'd1376}: begin data_out[0] <= Bit_1377; data_out[1] <= Bit_1378;data_out[2] <= Bit_1379; data_out[3] <= Bit_1380; end
		{1'b1, 16'd1380}: begin data_out[0] <= Bit_1381; data_out[1] <= Bit_1382;data_out[2] <= Bit_1383; data_out[3] <= Bit_1384; end
		{1'b1, 16'd1384}: begin data_out[0] <= Bit_1385; data_out[1] <= Bit_1386;data_out[2] <= Bit_1387; data_out[3] <= Bit_1388; end
		{1'b1, 16'd1388}: begin data_out[0] <= Bit_1389; data_out[1] <= Bit_1390;data_out[2] <= Bit_1391; data_out[3] <= Bit_1392; end
		{1'b1, 16'd1392}: begin data_out[0] <= Bit_1393; data_out[1] <= Bit_1394;data_out[2] <= Bit_1395; data_out[3] <= Bit_1396; end
		{1'b1, 16'd1396}: begin data_out[0] <= Bit_1397; data_out[1] <= Bit_1398;data_out[2] <= Bit_1399; data_out[3] <= Bit_1400; end
		{1'b1, 16'd1400}: begin data_out[0] <= Bit_1401; data_out[1] <= Bit_1402;data_out[2] <= Bit_1403; data_out[3] <= Bit_1404; end
		{1'b1, 16'd1404}: begin data_out[0] <= Bit_1405; data_out[1] <= Bit_1406;data_out[2] <= Bit_1407; data_out[3] <= Bit_1408; end
		{1'b1, 16'd1408}: begin data_out[0] <= Bit_1409; data_out[1] <= Bit_1410;data_out[2] <= Bit_1411; data_out[3] <= Bit_1412; end
		{1'b1, 16'd1412}: begin data_out[0] <= Bit_1413; data_out[1] <= Bit_1414;data_out[2] <= Bit_1415; data_out[3] <= Bit_1416; end
		{1'b1, 16'd1416}: begin data_out[0] <= Bit_1417; data_out[1] <= Bit_1418;data_out[2] <= Bit_1419; data_out[3] <= Bit_1420; end
		{1'b1, 16'd1420}: begin data_out[0] <= Bit_1421; data_out[1] <= Bit_1422;data_out[2] <= Bit_1423; data_out[3] <= Bit_1424; end
		{1'b1, 16'd1424}: begin data_out[0] <= Bit_1425; data_out[1] <= Bit_1426;data_out[2] <= Bit_1427; data_out[3] <= Bit_1428; end
		{1'b1, 16'd1428}: begin data_out[0] <= Bit_1429; data_out[1] <= Bit_1430;data_out[2] <= Bit_1431; data_out[3] <= Bit_1432; end
		{1'b1, 16'd1432}: begin data_out[0] <= Bit_1433; data_out[1] <= Bit_1434;data_out[2] <= Bit_1435; data_out[3] <= Bit_1436; end
		{1'b1, 16'd1436}: begin data_out[0] <= Bit_1437; data_out[1] <= Bit_1438;data_out[2] <= Bit_1439; data_out[3] <= Bit_1440; end
	endcase
end

always @ (posedge clk) begin
if (out_valid == 1) begin
if (out_index < code_length - 4)
out_index <= out_index + 4;
else
out_valid <= 0;
end
end

always @ (posedge clk or negedge rst) begin
	if (!rst) begin
		cnt <= 0;
		iter <= 0;
		out_valid <= 0;
		out_index <= 0;
		data_out <= 4'd0;
		Check_1 <= 1;
		Check_2 <= 1;
		Check_3 <= 1;
		Check_4 <= 1;
		Check_5 <= 1;
		Check_6 <= 1;
		Check_7 <= 1;
		Check_8 <= 1;
		Check_9 <= 1;
		Check_10 <= 1;
		Check_11 <= 1;
		Check_12 <= 1;
		Check_13 <= 1;
		Check_14 <= 1;
		Check_15 <= 1;
		Check_16 <= 1;
		Check_17 <= 1;
		Check_18 <= 1;
		Check_19 <= 1;
		Check_20 <= 1;
		Check_21 <= 1;
		Check_22 <= 1;
		Check_23 <= 1;
		Check_24 <= 1;
		Check_25 <= 1;
		Check_26 <= 1;
		Check_27 <= 1;
		Check_28 <= 1;
		Check_29 <= 1;
		Check_30 <= 1;
		Check_31 <= 1;
		Check_32 <= 1;
		Check_33 <= 1;
		Check_34 <= 1;
		Check_35 <= 1;
		Check_36 <= 1;
		Check_37 <= 1;
		Check_38 <= 1;
		Check_39 <= 1;
		Check_40 <= 1;
		Check_41 <= 1;
		Check_42 <= 1;
		Check_43 <= 1;
		Check_44 <= 1;
		Check_45 <= 1;
		Check_46 <= 1;
		Check_47 <= 1;
		Check_48 <= 1;
		Check_49 <= 1;
		Check_50 <= 1;
		Check_51 <= 1;
		Check_52 <= 1;
		Check_53 <= 1;
		Check_54 <= 1;
		Check_55 <= 1;
		Check_56 <= 1;
		Check_57 <= 1;
		Check_58 <= 1;
		Check_59 <= 1;
		Check_60 <= 1;
		Check_61 <= 1;
		Check_62 <= 1;
		Check_63 <= 1;
		Check_64 <= 1;
		Check_65 <= 1;
		Check_66 <= 1;
		Check_67 <= 1;
		Check_68 <= 1;
		Check_69 <= 1;
		Check_70 <= 1;
		Check_71 <= 1;
		Check_72 <= 1;
		Check_73 <= 1;
		Check_74 <= 1;
		Check_75 <= 1;
		Check_76 <= 1;
		Check_77 <= 1;
		Check_78 <= 1;
		Check_79 <= 1;
		Check_80 <= 1;
		Check_81 <= 1;
		Check_82 <= 1;
		Check_83 <= 1;
		Check_84 <= 1;
		Check_85 <= 1;
		Check_86 <= 1;
		Check_87 <= 1;
		Check_88 <= 1;
		Check_89 <= 1;
		Check_90 <= 1;
		Check_91 <= 1;
		Check_92 <= 1;
		Check_93 <= 1;
		Check_94 <= 1;
		Check_95 <= 1;
		Check_96 <= 1;
		Check_97 <= 1;
		Check_98 <= 1;
		Check_99 <= 1;
		Check_100 <= 1;
		Check_101 <= 1;
		Check_102 <= 1;
		Check_103 <= 1;
		Check_104 <= 1;
		Check_105 <= 1;
		Check_106 <= 1;
		Check_107 <= 1;
		Check_108 <= 1;
		Check_109 <= 1;
		Check_110 <= 1;
		Check_111 <= 1;
		Check_112 <= 1;
		Check_113 <= 1;
		Check_114 <= 1;
		Check_115 <= 1;
		Check_116 <= 1;
		Check_117 <= 1;
		Check_118 <= 1;
		Check_119 <= 1;
		Check_120 <= 1;
		Check_121 <= 1;
		Check_122 <= 1;
		Check_123 <= 1;
		Check_124 <= 1;
		Check_125 <= 1;
		Check_126 <= 1;
		Check_127 <= 1;
		Check_128 <= 1;
		Check_129 <= 1;
		Check_130 <= 1;
		Check_131 <= 1;
		Check_132 <= 1;
		Check_133 <= 1;
		Check_134 <= 1;
		Check_135 <= 1;
		Check_136 <= 1;
		Check_137 <= 1;
		Check_138 <= 1;
		Check_139 <= 1;
		Check_140 <= 1;
		Check_141 <= 1;
		Check_142 <= 1;
		Check_143 <= 1;
		Check_144 <= 1;
		Check_145 <= 1;
		Check_146 <= 1;
		Check_147 <= 1;
		Check_148 <= 1;
		Check_149 <= 1;
		Check_150 <= 1;
		Check_151 <= 1;
		Check_152 <= 1;
		Check_153 <= 1;
		Check_154 <= 1;
		Check_155 <= 1;
		Check_156 <= 1;
		Check_157 <= 1;
		Check_158 <= 1;
		Check_159 <= 1;
		Check_160 <= 1;
		Check_161 <= 1;
		Check_162 <= 1;
		Check_163 <= 1;
		Check_164 <= 1;
		Check_165 <= 1;
		Check_166 <= 1;
		Check_167 <= 1;
		Check_168 <= 1;
		Check_169 <= 1;
		Check_170 <= 1;
		Check_171 <= 1;
		Check_172 <= 1;
		Check_173 <= 1;
		Check_174 <= 1;
		Check_175 <= 1;
		Check_176 <= 1;
		Check_177 <= 1;
		Check_178 <= 1;
		Check_179 <= 1;
		Check_180 <= 1;
		Check_181 <= 1;
		Check_182 <= 1;
		Check_183 <= 1;
		Check_184 <= 1;
		Check_185 <= 1;
		Check_186 <= 1;
		Check_187 <= 1;
		Check_188 <= 1;
		Check_189 <= 1;
		Check_190 <= 1;
		Check_191 <= 1;
		Check_192 <= 1;
		Check_193 <= 1;
		Check_194 <= 1;
		Check_195 <= 1;
		Check_196 <= 1;
		Check_197 <= 1;
		Check_198 <= 1;
		Check_199 <= 1;
		Check_200 <= 1;
		Check_201 <= 1;
		Check_202 <= 1;
		Check_203 <= 1;
		Check_204 <= 1;
		Check_205 <= 1;
		Check_206 <= 1;
		Check_207 <= 1;
		Check_208 <= 1;
		Check_209 <= 1;
		Check_210 <= 1;
		Check_211 <= 1;
		Check_212 <= 1;
		Check_213 <= 1;
		Check_214 <= 1;
		Check_215 <= 1;
		Check_216 <= 1;
		Check_217 <= 1;
		Check_218 <= 1;
		Check_219 <= 1;
		Check_220 <= 1;
		Check_221 <= 1;
		Check_222 <= 1;
		Check_223 <= 1;
		Check_224 <= 1;
		Check_225 <= 1;
		Check_226 <= 1;
		Check_227 <= 1;
		Check_228 <= 1;
		Check_229 <= 1;
		Check_230 <= 1;
		Check_231 <= 1;
		Check_232 <= 1;
		Check_233 <= 1;
		Check_234 <= 1;
		Check_235 <= 1;
		Check_236 <= 1;
		Check_237 <= 1;
		Check_238 <= 1;
		Check_239 <= 1;
		Check_240 <= 1;
		Check_241 <= 1;
		Check_242 <= 1;
		Check_243 <= 1;
		Check_244 <= 1;
		Check_245 <= 1;
		Check_246 <= 1;
		Check_247 <= 1;
		Check_248 <= 1;
		Check_249 <= 1;
		Check_250 <= 1;
		Check_251 <= 1;
		Check_252 <= 1;
		Check_253 <= 1;
		Check_254 <= 1;
		Check_255 <= 1;
		Check_256 <= 1;
		Check_257 <= 1;
		Check_258 <= 1;
		Check_259 <= 1;
		Check_260 <= 1;
		Check_261 <= 1;
		Check_262 <= 1;
		Check_263 <= 1;
		Check_264 <= 1;
		Check_265 <= 1;
		Check_266 <= 1;
		Check_267 <= 1;
		Check_268 <= 1;
		Check_269 <= 1;
		Check_270 <= 1;
		Check_271 <= 1;
		Check_272 <= 1;
		Check_273 <= 1;
		Check_274 <= 1;
		Check_275 <= 1;
		Check_276 <= 1;
		Check_277 <= 1;
		Check_278 <= 1;
		Check_279 <= 1;
		Check_280 <= 1;
		Check_281 <= 1;
		Check_282 <= 1;
		Check_283 <= 1;
		Check_284 <= 1;
		Check_285 <= 1;
		Check_286 <= 1;
		Check_287 <= 1;
		Check_288 <= 1;
		Check_Sum <= 1;
	end
	else begin
		if (out_valid == 0) begin
			if (8'd0 < cnt && cnt < 8'd15)
			cnt <= cnt + 1;
			else if (cnt == 8'd15) begin
				Check_1 <= Bit_5 ^ Bit_89 ^ Bit_109 ^ Bit_170 ^ Bit_232 ^ Bit_275 ^ Bit_375 ^ Bit_429 ^ Bit_526 ^ Bit_762 ^ Bit_810 ^ Bit_858 ^ Bit_899 ^ Bit_940 ^ Bit_974 ^ Bit_1013 ^ Bit_1087 ^ Bit_1146 ^ Bit_1153;
				Check_2 <= Bit_14 ^ Bit_63 ^ Bit_119 ^ Bit_167 ^ Bit_196 ^ Bit_265 ^ Bit_316 ^ Bit_423 ^ Bit_512 ^ Bit_672 ^ Bit_685 ^ Bit_853 ^ Bit_895 ^ Bit_958 ^ Bit_989 ^ Bit_1021 ^ Bit_1088 ^ Bit_1119 ^ Bit_1153 ^ Bit_1154;
				Check_3 <= Bit_9 ^ Bit_84 ^ Bit_101 ^ Bit_183 ^ Bit_201 ^ Bit_268 ^ Bit_365 ^ Bit_420 ^ Bit_531 ^ Bit_588 ^ Bit_664 ^ Bit_768 ^ Bit_899 ^ Bit_943 ^ Bit_968 ^ Bit_1028 ^ Bit_1058 ^ Bit_1151 ^ Bit_1154 ^ Bit_1155;
				Check_4 <= Bit_28 ^ Bit_87 ^ Bit_126 ^ Bit_182 ^ Bit_199 ^ Bit_253 ^ Bit_477 ^ Bit_517 ^ Bit_553 ^ Bit_615 ^ Bit_640 ^ Bit_686 ^ Bit_903 ^ Bit_927 ^ Bit_963 ^ Bit_1041 ^ Bit_1068 ^ Bit_1132 ^ Bit_1155 ^ Bit_1156;
				Check_5 <= Bit_47 ^ Bit_57 ^ Bit_140 ^ Bit_163 ^ Bit_227 ^ Bit_245 ^ Bit_294 ^ Bit_361 ^ Bit_440 ^ Bit_674 ^ Bit_738 ^ Bit_792 ^ Bit_870 ^ Bit_918 ^ Bit_961 ^ Bit_1013 ^ Bit_1062 ^ Bit_1110 ^ Bit_1156 ^ Bit_1157;
				Check_6 <= Bit_30 ^ Bit_54 ^ Bit_142 ^ Bit_162 ^ Bit_196 ^ Bit_275 ^ Bit_328 ^ Bit_480 ^ Bit_529 ^ Bit_610 ^ Bit_814 ^ Bit_842 ^ Bit_875 ^ Bit_937 ^ Bit_972 ^ Bit_1039 ^ Bit_1103 ^ Bit_1105 ^ Bit_1157 ^ Bit_1158;
				Check_7 <= Bit_6 ^ Bit_90 ^ Bit_110 ^ Bit_171 ^ Bit_233 ^ Bit_276 ^ Bit_376 ^ Bit_430 ^ Bit_527 ^ Bit_763 ^ Bit_811 ^ Bit_859 ^ Bit_900 ^ Bit_941 ^ Bit_975 ^ Bit_1014 ^ Bit_1088 ^ Bit_1147 ^ Bit_1158 ^ Bit_1159;
				Check_8 <= Bit_15 ^ Bit_64 ^ Bit_120 ^ Bit_168 ^ Bit_197 ^ Bit_266 ^ Bit_317 ^ Bit_424 ^ Bit_513 ^ Bit_625 ^ Bit_686 ^ Bit_854 ^ Bit_896 ^ Bit_959 ^ Bit_990 ^ Bit_1022 ^ Bit_1089 ^ Bit_1120 ^ Bit_1159 ^ Bit_1160;
				Check_9 <= Bit_10 ^ Bit_85 ^ Bit_102 ^ Bit_184 ^ Bit_202 ^ Bit_269 ^ Bit_366 ^ Bit_421 ^ Bit_532 ^ Bit_589 ^ Bit_665 ^ Bit_721 ^ Bit_900 ^ Bit_944 ^ Bit_969 ^ Bit_1029 ^ Bit_1059 ^ Bit_1152 ^ Bit_1160 ^ Bit_1161;
				Check_10 <= Bit_29 ^ Bit_88 ^ Bit_127 ^ Bit_183 ^ Bit_200 ^ Bit_254 ^ Bit_478 ^ Bit_518 ^ Bit_554 ^ Bit_616 ^ Bit_641 ^ Bit_687 ^ Bit_904 ^ Bit_928 ^ Bit_964 ^ Bit_1042 ^ Bit_1069 ^ Bit_1133 ^ Bit_1161 ^ Bit_1162;
				Check_11 <= Bit_48 ^ Bit_58 ^ Bit_141 ^ Bit_164 ^ Bit_228 ^ Bit_246 ^ Bit_295 ^ Bit_362 ^ Bit_441 ^ Bit_675 ^ Bit_739 ^ Bit_793 ^ Bit_871 ^ Bit_919 ^ Bit_962 ^ Bit_1014 ^ Bit_1063 ^ Bit_1111 ^ Bit_1162 ^ Bit_1163;
				Check_12 <= Bit_31 ^ Bit_55 ^ Bit_143 ^ Bit_163 ^ Bit_197 ^ Bit_276 ^ Bit_329 ^ Bit_433 ^ Bit_530 ^ Bit_611 ^ Bit_815 ^ Bit_843 ^ Bit_876 ^ Bit_938 ^ Bit_973 ^ Bit_1040 ^ Bit_1104 ^ Bit_1106 ^ Bit_1163 ^ Bit_1164;
				Check_13 <= Bit_7 ^ Bit_91 ^ Bit_111 ^ Bit_172 ^ Bit_234 ^ Bit_277 ^ Bit_377 ^ Bit_431 ^ Bit_528 ^ Bit_764 ^ Bit_812 ^ Bit_860 ^ Bit_901 ^ Bit_942 ^ Bit_976 ^ Bit_1015 ^ Bit_1089 ^ Bit_1148 ^ Bit_1164 ^ Bit_1165;
				Check_14 <= Bit_16 ^ Bit_65 ^ Bit_121 ^ Bit_169 ^ Bit_198 ^ Bit_267 ^ Bit_318 ^ Bit_425 ^ Bit_514 ^ Bit_626 ^ Bit_687 ^ Bit_855 ^ Bit_897 ^ Bit_960 ^ Bit_991 ^ Bit_1023 ^ Bit_1090 ^ Bit_1121 ^ Bit_1165 ^ Bit_1166;
				Check_15 <= Bit_11 ^ Bit_86 ^ Bit_103 ^ Bit_185 ^ Bit_203 ^ Bit_270 ^ Bit_367 ^ Bit_422 ^ Bit_533 ^ Bit_590 ^ Bit_666 ^ Bit_722 ^ Bit_901 ^ Bit_945 ^ Bit_970 ^ Bit_1030 ^ Bit_1060 ^ Bit_1105 ^ Bit_1166 ^ Bit_1167;
				Check_16 <= Bit_30 ^ Bit_89 ^ Bit_128 ^ Bit_184 ^ Bit_201 ^ Bit_255 ^ Bit_479 ^ Bit_519 ^ Bit_555 ^ Bit_617 ^ Bit_642 ^ Bit_688 ^ Bit_905 ^ Bit_929 ^ Bit_965 ^ Bit_1043 ^ Bit_1070 ^ Bit_1134 ^ Bit_1167 ^ Bit_1168;
				Check_17 <= Bit_1 ^ Bit_59 ^ Bit_142 ^ Bit_165 ^ Bit_229 ^ Bit_247 ^ Bit_296 ^ Bit_363 ^ Bit_442 ^ Bit_676 ^ Bit_740 ^ Bit_794 ^ Bit_872 ^ Bit_920 ^ Bit_963 ^ Bit_1015 ^ Bit_1064 ^ Bit_1112 ^ Bit_1168 ^ Bit_1169;
				Check_18 <= Bit_32 ^ Bit_56 ^ Bit_144 ^ Bit_164 ^ Bit_198 ^ Bit_277 ^ Bit_330 ^ Bit_434 ^ Bit_531 ^ Bit_612 ^ Bit_816 ^ Bit_844 ^ Bit_877 ^ Bit_939 ^ Bit_974 ^ Bit_1041 ^ Bit_1057 ^ Bit_1107 ^ Bit_1169 ^ Bit_1170;
				Check_19 <= Bit_8 ^ Bit_92 ^ Bit_112 ^ Bit_173 ^ Bit_235 ^ Bit_278 ^ Bit_378 ^ Bit_432 ^ Bit_481 ^ Bit_765 ^ Bit_813 ^ Bit_861 ^ Bit_902 ^ Bit_943 ^ Bit_977 ^ Bit_1016 ^ Bit_1090 ^ Bit_1149 ^ Bit_1170 ^ Bit_1171;
				Check_20 <= Bit_17 ^ Bit_66 ^ Bit_122 ^ Bit_170 ^ Bit_199 ^ Bit_268 ^ Bit_319 ^ Bit_426 ^ Bit_515 ^ Bit_627 ^ Bit_688 ^ Bit_856 ^ Bit_898 ^ Bit_913 ^ Bit_992 ^ Bit_1024 ^ Bit_1091 ^ Bit_1122 ^ Bit_1171 ^ Bit_1172;
				Check_21 <= Bit_12 ^ Bit_87 ^ Bit_104 ^ Bit_186 ^ Bit_204 ^ Bit_271 ^ Bit_368 ^ Bit_423 ^ Bit_534 ^ Bit_591 ^ Bit_667 ^ Bit_723 ^ Bit_902 ^ Bit_946 ^ Bit_971 ^ Bit_1031 ^ Bit_1061 ^ Bit_1106 ^ Bit_1172 ^ Bit_1173;
				Check_22 <= Bit_31 ^ Bit_90 ^ Bit_129 ^ Bit_185 ^ Bit_202 ^ Bit_256 ^ Bit_480 ^ Bit_520 ^ Bit_556 ^ Bit_618 ^ Bit_643 ^ Bit_689 ^ Bit_906 ^ Bit_930 ^ Bit_966 ^ Bit_1044 ^ Bit_1071 ^ Bit_1135 ^ Bit_1173 ^ Bit_1174;
				Check_23 <= Bit_2 ^ Bit_60 ^ Bit_143 ^ Bit_166 ^ Bit_230 ^ Bit_248 ^ Bit_297 ^ Bit_364 ^ Bit_443 ^ Bit_677 ^ Bit_741 ^ Bit_795 ^ Bit_873 ^ Bit_921 ^ Bit_964 ^ Bit_1016 ^ Bit_1065 ^ Bit_1113 ^ Bit_1174 ^ Bit_1175;
				Check_24 <= Bit_33 ^ Bit_57 ^ Bit_97 ^ Bit_165 ^ Bit_199 ^ Bit_278 ^ Bit_331 ^ Bit_435 ^ Bit_532 ^ Bit_613 ^ Bit_769 ^ Bit_845 ^ Bit_878 ^ Bit_940 ^ Bit_975 ^ Bit_1042 ^ Bit_1058 ^ Bit_1108 ^ Bit_1175 ^ Bit_1176;
				Check_25 <= Bit_9 ^ Bit_93 ^ Bit_113 ^ Bit_174 ^ Bit_236 ^ Bit_279 ^ Bit_379 ^ Bit_385 ^ Bit_482 ^ Bit_766 ^ Bit_814 ^ Bit_862 ^ Bit_903 ^ Bit_944 ^ Bit_978 ^ Bit_1017 ^ Bit_1091 ^ Bit_1150 ^ Bit_1176 ^ Bit_1177;
				Check_26 <= Bit_18 ^ Bit_67 ^ Bit_123 ^ Bit_171 ^ Bit_200 ^ Bit_269 ^ Bit_320 ^ Bit_427 ^ Bit_516 ^ Bit_628 ^ Bit_689 ^ Bit_857 ^ Bit_899 ^ Bit_914 ^ Bit_993 ^ Bit_1025 ^ Bit_1092 ^ Bit_1123 ^ Bit_1177 ^ Bit_1178;
				Check_27 <= Bit_13 ^ Bit_88 ^ Bit_105 ^ Bit_187 ^ Bit_205 ^ Bit_272 ^ Bit_369 ^ Bit_424 ^ Bit_535 ^ Bit_592 ^ Bit_668 ^ Bit_724 ^ Bit_903 ^ Bit_947 ^ Bit_972 ^ Bit_1032 ^ Bit_1062 ^ Bit_1107 ^ Bit_1178 ^ Bit_1179;
				Check_28 <= Bit_32 ^ Bit_91 ^ Bit_130 ^ Bit_186 ^ Bit_203 ^ Bit_257 ^ Bit_433 ^ Bit_521 ^ Bit_557 ^ Bit_619 ^ Bit_644 ^ Bit_690 ^ Bit_907 ^ Bit_931 ^ Bit_967 ^ Bit_1045 ^ Bit_1072 ^ Bit_1136 ^ Bit_1179 ^ Bit_1180;
				Check_29 <= Bit_3 ^ Bit_61 ^ Bit_144 ^ Bit_167 ^ Bit_231 ^ Bit_249 ^ Bit_298 ^ Bit_365 ^ Bit_444 ^ Bit_678 ^ Bit_742 ^ Bit_796 ^ Bit_874 ^ Bit_922 ^ Bit_965 ^ Bit_1017 ^ Bit_1066 ^ Bit_1114 ^ Bit_1180 ^ Bit_1181;
				Check_30 <= Bit_34 ^ Bit_58 ^ Bit_98 ^ Bit_166 ^ Bit_200 ^ Bit_279 ^ Bit_332 ^ Bit_436 ^ Bit_533 ^ Bit_614 ^ Bit_770 ^ Bit_846 ^ Bit_879 ^ Bit_941 ^ Bit_976 ^ Bit_1043 ^ Bit_1059 ^ Bit_1109 ^ Bit_1181 ^ Bit_1182;
				Check_31 <= Bit_10 ^ Bit_94 ^ Bit_114 ^ Bit_175 ^ Bit_237 ^ Bit_280 ^ Bit_380 ^ Bit_386 ^ Bit_483 ^ Bit_767 ^ Bit_815 ^ Bit_863 ^ Bit_904 ^ Bit_945 ^ Bit_979 ^ Bit_1018 ^ Bit_1092 ^ Bit_1151 ^ Bit_1182 ^ Bit_1183;
				Check_32 <= Bit_19 ^ Bit_68 ^ Bit_124 ^ Bit_172 ^ Bit_201 ^ Bit_270 ^ Bit_321 ^ Bit_428 ^ Bit_517 ^ Bit_629 ^ Bit_690 ^ Bit_858 ^ Bit_900 ^ Bit_915 ^ Bit_994 ^ Bit_1026 ^ Bit_1093 ^ Bit_1124 ^ Bit_1183 ^ Bit_1184;
				Check_33 <= Bit_14 ^ Bit_89 ^ Bit_106 ^ Bit_188 ^ Bit_206 ^ Bit_273 ^ Bit_370 ^ Bit_425 ^ Bit_536 ^ Bit_593 ^ Bit_669 ^ Bit_725 ^ Bit_904 ^ Bit_948 ^ Bit_973 ^ Bit_1033 ^ Bit_1063 ^ Bit_1108 ^ Bit_1184 ^ Bit_1185;
				Check_34 <= Bit_33 ^ Bit_92 ^ Bit_131 ^ Bit_187 ^ Bit_204 ^ Bit_258 ^ Bit_434 ^ Bit_522 ^ Bit_558 ^ Bit_620 ^ Bit_645 ^ Bit_691 ^ Bit_908 ^ Bit_932 ^ Bit_968 ^ Bit_1046 ^ Bit_1073 ^ Bit_1137 ^ Bit_1185 ^ Bit_1186;
				Check_35 <= Bit_4 ^ Bit_62 ^ Bit_97 ^ Bit_168 ^ Bit_232 ^ Bit_250 ^ Bit_299 ^ Bit_366 ^ Bit_445 ^ Bit_679 ^ Bit_743 ^ Bit_797 ^ Bit_875 ^ Bit_923 ^ Bit_966 ^ Bit_1018 ^ Bit_1067 ^ Bit_1115 ^ Bit_1186 ^ Bit_1187;
				Check_36 <= Bit_35 ^ Bit_59 ^ Bit_99 ^ Bit_167 ^ Bit_201 ^ Bit_280 ^ Bit_333 ^ Bit_437 ^ Bit_534 ^ Bit_615 ^ Bit_771 ^ Bit_847 ^ Bit_880 ^ Bit_942 ^ Bit_977 ^ Bit_1044 ^ Bit_1060 ^ Bit_1110 ^ Bit_1187 ^ Bit_1188;
				Check_37 <= Bit_11 ^ Bit_95 ^ Bit_115 ^ Bit_176 ^ Bit_238 ^ Bit_281 ^ Bit_381 ^ Bit_387 ^ Bit_484 ^ Bit_768 ^ Bit_816 ^ Bit_864 ^ Bit_905 ^ Bit_946 ^ Bit_980 ^ Bit_1019 ^ Bit_1093 ^ Bit_1152 ^ Bit_1188 ^ Bit_1189;
				Check_38 <= Bit_20 ^ Bit_69 ^ Bit_125 ^ Bit_173 ^ Bit_202 ^ Bit_271 ^ Bit_322 ^ Bit_429 ^ Bit_518 ^ Bit_630 ^ Bit_691 ^ Bit_859 ^ Bit_901 ^ Bit_916 ^ Bit_995 ^ Bit_1027 ^ Bit_1094 ^ Bit_1125 ^ Bit_1189 ^ Bit_1190;
				Check_39 <= Bit_15 ^ Bit_90 ^ Bit_107 ^ Bit_189 ^ Bit_207 ^ Bit_274 ^ Bit_371 ^ Bit_426 ^ Bit_537 ^ Bit_594 ^ Bit_670 ^ Bit_726 ^ Bit_905 ^ Bit_949 ^ Bit_974 ^ Bit_1034 ^ Bit_1064 ^ Bit_1109 ^ Bit_1190 ^ Bit_1191;
				Check_40 <= Bit_34 ^ Bit_93 ^ Bit_132 ^ Bit_188 ^ Bit_205 ^ Bit_259 ^ Bit_435 ^ Bit_523 ^ Bit_559 ^ Bit_621 ^ Bit_646 ^ Bit_692 ^ Bit_909 ^ Bit_933 ^ Bit_969 ^ Bit_1047 ^ Bit_1074 ^ Bit_1138 ^ Bit_1191 ^ Bit_1192;
				Check_41 <= Bit_5 ^ Bit_63 ^ Bit_98 ^ Bit_169 ^ Bit_233 ^ Bit_251 ^ Bit_300 ^ Bit_367 ^ Bit_446 ^ Bit_680 ^ Bit_744 ^ Bit_798 ^ Bit_876 ^ Bit_924 ^ Bit_967 ^ Bit_1019 ^ Bit_1068 ^ Bit_1116 ^ Bit_1192 ^ Bit_1193;
				Check_42 <= Bit_36 ^ Bit_60 ^ Bit_100 ^ Bit_168 ^ Bit_202 ^ Bit_281 ^ Bit_334 ^ Bit_438 ^ Bit_535 ^ Bit_616 ^ Bit_772 ^ Bit_848 ^ Bit_881 ^ Bit_943 ^ Bit_978 ^ Bit_1045 ^ Bit_1061 ^ Bit_1111 ^ Bit_1193 ^ Bit_1194;
				Check_43 <= Bit_12 ^ Bit_96 ^ Bit_116 ^ Bit_177 ^ Bit_239 ^ Bit_282 ^ Bit_382 ^ Bit_388 ^ Bit_485 ^ Bit_721 ^ Bit_769 ^ Bit_817 ^ Bit_906 ^ Bit_947 ^ Bit_981 ^ Bit_1020 ^ Bit_1094 ^ Bit_1105 ^ Bit_1194 ^ Bit_1195;
				Check_44 <= Bit_21 ^ Bit_70 ^ Bit_126 ^ Bit_174 ^ Bit_203 ^ Bit_272 ^ Bit_323 ^ Bit_430 ^ Bit_519 ^ Bit_631 ^ Bit_692 ^ Bit_860 ^ Bit_902 ^ Bit_917 ^ Bit_996 ^ Bit_1028 ^ Bit_1095 ^ Bit_1126 ^ Bit_1195 ^ Bit_1196;
				Check_45 <= Bit_16 ^ Bit_91 ^ Bit_108 ^ Bit_190 ^ Bit_208 ^ Bit_275 ^ Bit_372 ^ Bit_427 ^ Bit_538 ^ Bit_595 ^ Bit_671 ^ Bit_727 ^ Bit_906 ^ Bit_950 ^ Bit_975 ^ Bit_1035 ^ Bit_1065 ^ Bit_1110 ^ Bit_1196 ^ Bit_1197;
				Check_46 <= Bit_35 ^ Bit_94 ^ Bit_133 ^ Bit_189 ^ Bit_206 ^ Bit_260 ^ Bit_436 ^ Bit_524 ^ Bit_560 ^ Bit_622 ^ Bit_647 ^ Bit_693 ^ Bit_910 ^ Bit_934 ^ Bit_970 ^ Bit_1048 ^ Bit_1075 ^ Bit_1139 ^ Bit_1197 ^ Bit_1198;
				Check_47 <= Bit_6 ^ Bit_64 ^ Bit_99 ^ Bit_170 ^ Bit_234 ^ Bit_252 ^ Bit_301 ^ Bit_368 ^ Bit_447 ^ Bit_681 ^ Bit_745 ^ Bit_799 ^ Bit_877 ^ Bit_925 ^ Bit_968 ^ Bit_1020 ^ Bit_1069 ^ Bit_1117 ^ Bit_1198 ^ Bit_1199;
				Check_48 <= Bit_37 ^ Bit_61 ^ Bit_101 ^ Bit_169 ^ Bit_203 ^ Bit_282 ^ Bit_335 ^ Bit_439 ^ Bit_536 ^ Bit_617 ^ Bit_773 ^ Bit_849 ^ Bit_882 ^ Bit_944 ^ Bit_979 ^ Bit_1046 ^ Bit_1062 ^ Bit_1112 ^ Bit_1199 ^ Bit_1200;
				Check_49 <= Bit_13 ^ Bit_49 ^ Bit_117 ^ Bit_178 ^ Bit_240 ^ Bit_283 ^ Bit_383 ^ Bit_389 ^ Bit_486 ^ Bit_722 ^ Bit_770 ^ Bit_818 ^ Bit_907 ^ Bit_948 ^ Bit_982 ^ Bit_1021 ^ Bit_1095 ^ Bit_1106 ^ Bit_1200 ^ Bit_1201;
				Check_50 <= Bit_22 ^ Bit_71 ^ Bit_127 ^ Bit_175 ^ Bit_204 ^ Bit_273 ^ Bit_324 ^ Bit_431 ^ Bit_520 ^ Bit_632 ^ Bit_693 ^ Bit_861 ^ Bit_903 ^ Bit_918 ^ Bit_997 ^ Bit_1029 ^ Bit_1096 ^ Bit_1127 ^ Bit_1201 ^ Bit_1202;
				Check_51 <= Bit_17 ^ Bit_92 ^ Bit_109 ^ Bit_191 ^ Bit_209 ^ Bit_276 ^ Bit_373 ^ Bit_428 ^ Bit_539 ^ Bit_596 ^ Bit_672 ^ Bit_728 ^ Bit_907 ^ Bit_951 ^ Bit_976 ^ Bit_1036 ^ Bit_1066 ^ Bit_1111 ^ Bit_1202 ^ Bit_1203;
				Check_52 <= Bit_36 ^ Bit_95 ^ Bit_134 ^ Bit_190 ^ Bit_207 ^ Bit_261 ^ Bit_437 ^ Bit_525 ^ Bit_561 ^ Bit_623 ^ Bit_648 ^ Bit_694 ^ Bit_911 ^ Bit_935 ^ Bit_971 ^ Bit_1049 ^ Bit_1076 ^ Bit_1140 ^ Bit_1203 ^ Bit_1204;
				Check_53 <= Bit_7 ^ Bit_65 ^ Bit_100 ^ Bit_171 ^ Bit_235 ^ Bit_253 ^ Bit_302 ^ Bit_369 ^ Bit_448 ^ Bit_682 ^ Bit_746 ^ Bit_800 ^ Bit_878 ^ Bit_926 ^ Bit_969 ^ Bit_1021 ^ Bit_1070 ^ Bit_1118 ^ Bit_1204 ^ Bit_1205;
				Check_54 <= Bit_38 ^ Bit_62 ^ Bit_102 ^ Bit_170 ^ Bit_204 ^ Bit_283 ^ Bit_336 ^ Bit_440 ^ Bit_537 ^ Bit_618 ^ Bit_774 ^ Bit_850 ^ Bit_883 ^ Bit_945 ^ Bit_980 ^ Bit_1047 ^ Bit_1063 ^ Bit_1113 ^ Bit_1205 ^ Bit_1206;
				Check_55 <= Bit_14 ^ Bit_50 ^ Bit_118 ^ Bit_179 ^ Bit_193 ^ Bit_284 ^ Bit_384 ^ Bit_390 ^ Bit_487 ^ Bit_723 ^ Bit_771 ^ Bit_819 ^ Bit_908 ^ Bit_949 ^ Bit_983 ^ Bit_1022 ^ Bit_1096 ^ Bit_1107 ^ Bit_1206 ^ Bit_1207;
				Check_56 <= Bit_23 ^ Bit_72 ^ Bit_128 ^ Bit_176 ^ Bit_205 ^ Bit_274 ^ Bit_325 ^ Bit_432 ^ Bit_521 ^ Bit_633 ^ Bit_694 ^ Bit_862 ^ Bit_904 ^ Bit_919 ^ Bit_998 ^ Bit_1030 ^ Bit_1097 ^ Bit_1128 ^ Bit_1207 ^ Bit_1208;
				Check_57 <= Bit_18 ^ Bit_93 ^ Bit_110 ^ Bit_192 ^ Bit_210 ^ Bit_277 ^ Bit_374 ^ Bit_429 ^ Bit_540 ^ Bit_597 ^ Bit_625 ^ Bit_729 ^ Bit_908 ^ Bit_952 ^ Bit_977 ^ Bit_1037 ^ Bit_1067 ^ Bit_1112 ^ Bit_1208 ^ Bit_1209;
				Check_58 <= Bit_37 ^ Bit_96 ^ Bit_135 ^ Bit_191 ^ Bit_208 ^ Bit_262 ^ Bit_438 ^ Bit_526 ^ Bit_562 ^ Bit_624 ^ Bit_649 ^ Bit_695 ^ Bit_912 ^ Bit_936 ^ Bit_972 ^ Bit_1050 ^ Bit_1077 ^ Bit_1141 ^ Bit_1209 ^ Bit_1210;
				Check_59 <= Bit_8 ^ Bit_66 ^ Bit_101 ^ Bit_172 ^ Bit_236 ^ Bit_254 ^ Bit_303 ^ Bit_370 ^ Bit_449 ^ Bit_683 ^ Bit_747 ^ Bit_801 ^ Bit_879 ^ Bit_927 ^ Bit_970 ^ Bit_1022 ^ Bit_1071 ^ Bit_1119 ^ Bit_1210 ^ Bit_1211;
				Check_60 <= Bit_39 ^ Bit_63 ^ Bit_103 ^ Bit_171 ^ Bit_205 ^ Bit_284 ^ Bit_289 ^ Bit_441 ^ Bit_538 ^ Bit_619 ^ Bit_775 ^ Bit_851 ^ Bit_884 ^ Bit_946 ^ Bit_981 ^ Bit_1048 ^ Bit_1064 ^ Bit_1114 ^ Bit_1211 ^ Bit_1212;
				Check_61 <= Bit_15 ^ Bit_51 ^ Bit_119 ^ Bit_180 ^ Bit_194 ^ Bit_285 ^ Bit_337 ^ Bit_391 ^ Bit_488 ^ Bit_724 ^ Bit_772 ^ Bit_820 ^ Bit_909 ^ Bit_950 ^ Bit_984 ^ Bit_1023 ^ Bit_1097 ^ Bit_1108 ^ Bit_1212 ^ Bit_1213;
				Check_62 <= Bit_24 ^ Bit_73 ^ Bit_129 ^ Bit_177 ^ Bit_206 ^ Bit_275 ^ Bit_326 ^ Bit_385 ^ Bit_522 ^ Bit_634 ^ Bit_695 ^ Bit_863 ^ Bit_905 ^ Bit_920 ^ Bit_999 ^ Bit_1031 ^ Bit_1098 ^ Bit_1129 ^ Bit_1213 ^ Bit_1214;
				Check_63 <= Bit_19 ^ Bit_94 ^ Bit_111 ^ Bit_145 ^ Bit_211 ^ Bit_278 ^ Bit_375 ^ Bit_430 ^ Bit_541 ^ Bit_598 ^ Bit_626 ^ Bit_730 ^ Bit_909 ^ Bit_953 ^ Bit_978 ^ Bit_1038 ^ Bit_1068 ^ Bit_1113 ^ Bit_1214 ^ Bit_1215;
				Check_64 <= Bit_38 ^ Bit_49 ^ Bit_136 ^ Bit_192 ^ Bit_209 ^ Bit_263 ^ Bit_439 ^ Bit_527 ^ Bit_563 ^ Bit_577 ^ Bit_650 ^ Bit_696 ^ Bit_865 ^ Bit_937 ^ Bit_973 ^ Bit_1051 ^ Bit_1078 ^ Bit_1142 ^ Bit_1215 ^ Bit_1216;
				Check_65 <= Bit_9 ^ Bit_67 ^ Bit_102 ^ Bit_173 ^ Bit_237 ^ Bit_255 ^ Bit_304 ^ Bit_371 ^ Bit_450 ^ Bit_684 ^ Bit_748 ^ Bit_802 ^ Bit_880 ^ Bit_928 ^ Bit_971 ^ Bit_1023 ^ Bit_1072 ^ Bit_1120 ^ Bit_1216 ^ Bit_1217;
				Check_66 <= Bit_40 ^ Bit_64 ^ Bit_104 ^ Bit_172 ^ Bit_206 ^ Bit_285 ^ Bit_290 ^ Bit_442 ^ Bit_539 ^ Bit_620 ^ Bit_776 ^ Bit_852 ^ Bit_885 ^ Bit_947 ^ Bit_982 ^ Bit_1049 ^ Bit_1065 ^ Bit_1115 ^ Bit_1217 ^ Bit_1218;
				Check_67 <= Bit_16 ^ Bit_52 ^ Bit_120 ^ Bit_181 ^ Bit_195 ^ Bit_286 ^ Bit_338 ^ Bit_392 ^ Bit_489 ^ Bit_725 ^ Bit_773 ^ Bit_821 ^ Bit_910 ^ Bit_951 ^ Bit_985 ^ Bit_1024 ^ Bit_1098 ^ Bit_1109 ^ Bit_1218 ^ Bit_1219;
				Check_68 <= Bit_25 ^ Bit_74 ^ Bit_130 ^ Bit_178 ^ Bit_207 ^ Bit_276 ^ Bit_327 ^ Bit_386 ^ Bit_523 ^ Bit_635 ^ Bit_696 ^ Bit_864 ^ Bit_906 ^ Bit_921 ^ Bit_1000 ^ Bit_1032 ^ Bit_1099 ^ Bit_1130 ^ Bit_1219 ^ Bit_1220;
				Check_69 <= Bit_20 ^ Bit_95 ^ Bit_112 ^ Bit_146 ^ Bit_212 ^ Bit_279 ^ Bit_376 ^ Bit_431 ^ Bit_542 ^ Bit_599 ^ Bit_627 ^ Bit_731 ^ Bit_910 ^ Bit_954 ^ Bit_979 ^ Bit_1039 ^ Bit_1069 ^ Bit_1114 ^ Bit_1220 ^ Bit_1221;
				Check_70 <= Bit_39 ^ Bit_50 ^ Bit_137 ^ Bit_145 ^ Bit_210 ^ Bit_264 ^ Bit_440 ^ Bit_528 ^ Bit_564 ^ Bit_578 ^ Bit_651 ^ Bit_697 ^ Bit_866 ^ Bit_938 ^ Bit_974 ^ Bit_1052 ^ Bit_1079 ^ Bit_1143 ^ Bit_1221 ^ Bit_1222;
				Check_71 <= Bit_10 ^ Bit_68 ^ Bit_103 ^ Bit_174 ^ Bit_238 ^ Bit_256 ^ Bit_305 ^ Bit_372 ^ Bit_451 ^ Bit_685 ^ Bit_749 ^ Bit_803 ^ Bit_881 ^ Bit_929 ^ Bit_972 ^ Bit_1024 ^ Bit_1073 ^ Bit_1121 ^ Bit_1222 ^ Bit_1223;
				Check_72 <= Bit_41 ^ Bit_65 ^ Bit_105 ^ Bit_173 ^ Bit_207 ^ Bit_286 ^ Bit_291 ^ Bit_443 ^ Bit_540 ^ Bit_621 ^ Bit_777 ^ Bit_853 ^ Bit_886 ^ Bit_948 ^ Bit_983 ^ Bit_1050 ^ Bit_1066 ^ Bit_1116 ^ Bit_1223 ^ Bit_1224;
				Check_73 <= Bit_17 ^ Bit_53 ^ Bit_121 ^ Bit_182 ^ Bit_196 ^ Bit_287 ^ Bit_339 ^ Bit_393 ^ Bit_490 ^ Bit_726 ^ Bit_774 ^ Bit_822 ^ Bit_911 ^ Bit_952 ^ Bit_986 ^ Bit_1025 ^ Bit_1099 ^ Bit_1110 ^ Bit_1224 ^ Bit_1225;
				Check_74 <= Bit_26 ^ Bit_75 ^ Bit_131 ^ Bit_179 ^ Bit_208 ^ Bit_277 ^ Bit_328 ^ Bit_387 ^ Bit_524 ^ Bit_636 ^ Bit_697 ^ Bit_817 ^ Bit_907 ^ Bit_922 ^ Bit_1001 ^ Bit_1033 ^ Bit_1100 ^ Bit_1131 ^ Bit_1225 ^ Bit_1226;
				Check_75 <= Bit_21 ^ Bit_96 ^ Bit_113 ^ Bit_147 ^ Bit_213 ^ Bit_280 ^ Bit_377 ^ Bit_432 ^ Bit_543 ^ Bit_600 ^ Bit_628 ^ Bit_732 ^ Bit_911 ^ Bit_955 ^ Bit_980 ^ Bit_1040 ^ Bit_1070 ^ Bit_1115 ^ Bit_1226 ^ Bit_1227;
				Check_76 <= Bit_40 ^ Bit_51 ^ Bit_138 ^ Bit_146 ^ Bit_211 ^ Bit_265 ^ Bit_441 ^ Bit_481 ^ Bit_565 ^ Bit_579 ^ Bit_652 ^ Bit_698 ^ Bit_867 ^ Bit_939 ^ Bit_975 ^ Bit_1053 ^ Bit_1080 ^ Bit_1144 ^ Bit_1227 ^ Bit_1228;
				Check_77 <= Bit_11 ^ Bit_69 ^ Bit_104 ^ Bit_175 ^ Bit_239 ^ Bit_257 ^ Bit_306 ^ Bit_373 ^ Bit_452 ^ Bit_686 ^ Bit_750 ^ Bit_804 ^ Bit_882 ^ Bit_930 ^ Bit_973 ^ Bit_1025 ^ Bit_1074 ^ Bit_1122 ^ Bit_1228 ^ Bit_1229;
				Check_78 <= Bit_42 ^ Bit_66 ^ Bit_106 ^ Bit_174 ^ Bit_208 ^ Bit_287 ^ Bit_292 ^ Bit_444 ^ Bit_541 ^ Bit_622 ^ Bit_778 ^ Bit_854 ^ Bit_887 ^ Bit_949 ^ Bit_984 ^ Bit_1051 ^ Bit_1067 ^ Bit_1117 ^ Bit_1229 ^ Bit_1230;
				Check_79 <= Bit_18 ^ Bit_54 ^ Bit_122 ^ Bit_183 ^ Bit_197 ^ Bit_288 ^ Bit_340 ^ Bit_394 ^ Bit_491 ^ Bit_727 ^ Bit_775 ^ Bit_823 ^ Bit_912 ^ Bit_953 ^ Bit_987 ^ Bit_1026 ^ Bit_1100 ^ Bit_1111 ^ Bit_1230 ^ Bit_1231;
				Check_80 <= Bit_27 ^ Bit_76 ^ Bit_132 ^ Bit_180 ^ Bit_209 ^ Bit_278 ^ Bit_329 ^ Bit_388 ^ Bit_525 ^ Bit_637 ^ Bit_698 ^ Bit_818 ^ Bit_908 ^ Bit_923 ^ Bit_1002 ^ Bit_1034 ^ Bit_1101 ^ Bit_1132 ^ Bit_1231 ^ Bit_1232;
				Check_81 <= Bit_22 ^ Bit_49 ^ Bit_114 ^ Bit_148 ^ Bit_214 ^ Bit_281 ^ Bit_378 ^ Bit_385 ^ Bit_544 ^ Bit_601 ^ Bit_629 ^ Bit_733 ^ Bit_912 ^ Bit_956 ^ Bit_981 ^ Bit_1041 ^ Bit_1071 ^ Bit_1116 ^ Bit_1232 ^ Bit_1233;
				Check_82 <= Bit_41 ^ Bit_52 ^ Bit_139 ^ Bit_147 ^ Bit_212 ^ Bit_266 ^ Bit_442 ^ Bit_482 ^ Bit_566 ^ Bit_580 ^ Bit_653 ^ Bit_699 ^ Bit_868 ^ Bit_940 ^ Bit_976 ^ Bit_1054 ^ Bit_1081 ^ Bit_1145 ^ Bit_1233 ^ Bit_1234;
				Check_83 <= Bit_12 ^ Bit_70 ^ Bit_105 ^ Bit_176 ^ Bit_240 ^ Bit_258 ^ Bit_307 ^ Bit_374 ^ Bit_453 ^ Bit_687 ^ Bit_751 ^ Bit_805 ^ Bit_883 ^ Bit_931 ^ Bit_974 ^ Bit_1026 ^ Bit_1075 ^ Bit_1123 ^ Bit_1234 ^ Bit_1235;
				Check_84 <= Bit_43 ^ Bit_67 ^ Bit_107 ^ Bit_175 ^ Bit_209 ^ Bit_288 ^ Bit_293 ^ Bit_445 ^ Bit_542 ^ Bit_623 ^ Bit_779 ^ Bit_855 ^ Bit_888 ^ Bit_950 ^ Bit_985 ^ Bit_1052 ^ Bit_1068 ^ Bit_1118 ^ Bit_1235 ^ Bit_1236;
				Check_85 <= Bit_19 ^ Bit_55 ^ Bit_123 ^ Bit_184 ^ Bit_198 ^ Bit_241 ^ Bit_341 ^ Bit_395 ^ Bit_492 ^ Bit_728 ^ Bit_776 ^ Bit_824 ^ Bit_865 ^ Bit_954 ^ Bit_988 ^ Bit_1027 ^ Bit_1101 ^ Bit_1112 ^ Bit_1236 ^ Bit_1237;
				Check_86 <= Bit_28 ^ Bit_77 ^ Bit_133 ^ Bit_181 ^ Bit_210 ^ Bit_279 ^ Bit_330 ^ Bit_389 ^ Bit_526 ^ Bit_638 ^ Bit_699 ^ Bit_819 ^ Bit_909 ^ Bit_924 ^ Bit_1003 ^ Bit_1035 ^ Bit_1102 ^ Bit_1133 ^ Bit_1237 ^ Bit_1238;
				Check_87 <= Bit_23 ^ Bit_50 ^ Bit_115 ^ Bit_149 ^ Bit_215 ^ Bit_282 ^ Bit_379 ^ Bit_386 ^ Bit_545 ^ Bit_602 ^ Bit_630 ^ Bit_734 ^ Bit_865 ^ Bit_957 ^ Bit_982 ^ Bit_1042 ^ Bit_1072 ^ Bit_1117 ^ Bit_1238 ^ Bit_1239;
				Check_88 <= Bit_42 ^ Bit_53 ^ Bit_140 ^ Bit_148 ^ Bit_213 ^ Bit_267 ^ Bit_443 ^ Bit_483 ^ Bit_567 ^ Bit_581 ^ Bit_654 ^ Bit_700 ^ Bit_869 ^ Bit_941 ^ Bit_977 ^ Bit_1055 ^ Bit_1082 ^ Bit_1146 ^ Bit_1239 ^ Bit_1240;
				Check_89 <= Bit_13 ^ Bit_71 ^ Bit_106 ^ Bit_177 ^ Bit_193 ^ Bit_259 ^ Bit_308 ^ Bit_375 ^ Bit_454 ^ Bit_688 ^ Bit_752 ^ Bit_806 ^ Bit_884 ^ Bit_932 ^ Bit_975 ^ Bit_1027 ^ Bit_1076 ^ Bit_1124 ^ Bit_1240 ^ Bit_1241;
				Check_90 <= Bit_44 ^ Bit_68 ^ Bit_108 ^ Bit_176 ^ Bit_210 ^ Bit_241 ^ Bit_294 ^ Bit_446 ^ Bit_543 ^ Bit_624 ^ Bit_780 ^ Bit_856 ^ Bit_889 ^ Bit_951 ^ Bit_986 ^ Bit_1053 ^ Bit_1069 ^ Bit_1119 ^ Bit_1241 ^ Bit_1242;
				Check_91 <= Bit_20 ^ Bit_56 ^ Bit_124 ^ Bit_185 ^ Bit_199 ^ Bit_242 ^ Bit_342 ^ Bit_396 ^ Bit_493 ^ Bit_729 ^ Bit_777 ^ Bit_825 ^ Bit_866 ^ Bit_955 ^ Bit_989 ^ Bit_1028 ^ Bit_1102 ^ Bit_1113 ^ Bit_1242 ^ Bit_1243;
				Check_92 <= Bit_29 ^ Bit_78 ^ Bit_134 ^ Bit_182 ^ Bit_211 ^ Bit_280 ^ Bit_331 ^ Bit_390 ^ Bit_527 ^ Bit_639 ^ Bit_700 ^ Bit_820 ^ Bit_910 ^ Bit_925 ^ Bit_1004 ^ Bit_1036 ^ Bit_1103 ^ Bit_1134 ^ Bit_1243 ^ Bit_1244;
				Check_93 <= Bit_24 ^ Bit_51 ^ Bit_116 ^ Bit_150 ^ Bit_216 ^ Bit_283 ^ Bit_380 ^ Bit_387 ^ Bit_546 ^ Bit_603 ^ Bit_631 ^ Bit_735 ^ Bit_866 ^ Bit_958 ^ Bit_983 ^ Bit_1043 ^ Bit_1073 ^ Bit_1118 ^ Bit_1244 ^ Bit_1245;
				Check_94 <= Bit_43 ^ Bit_54 ^ Bit_141 ^ Bit_149 ^ Bit_214 ^ Bit_268 ^ Bit_444 ^ Bit_484 ^ Bit_568 ^ Bit_582 ^ Bit_655 ^ Bit_701 ^ Bit_870 ^ Bit_942 ^ Bit_978 ^ Bit_1056 ^ Bit_1083 ^ Bit_1147 ^ Bit_1245 ^ Bit_1246;
				Check_95 <= Bit_14 ^ Bit_72 ^ Bit_107 ^ Bit_178 ^ Bit_194 ^ Bit_260 ^ Bit_309 ^ Bit_376 ^ Bit_455 ^ Bit_689 ^ Bit_753 ^ Bit_807 ^ Bit_885 ^ Bit_933 ^ Bit_976 ^ Bit_1028 ^ Bit_1077 ^ Bit_1125 ^ Bit_1246 ^ Bit_1247;
				Check_96 <= Bit_45 ^ Bit_69 ^ Bit_109 ^ Bit_177 ^ Bit_211 ^ Bit_242 ^ Bit_295 ^ Bit_447 ^ Bit_544 ^ Bit_577 ^ Bit_781 ^ Bit_857 ^ Bit_890 ^ Bit_952 ^ Bit_987 ^ Bit_1054 ^ Bit_1070 ^ Bit_1120 ^ Bit_1247 ^ Bit_1248;
				Check_97 <= Bit_21 ^ Bit_57 ^ Bit_125 ^ Bit_186 ^ Bit_200 ^ Bit_243 ^ Bit_343 ^ Bit_397 ^ Bit_494 ^ Bit_730 ^ Bit_778 ^ Bit_826 ^ Bit_867 ^ Bit_956 ^ Bit_990 ^ Bit_1029 ^ Bit_1103 ^ Bit_1114 ^ Bit_1248 ^ Bit_1249;
				Check_98 <= Bit_30 ^ Bit_79 ^ Bit_135 ^ Bit_183 ^ Bit_212 ^ Bit_281 ^ Bit_332 ^ Bit_391 ^ Bit_528 ^ Bit_640 ^ Bit_701 ^ Bit_821 ^ Bit_911 ^ Bit_926 ^ Bit_1005 ^ Bit_1037 ^ Bit_1104 ^ Bit_1135 ^ Bit_1249 ^ Bit_1250;
				Check_99 <= Bit_25 ^ Bit_52 ^ Bit_117 ^ Bit_151 ^ Bit_217 ^ Bit_284 ^ Bit_381 ^ Bit_388 ^ Bit_547 ^ Bit_604 ^ Bit_632 ^ Bit_736 ^ Bit_867 ^ Bit_959 ^ Bit_984 ^ Bit_1044 ^ Bit_1074 ^ Bit_1119 ^ Bit_1250 ^ Bit_1251;
				Check_100 <= Bit_44 ^ Bit_55 ^ Bit_142 ^ Bit_150 ^ Bit_215 ^ Bit_269 ^ Bit_445 ^ Bit_485 ^ Bit_569 ^ Bit_583 ^ Bit_656 ^ Bit_702 ^ Bit_871 ^ Bit_943 ^ Bit_979 ^ Bit_1009 ^ Bit_1084 ^ Bit_1148 ^ Bit_1251 ^ Bit_1252;
				Check_101 <= Bit_15 ^ Bit_73 ^ Bit_108 ^ Bit_179 ^ Bit_195 ^ Bit_261 ^ Bit_310 ^ Bit_377 ^ Bit_456 ^ Bit_690 ^ Bit_754 ^ Bit_808 ^ Bit_886 ^ Bit_934 ^ Bit_977 ^ Bit_1029 ^ Bit_1078 ^ Bit_1126 ^ Bit_1252 ^ Bit_1253;
				Check_102 <= Bit_46 ^ Bit_70 ^ Bit_110 ^ Bit_178 ^ Bit_212 ^ Bit_243 ^ Bit_296 ^ Bit_448 ^ Bit_545 ^ Bit_578 ^ Bit_782 ^ Bit_858 ^ Bit_891 ^ Bit_953 ^ Bit_988 ^ Bit_1055 ^ Bit_1071 ^ Bit_1121 ^ Bit_1253 ^ Bit_1254;
				Check_103 <= Bit_22 ^ Bit_58 ^ Bit_126 ^ Bit_187 ^ Bit_201 ^ Bit_244 ^ Bit_344 ^ Bit_398 ^ Bit_495 ^ Bit_731 ^ Bit_779 ^ Bit_827 ^ Bit_868 ^ Bit_957 ^ Bit_991 ^ Bit_1030 ^ Bit_1104 ^ Bit_1115 ^ Bit_1254 ^ Bit_1255;
				Check_104 <= Bit_31 ^ Bit_80 ^ Bit_136 ^ Bit_184 ^ Bit_213 ^ Bit_282 ^ Bit_333 ^ Bit_392 ^ Bit_481 ^ Bit_641 ^ Bit_702 ^ Bit_822 ^ Bit_912 ^ Bit_927 ^ Bit_1006 ^ Bit_1038 ^ Bit_1057 ^ Bit_1136 ^ Bit_1255 ^ Bit_1256;
				Check_105 <= Bit_26 ^ Bit_53 ^ Bit_118 ^ Bit_152 ^ Bit_218 ^ Bit_285 ^ Bit_382 ^ Bit_389 ^ Bit_548 ^ Bit_605 ^ Bit_633 ^ Bit_737 ^ Bit_868 ^ Bit_960 ^ Bit_985 ^ Bit_1045 ^ Bit_1075 ^ Bit_1120 ^ Bit_1256 ^ Bit_1257;
				Check_106 <= Bit_45 ^ Bit_56 ^ Bit_143 ^ Bit_151 ^ Bit_216 ^ Bit_270 ^ Bit_446 ^ Bit_486 ^ Bit_570 ^ Bit_584 ^ Bit_657 ^ Bit_703 ^ Bit_872 ^ Bit_944 ^ Bit_980 ^ Bit_1010 ^ Bit_1085 ^ Bit_1149 ^ Bit_1257 ^ Bit_1258;
				Check_107 <= Bit_16 ^ Bit_74 ^ Bit_109 ^ Bit_180 ^ Bit_196 ^ Bit_262 ^ Bit_311 ^ Bit_378 ^ Bit_457 ^ Bit_691 ^ Bit_755 ^ Bit_809 ^ Bit_887 ^ Bit_935 ^ Bit_978 ^ Bit_1030 ^ Bit_1079 ^ Bit_1127 ^ Bit_1258 ^ Bit_1259;
				Check_108 <= Bit_47 ^ Bit_71 ^ Bit_111 ^ Bit_179 ^ Bit_213 ^ Bit_244 ^ Bit_297 ^ Bit_449 ^ Bit_546 ^ Bit_579 ^ Bit_783 ^ Bit_859 ^ Bit_892 ^ Bit_954 ^ Bit_989 ^ Bit_1056 ^ Bit_1072 ^ Bit_1122 ^ Bit_1259 ^ Bit_1260;
				Check_109 <= Bit_23 ^ Bit_59 ^ Bit_127 ^ Bit_188 ^ Bit_202 ^ Bit_245 ^ Bit_345 ^ Bit_399 ^ Bit_496 ^ Bit_732 ^ Bit_780 ^ Bit_828 ^ Bit_869 ^ Bit_958 ^ Bit_992 ^ Bit_1031 ^ Bit_1057 ^ Bit_1116 ^ Bit_1260 ^ Bit_1261;
				Check_110 <= Bit_32 ^ Bit_81 ^ Bit_137 ^ Bit_185 ^ Bit_214 ^ Bit_283 ^ Bit_334 ^ Bit_393 ^ Bit_482 ^ Bit_642 ^ Bit_703 ^ Bit_823 ^ Bit_865 ^ Bit_928 ^ Bit_1007 ^ Bit_1039 ^ Bit_1058 ^ Bit_1137 ^ Bit_1261 ^ Bit_1262;
				Check_111 <= Bit_27 ^ Bit_54 ^ Bit_119 ^ Bit_153 ^ Bit_219 ^ Bit_286 ^ Bit_383 ^ Bit_390 ^ Bit_549 ^ Bit_606 ^ Bit_634 ^ Bit_738 ^ Bit_869 ^ Bit_913 ^ Bit_986 ^ Bit_1046 ^ Bit_1076 ^ Bit_1121 ^ Bit_1262 ^ Bit_1263;
				Check_112 <= Bit_46 ^ Bit_57 ^ Bit_144 ^ Bit_152 ^ Bit_217 ^ Bit_271 ^ Bit_447 ^ Bit_487 ^ Bit_571 ^ Bit_585 ^ Bit_658 ^ Bit_704 ^ Bit_873 ^ Bit_945 ^ Bit_981 ^ Bit_1011 ^ Bit_1086 ^ Bit_1150 ^ Bit_1263 ^ Bit_1264;
				Check_113 <= Bit_17 ^ Bit_75 ^ Bit_110 ^ Bit_181 ^ Bit_197 ^ Bit_263 ^ Bit_312 ^ Bit_379 ^ Bit_458 ^ Bit_692 ^ Bit_756 ^ Bit_810 ^ Bit_888 ^ Bit_936 ^ Bit_979 ^ Bit_1031 ^ Bit_1080 ^ Bit_1128 ^ Bit_1264 ^ Bit_1265;
				Check_114 <= Bit_48 ^ Bit_72 ^ Bit_112 ^ Bit_180 ^ Bit_214 ^ Bit_245 ^ Bit_298 ^ Bit_450 ^ Bit_547 ^ Bit_580 ^ Bit_784 ^ Bit_860 ^ Bit_893 ^ Bit_955 ^ Bit_990 ^ Bit_1009 ^ Bit_1073 ^ Bit_1123 ^ Bit_1265 ^ Bit_1266;
				Check_115 <= Bit_24 ^ Bit_60 ^ Bit_128 ^ Bit_189 ^ Bit_203 ^ Bit_246 ^ Bit_346 ^ Bit_400 ^ Bit_497 ^ Bit_733 ^ Bit_781 ^ Bit_829 ^ Bit_870 ^ Bit_959 ^ Bit_993 ^ Bit_1032 ^ Bit_1058 ^ Bit_1117 ^ Bit_1266 ^ Bit_1267;
				Check_116 <= Bit_33 ^ Bit_82 ^ Bit_138 ^ Bit_186 ^ Bit_215 ^ Bit_284 ^ Bit_335 ^ Bit_394 ^ Bit_483 ^ Bit_643 ^ Bit_704 ^ Bit_824 ^ Bit_866 ^ Bit_929 ^ Bit_1008 ^ Bit_1040 ^ Bit_1059 ^ Bit_1138 ^ Bit_1267 ^ Bit_1268;
				Check_117 <= Bit_28 ^ Bit_55 ^ Bit_120 ^ Bit_154 ^ Bit_220 ^ Bit_287 ^ Bit_384 ^ Bit_391 ^ Bit_550 ^ Bit_607 ^ Bit_635 ^ Bit_739 ^ Bit_870 ^ Bit_914 ^ Bit_987 ^ Bit_1047 ^ Bit_1077 ^ Bit_1122 ^ Bit_1268 ^ Bit_1269;
				Check_118 <= Bit_47 ^ Bit_58 ^ Bit_97 ^ Bit_153 ^ Bit_218 ^ Bit_272 ^ Bit_448 ^ Bit_488 ^ Bit_572 ^ Bit_586 ^ Bit_659 ^ Bit_705 ^ Bit_874 ^ Bit_946 ^ Bit_982 ^ Bit_1012 ^ Bit_1087 ^ Bit_1151 ^ Bit_1269 ^ Bit_1270;
				Check_119 <= Bit_18 ^ Bit_76 ^ Bit_111 ^ Bit_182 ^ Bit_198 ^ Bit_264 ^ Bit_313 ^ Bit_380 ^ Bit_459 ^ Bit_693 ^ Bit_757 ^ Bit_811 ^ Bit_889 ^ Bit_937 ^ Bit_980 ^ Bit_1032 ^ Bit_1081 ^ Bit_1129 ^ Bit_1270 ^ Bit_1271;
				Check_120 <= Bit_1 ^ Bit_73 ^ Bit_113 ^ Bit_181 ^ Bit_215 ^ Bit_246 ^ Bit_299 ^ Bit_451 ^ Bit_548 ^ Bit_581 ^ Bit_785 ^ Bit_861 ^ Bit_894 ^ Bit_956 ^ Bit_991 ^ Bit_1010 ^ Bit_1074 ^ Bit_1124 ^ Bit_1271 ^ Bit_1272;
				Check_121 <= Bit_25 ^ Bit_61 ^ Bit_129 ^ Bit_190 ^ Bit_204 ^ Bit_247 ^ Bit_347 ^ Bit_401 ^ Bit_498 ^ Bit_734 ^ Bit_782 ^ Bit_830 ^ Bit_871 ^ Bit_960 ^ Bit_994 ^ Bit_1033 ^ Bit_1059 ^ Bit_1118 ^ Bit_1272 ^ Bit_1273;
				Check_122 <= Bit_34 ^ Bit_83 ^ Bit_139 ^ Bit_187 ^ Bit_216 ^ Bit_285 ^ Bit_336 ^ Bit_395 ^ Bit_484 ^ Bit_644 ^ Bit_705 ^ Bit_825 ^ Bit_867 ^ Bit_930 ^ Bit_961 ^ Bit_1041 ^ Bit_1060 ^ Bit_1139 ^ Bit_1273 ^ Bit_1274;
				Check_123 <= Bit_29 ^ Bit_56 ^ Bit_121 ^ Bit_155 ^ Bit_221 ^ Bit_288 ^ Bit_337 ^ Bit_392 ^ Bit_551 ^ Bit_608 ^ Bit_636 ^ Bit_740 ^ Bit_871 ^ Bit_915 ^ Bit_988 ^ Bit_1048 ^ Bit_1078 ^ Bit_1123 ^ Bit_1274 ^ Bit_1275;
				Check_124 <= Bit_48 ^ Bit_59 ^ Bit_98 ^ Bit_154 ^ Bit_219 ^ Bit_273 ^ Bit_449 ^ Bit_489 ^ Bit_573 ^ Bit_587 ^ Bit_660 ^ Bit_706 ^ Bit_875 ^ Bit_947 ^ Bit_983 ^ Bit_1013 ^ Bit_1088 ^ Bit_1152 ^ Bit_1275 ^ Bit_1276;
				Check_125 <= Bit_19 ^ Bit_77 ^ Bit_112 ^ Bit_183 ^ Bit_199 ^ Bit_265 ^ Bit_314 ^ Bit_381 ^ Bit_460 ^ Bit_694 ^ Bit_758 ^ Bit_812 ^ Bit_890 ^ Bit_938 ^ Bit_981 ^ Bit_1033 ^ Bit_1082 ^ Bit_1130 ^ Bit_1276 ^ Bit_1277;
				Check_126 <= Bit_2 ^ Bit_74 ^ Bit_114 ^ Bit_182 ^ Bit_216 ^ Bit_247 ^ Bit_300 ^ Bit_452 ^ Bit_549 ^ Bit_582 ^ Bit_786 ^ Bit_862 ^ Bit_895 ^ Bit_957 ^ Bit_992 ^ Bit_1011 ^ Bit_1075 ^ Bit_1125 ^ Bit_1277 ^ Bit_1278;
				Check_127 <= Bit_26 ^ Bit_62 ^ Bit_130 ^ Bit_191 ^ Bit_205 ^ Bit_248 ^ Bit_348 ^ Bit_402 ^ Bit_499 ^ Bit_735 ^ Bit_783 ^ Bit_831 ^ Bit_872 ^ Bit_913 ^ Bit_995 ^ Bit_1034 ^ Bit_1060 ^ Bit_1119 ^ Bit_1278 ^ Bit_1279;
				Check_128 <= Bit_35 ^ Bit_84 ^ Bit_140 ^ Bit_188 ^ Bit_217 ^ Bit_286 ^ Bit_289 ^ Bit_396 ^ Bit_485 ^ Bit_645 ^ Bit_706 ^ Bit_826 ^ Bit_868 ^ Bit_931 ^ Bit_962 ^ Bit_1042 ^ Bit_1061 ^ Bit_1140 ^ Bit_1279 ^ Bit_1280;
				Check_129 <= Bit_30 ^ Bit_57 ^ Bit_122 ^ Bit_156 ^ Bit_222 ^ Bit_241 ^ Bit_338 ^ Bit_393 ^ Bit_552 ^ Bit_609 ^ Bit_637 ^ Bit_741 ^ Bit_872 ^ Bit_916 ^ Bit_989 ^ Bit_1049 ^ Bit_1079 ^ Bit_1124 ^ Bit_1280 ^ Bit_1281;
				Check_130 <= Bit_1 ^ Bit_60 ^ Bit_99 ^ Bit_155 ^ Bit_220 ^ Bit_274 ^ Bit_450 ^ Bit_490 ^ Bit_574 ^ Bit_588 ^ Bit_661 ^ Bit_707 ^ Bit_876 ^ Bit_948 ^ Bit_984 ^ Bit_1014 ^ Bit_1089 ^ Bit_1105 ^ Bit_1281 ^ Bit_1282;
				Check_131 <= Bit_20 ^ Bit_78 ^ Bit_113 ^ Bit_184 ^ Bit_200 ^ Bit_266 ^ Bit_315 ^ Bit_382 ^ Bit_461 ^ Bit_695 ^ Bit_759 ^ Bit_813 ^ Bit_891 ^ Bit_939 ^ Bit_982 ^ Bit_1034 ^ Bit_1083 ^ Bit_1131 ^ Bit_1282 ^ Bit_1283;
				Check_132 <= Bit_3 ^ Bit_75 ^ Bit_115 ^ Bit_183 ^ Bit_217 ^ Bit_248 ^ Bit_301 ^ Bit_453 ^ Bit_550 ^ Bit_583 ^ Bit_787 ^ Bit_863 ^ Bit_896 ^ Bit_958 ^ Bit_993 ^ Bit_1012 ^ Bit_1076 ^ Bit_1126 ^ Bit_1283 ^ Bit_1284;
				Check_133 <= Bit_27 ^ Bit_63 ^ Bit_131 ^ Bit_192 ^ Bit_206 ^ Bit_249 ^ Bit_349 ^ Bit_403 ^ Bit_500 ^ Bit_736 ^ Bit_784 ^ Bit_832 ^ Bit_873 ^ Bit_914 ^ Bit_996 ^ Bit_1035 ^ Bit_1061 ^ Bit_1120 ^ Bit_1284 ^ Bit_1285;
				Check_134 <= Bit_36 ^ Bit_85 ^ Bit_141 ^ Bit_189 ^ Bit_218 ^ Bit_287 ^ Bit_290 ^ Bit_397 ^ Bit_486 ^ Bit_646 ^ Bit_707 ^ Bit_827 ^ Bit_869 ^ Bit_932 ^ Bit_963 ^ Bit_1043 ^ Bit_1062 ^ Bit_1141 ^ Bit_1285 ^ Bit_1286;
				Check_135 <= Bit_31 ^ Bit_58 ^ Bit_123 ^ Bit_157 ^ Bit_223 ^ Bit_242 ^ Bit_339 ^ Bit_394 ^ Bit_553 ^ Bit_610 ^ Bit_638 ^ Bit_742 ^ Bit_873 ^ Bit_917 ^ Bit_990 ^ Bit_1050 ^ Bit_1080 ^ Bit_1125 ^ Bit_1286 ^ Bit_1287;
				Check_136 <= Bit_2 ^ Bit_61 ^ Bit_100 ^ Bit_156 ^ Bit_221 ^ Bit_275 ^ Bit_451 ^ Bit_491 ^ Bit_575 ^ Bit_589 ^ Bit_662 ^ Bit_708 ^ Bit_877 ^ Bit_949 ^ Bit_985 ^ Bit_1015 ^ Bit_1090 ^ Bit_1106 ^ Bit_1287 ^ Bit_1288;
				Check_137 <= Bit_21 ^ Bit_79 ^ Bit_114 ^ Bit_185 ^ Bit_201 ^ Bit_267 ^ Bit_316 ^ Bit_383 ^ Bit_462 ^ Bit_696 ^ Bit_760 ^ Bit_814 ^ Bit_892 ^ Bit_940 ^ Bit_983 ^ Bit_1035 ^ Bit_1084 ^ Bit_1132 ^ Bit_1288 ^ Bit_1289;
				Check_138 <= Bit_4 ^ Bit_76 ^ Bit_116 ^ Bit_184 ^ Bit_218 ^ Bit_249 ^ Bit_302 ^ Bit_454 ^ Bit_551 ^ Bit_584 ^ Bit_788 ^ Bit_864 ^ Bit_897 ^ Bit_959 ^ Bit_994 ^ Bit_1013 ^ Bit_1077 ^ Bit_1127 ^ Bit_1289 ^ Bit_1290;
				Check_139 <= Bit_28 ^ Bit_64 ^ Bit_132 ^ Bit_145 ^ Bit_207 ^ Bit_250 ^ Bit_350 ^ Bit_404 ^ Bit_501 ^ Bit_737 ^ Bit_785 ^ Bit_833 ^ Bit_874 ^ Bit_915 ^ Bit_997 ^ Bit_1036 ^ Bit_1062 ^ Bit_1121 ^ Bit_1290 ^ Bit_1291;
				Check_140 <= Bit_37 ^ Bit_86 ^ Bit_142 ^ Bit_190 ^ Bit_219 ^ Bit_288 ^ Bit_291 ^ Bit_398 ^ Bit_487 ^ Bit_647 ^ Bit_708 ^ Bit_828 ^ Bit_870 ^ Bit_933 ^ Bit_964 ^ Bit_1044 ^ Bit_1063 ^ Bit_1142 ^ Bit_1291 ^ Bit_1292;
				Check_141 <= Bit_32 ^ Bit_59 ^ Bit_124 ^ Bit_158 ^ Bit_224 ^ Bit_243 ^ Bit_340 ^ Bit_395 ^ Bit_554 ^ Bit_611 ^ Bit_639 ^ Bit_743 ^ Bit_874 ^ Bit_918 ^ Bit_991 ^ Bit_1051 ^ Bit_1081 ^ Bit_1126 ^ Bit_1292 ^ Bit_1293;
				Check_142 <= Bit_3 ^ Bit_62 ^ Bit_101 ^ Bit_157 ^ Bit_222 ^ Bit_276 ^ Bit_452 ^ Bit_492 ^ Bit_576 ^ Bit_590 ^ Bit_663 ^ Bit_709 ^ Bit_878 ^ Bit_950 ^ Bit_986 ^ Bit_1016 ^ Bit_1091 ^ Bit_1107 ^ Bit_1293 ^ Bit_1294;
				Check_143 <= Bit_22 ^ Bit_80 ^ Bit_115 ^ Bit_186 ^ Bit_202 ^ Bit_268 ^ Bit_317 ^ Bit_384 ^ Bit_463 ^ Bit_697 ^ Bit_761 ^ Bit_815 ^ Bit_893 ^ Bit_941 ^ Bit_984 ^ Bit_1036 ^ Bit_1085 ^ Bit_1133 ^ Bit_1294 ^ Bit_1295;
				Check_144 <= Bit_5 ^ Bit_77 ^ Bit_117 ^ Bit_185 ^ Bit_219 ^ Bit_250 ^ Bit_303 ^ Bit_455 ^ Bit_552 ^ Bit_585 ^ Bit_789 ^ Bit_817 ^ Bit_898 ^ Bit_960 ^ Bit_995 ^ Bit_1014 ^ Bit_1078 ^ Bit_1128 ^ Bit_1295 ^ Bit_1296;
				Check_145 <= Bit_29 ^ Bit_65 ^ Bit_133 ^ Bit_146 ^ Bit_208 ^ Bit_251 ^ Bit_351 ^ Bit_405 ^ Bit_502 ^ Bit_738 ^ Bit_786 ^ Bit_834 ^ Bit_875 ^ Bit_916 ^ Bit_998 ^ Bit_1037 ^ Bit_1063 ^ Bit_1122 ^ Bit_1296 ^ Bit_1297;
				Check_146 <= Bit_38 ^ Bit_87 ^ Bit_143 ^ Bit_191 ^ Bit_220 ^ Bit_241 ^ Bit_292 ^ Bit_399 ^ Bit_488 ^ Bit_648 ^ Bit_709 ^ Bit_829 ^ Bit_871 ^ Bit_934 ^ Bit_965 ^ Bit_1045 ^ Bit_1064 ^ Bit_1143 ^ Bit_1297 ^ Bit_1298;
				Check_147 <= Bit_33 ^ Bit_60 ^ Bit_125 ^ Bit_159 ^ Bit_225 ^ Bit_244 ^ Bit_341 ^ Bit_396 ^ Bit_555 ^ Bit_612 ^ Bit_640 ^ Bit_744 ^ Bit_875 ^ Bit_919 ^ Bit_992 ^ Bit_1052 ^ Bit_1082 ^ Bit_1127 ^ Bit_1298 ^ Bit_1299;
				Check_148 <= Bit_4 ^ Bit_63 ^ Bit_102 ^ Bit_158 ^ Bit_223 ^ Bit_277 ^ Bit_453 ^ Bit_493 ^ Bit_529 ^ Bit_591 ^ Bit_664 ^ Bit_710 ^ Bit_879 ^ Bit_951 ^ Bit_987 ^ Bit_1017 ^ Bit_1092 ^ Bit_1108 ^ Bit_1299 ^ Bit_1300;
				Check_149 <= Bit_23 ^ Bit_81 ^ Bit_116 ^ Bit_187 ^ Bit_203 ^ Bit_269 ^ Bit_318 ^ Bit_337 ^ Bit_464 ^ Bit_698 ^ Bit_762 ^ Bit_816 ^ Bit_894 ^ Bit_942 ^ Bit_985 ^ Bit_1037 ^ Bit_1086 ^ Bit_1134 ^ Bit_1300 ^ Bit_1301;
				Check_150 <= Bit_6 ^ Bit_78 ^ Bit_118 ^ Bit_186 ^ Bit_220 ^ Bit_251 ^ Bit_304 ^ Bit_456 ^ Bit_553 ^ Bit_586 ^ Bit_790 ^ Bit_818 ^ Bit_899 ^ Bit_913 ^ Bit_996 ^ Bit_1015 ^ Bit_1079 ^ Bit_1129 ^ Bit_1301 ^ Bit_1302;
				Check_151 <= Bit_30 ^ Bit_66 ^ Bit_134 ^ Bit_147 ^ Bit_209 ^ Bit_252 ^ Bit_352 ^ Bit_406 ^ Bit_503 ^ Bit_739 ^ Bit_787 ^ Bit_835 ^ Bit_876 ^ Bit_917 ^ Bit_999 ^ Bit_1038 ^ Bit_1064 ^ Bit_1123 ^ Bit_1302 ^ Bit_1303;
				Check_152 <= Bit_39 ^ Bit_88 ^ Bit_144 ^ Bit_192 ^ Bit_221 ^ Bit_242 ^ Bit_293 ^ Bit_400 ^ Bit_489 ^ Bit_649 ^ Bit_710 ^ Bit_830 ^ Bit_872 ^ Bit_935 ^ Bit_966 ^ Bit_1046 ^ Bit_1065 ^ Bit_1144 ^ Bit_1303 ^ Bit_1304;
				Check_153 <= Bit_34 ^ Bit_61 ^ Bit_126 ^ Bit_160 ^ Bit_226 ^ Bit_245 ^ Bit_342 ^ Bit_397 ^ Bit_556 ^ Bit_613 ^ Bit_641 ^ Bit_745 ^ Bit_876 ^ Bit_920 ^ Bit_993 ^ Bit_1053 ^ Bit_1083 ^ Bit_1128 ^ Bit_1304 ^ Bit_1305;
				Check_154 <= Bit_5 ^ Bit_64 ^ Bit_103 ^ Bit_159 ^ Bit_224 ^ Bit_278 ^ Bit_454 ^ Bit_494 ^ Bit_530 ^ Bit_592 ^ Bit_665 ^ Bit_711 ^ Bit_880 ^ Bit_952 ^ Bit_988 ^ Bit_1018 ^ Bit_1093 ^ Bit_1109 ^ Bit_1305 ^ Bit_1306;
				Check_155 <= Bit_24 ^ Bit_82 ^ Bit_117 ^ Bit_188 ^ Bit_204 ^ Bit_270 ^ Bit_319 ^ Bit_338 ^ Bit_465 ^ Bit_699 ^ Bit_763 ^ Bit_769 ^ Bit_895 ^ Bit_943 ^ Bit_986 ^ Bit_1038 ^ Bit_1087 ^ Bit_1135 ^ Bit_1306 ^ Bit_1307;
				Check_156 <= Bit_7 ^ Bit_79 ^ Bit_119 ^ Bit_187 ^ Bit_221 ^ Bit_252 ^ Bit_305 ^ Bit_457 ^ Bit_554 ^ Bit_587 ^ Bit_791 ^ Bit_819 ^ Bit_900 ^ Bit_914 ^ Bit_997 ^ Bit_1016 ^ Bit_1080 ^ Bit_1130 ^ Bit_1307 ^ Bit_1308;
				Check_157 <= Bit_31 ^ Bit_67 ^ Bit_135 ^ Bit_148 ^ Bit_210 ^ Bit_253 ^ Bit_353 ^ Bit_407 ^ Bit_504 ^ Bit_740 ^ Bit_788 ^ Bit_836 ^ Bit_877 ^ Bit_918 ^ Bit_1000 ^ Bit_1039 ^ Bit_1065 ^ Bit_1124 ^ Bit_1308 ^ Bit_1309;
				Check_158 <= Bit_40 ^ Bit_89 ^ Bit_97 ^ Bit_145 ^ Bit_222 ^ Bit_243 ^ Bit_294 ^ Bit_401 ^ Bit_490 ^ Bit_650 ^ Bit_711 ^ Bit_831 ^ Bit_873 ^ Bit_936 ^ Bit_967 ^ Bit_1047 ^ Bit_1066 ^ Bit_1145 ^ Bit_1309 ^ Bit_1310;
				Check_159 <= Bit_35 ^ Bit_62 ^ Bit_127 ^ Bit_161 ^ Bit_227 ^ Bit_246 ^ Bit_343 ^ Bit_398 ^ Bit_557 ^ Bit_614 ^ Bit_642 ^ Bit_746 ^ Bit_877 ^ Bit_921 ^ Bit_994 ^ Bit_1054 ^ Bit_1084 ^ Bit_1129 ^ Bit_1310 ^ Bit_1311;
				Check_160 <= Bit_6 ^ Bit_65 ^ Bit_104 ^ Bit_160 ^ Bit_225 ^ Bit_279 ^ Bit_455 ^ Bit_495 ^ Bit_531 ^ Bit_593 ^ Bit_666 ^ Bit_712 ^ Bit_881 ^ Bit_953 ^ Bit_989 ^ Bit_1019 ^ Bit_1094 ^ Bit_1110 ^ Bit_1311 ^ Bit_1312;
				Check_161 <= Bit_25 ^ Bit_83 ^ Bit_118 ^ Bit_189 ^ Bit_205 ^ Bit_271 ^ Bit_320 ^ Bit_339 ^ Bit_466 ^ Bit_700 ^ Bit_764 ^ Bit_770 ^ Bit_896 ^ Bit_944 ^ Bit_987 ^ Bit_1039 ^ Bit_1088 ^ Bit_1136 ^ Bit_1312 ^ Bit_1313;
				Check_162 <= Bit_8 ^ Bit_80 ^ Bit_120 ^ Bit_188 ^ Bit_222 ^ Bit_253 ^ Bit_306 ^ Bit_458 ^ Bit_555 ^ Bit_588 ^ Bit_792 ^ Bit_820 ^ Bit_901 ^ Bit_915 ^ Bit_998 ^ Bit_1017 ^ Bit_1081 ^ Bit_1131 ^ Bit_1313 ^ Bit_1314;
				Check_163 <= Bit_32 ^ Bit_68 ^ Bit_136 ^ Bit_149 ^ Bit_211 ^ Bit_254 ^ Bit_354 ^ Bit_408 ^ Bit_505 ^ Bit_741 ^ Bit_789 ^ Bit_837 ^ Bit_878 ^ Bit_919 ^ Bit_1001 ^ Bit_1040 ^ Bit_1066 ^ Bit_1125 ^ Bit_1314 ^ Bit_1315;
				Check_164 <= Bit_41 ^ Bit_90 ^ Bit_98 ^ Bit_146 ^ Bit_223 ^ Bit_244 ^ Bit_295 ^ Bit_402 ^ Bit_491 ^ Bit_651 ^ Bit_712 ^ Bit_832 ^ Bit_874 ^ Bit_937 ^ Bit_968 ^ Bit_1048 ^ Bit_1067 ^ Bit_1146 ^ Bit_1315 ^ Bit_1316;
				Check_165 <= Bit_36 ^ Bit_63 ^ Bit_128 ^ Bit_162 ^ Bit_228 ^ Bit_247 ^ Bit_344 ^ Bit_399 ^ Bit_558 ^ Bit_615 ^ Bit_643 ^ Bit_747 ^ Bit_878 ^ Bit_922 ^ Bit_995 ^ Bit_1055 ^ Bit_1085 ^ Bit_1130 ^ Bit_1316 ^ Bit_1317;
				Check_166 <= Bit_7 ^ Bit_66 ^ Bit_105 ^ Bit_161 ^ Bit_226 ^ Bit_280 ^ Bit_456 ^ Bit_496 ^ Bit_532 ^ Bit_594 ^ Bit_667 ^ Bit_713 ^ Bit_882 ^ Bit_954 ^ Bit_990 ^ Bit_1020 ^ Bit_1095 ^ Bit_1111 ^ Bit_1317 ^ Bit_1318;
				Check_167 <= Bit_26 ^ Bit_84 ^ Bit_119 ^ Bit_190 ^ Bit_206 ^ Bit_272 ^ Bit_321 ^ Bit_340 ^ Bit_467 ^ Bit_701 ^ Bit_765 ^ Bit_771 ^ Bit_897 ^ Bit_945 ^ Bit_988 ^ Bit_1040 ^ Bit_1089 ^ Bit_1137 ^ Bit_1318 ^ Bit_1319;
				Check_168 <= Bit_9 ^ Bit_81 ^ Bit_121 ^ Bit_189 ^ Bit_223 ^ Bit_254 ^ Bit_307 ^ Bit_459 ^ Bit_556 ^ Bit_589 ^ Bit_793 ^ Bit_821 ^ Bit_902 ^ Bit_916 ^ Bit_999 ^ Bit_1018 ^ Bit_1082 ^ Bit_1132 ^ Bit_1319 ^ Bit_1320;
				Check_169 <= Bit_33 ^ Bit_69 ^ Bit_137 ^ Bit_150 ^ Bit_212 ^ Bit_255 ^ Bit_355 ^ Bit_409 ^ Bit_506 ^ Bit_742 ^ Bit_790 ^ Bit_838 ^ Bit_879 ^ Bit_920 ^ Bit_1002 ^ Bit_1041 ^ Bit_1067 ^ Bit_1126 ^ Bit_1320 ^ Bit_1321;
				Check_170 <= Bit_42 ^ Bit_91 ^ Bit_99 ^ Bit_147 ^ Bit_224 ^ Bit_245 ^ Bit_296 ^ Bit_403 ^ Bit_492 ^ Bit_652 ^ Bit_713 ^ Bit_833 ^ Bit_875 ^ Bit_938 ^ Bit_969 ^ Bit_1049 ^ Bit_1068 ^ Bit_1147 ^ Bit_1321 ^ Bit_1322;
				Check_171 <= Bit_37 ^ Bit_64 ^ Bit_129 ^ Bit_163 ^ Bit_229 ^ Bit_248 ^ Bit_345 ^ Bit_400 ^ Bit_559 ^ Bit_616 ^ Bit_644 ^ Bit_748 ^ Bit_879 ^ Bit_923 ^ Bit_996 ^ Bit_1056 ^ Bit_1086 ^ Bit_1131 ^ Bit_1322 ^ Bit_1323;
				Check_172 <= Bit_8 ^ Bit_67 ^ Bit_106 ^ Bit_162 ^ Bit_227 ^ Bit_281 ^ Bit_457 ^ Bit_497 ^ Bit_533 ^ Bit_595 ^ Bit_668 ^ Bit_714 ^ Bit_883 ^ Bit_955 ^ Bit_991 ^ Bit_1021 ^ Bit_1096 ^ Bit_1112 ^ Bit_1323 ^ Bit_1324;
				Check_173 <= Bit_27 ^ Bit_85 ^ Bit_120 ^ Bit_191 ^ Bit_207 ^ Bit_273 ^ Bit_322 ^ Bit_341 ^ Bit_468 ^ Bit_702 ^ Bit_766 ^ Bit_772 ^ Bit_898 ^ Bit_946 ^ Bit_989 ^ Bit_1041 ^ Bit_1090 ^ Bit_1138 ^ Bit_1324 ^ Bit_1325;
				Check_174 <= Bit_10 ^ Bit_82 ^ Bit_122 ^ Bit_190 ^ Bit_224 ^ Bit_255 ^ Bit_308 ^ Bit_460 ^ Bit_557 ^ Bit_590 ^ Bit_794 ^ Bit_822 ^ Bit_903 ^ Bit_917 ^ Bit_1000 ^ Bit_1019 ^ Bit_1083 ^ Bit_1133 ^ Bit_1325 ^ Bit_1326;
				Check_175 <= Bit_34 ^ Bit_70 ^ Bit_138 ^ Bit_151 ^ Bit_213 ^ Bit_256 ^ Bit_356 ^ Bit_410 ^ Bit_507 ^ Bit_743 ^ Bit_791 ^ Bit_839 ^ Bit_880 ^ Bit_921 ^ Bit_1003 ^ Bit_1042 ^ Bit_1068 ^ Bit_1127 ^ Bit_1326 ^ Bit_1327;
				Check_176 <= Bit_43 ^ Bit_92 ^ Bit_100 ^ Bit_148 ^ Bit_225 ^ Bit_246 ^ Bit_297 ^ Bit_404 ^ Bit_493 ^ Bit_653 ^ Bit_714 ^ Bit_834 ^ Bit_876 ^ Bit_939 ^ Bit_970 ^ Bit_1050 ^ Bit_1069 ^ Bit_1148 ^ Bit_1327 ^ Bit_1328;
				Check_177 <= Bit_38 ^ Bit_65 ^ Bit_130 ^ Bit_164 ^ Bit_230 ^ Bit_249 ^ Bit_346 ^ Bit_401 ^ Bit_560 ^ Bit_617 ^ Bit_645 ^ Bit_749 ^ Bit_880 ^ Bit_924 ^ Bit_997 ^ Bit_1009 ^ Bit_1087 ^ Bit_1132 ^ Bit_1328 ^ Bit_1329;
				Check_178 <= Bit_9 ^ Bit_68 ^ Bit_107 ^ Bit_163 ^ Bit_228 ^ Bit_282 ^ Bit_458 ^ Bit_498 ^ Bit_534 ^ Bit_596 ^ Bit_669 ^ Bit_715 ^ Bit_884 ^ Bit_956 ^ Bit_992 ^ Bit_1022 ^ Bit_1097 ^ Bit_1113 ^ Bit_1329 ^ Bit_1330;
				Check_179 <= Bit_28 ^ Bit_86 ^ Bit_121 ^ Bit_192 ^ Bit_208 ^ Bit_274 ^ Bit_323 ^ Bit_342 ^ Bit_469 ^ Bit_703 ^ Bit_767 ^ Bit_773 ^ Bit_899 ^ Bit_947 ^ Bit_990 ^ Bit_1042 ^ Bit_1091 ^ Bit_1139 ^ Bit_1330 ^ Bit_1331;
				Check_180 <= Bit_11 ^ Bit_83 ^ Bit_123 ^ Bit_191 ^ Bit_225 ^ Bit_256 ^ Bit_309 ^ Bit_461 ^ Bit_558 ^ Bit_591 ^ Bit_795 ^ Bit_823 ^ Bit_904 ^ Bit_918 ^ Bit_1001 ^ Bit_1020 ^ Bit_1084 ^ Bit_1134 ^ Bit_1331 ^ Bit_1332;
				Check_181 <= Bit_35 ^ Bit_71 ^ Bit_139 ^ Bit_152 ^ Bit_214 ^ Bit_257 ^ Bit_357 ^ Bit_411 ^ Bit_508 ^ Bit_744 ^ Bit_792 ^ Bit_840 ^ Bit_881 ^ Bit_922 ^ Bit_1004 ^ Bit_1043 ^ Bit_1069 ^ Bit_1128 ^ Bit_1332 ^ Bit_1333;
				Check_182 <= Bit_44 ^ Bit_93 ^ Bit_101 ^ Bit_149 ^ Bit_226 ^ Bit_247 ^ Bit_298 ^ Bit_405 ^ Bit_494 ^ Bit_654 ^ Bit_715 ^ Bit_835 ^ Bit_877 ^ Bit_940 ^ Bit_971 ^ Bit_1051 ^ Bit_1070 ^ Bit_1149 ^ Bit_1333 ^ Bit_1334;
				Check_183 <= Bit_39 ^ Bit_66 ^ Bit_131 ^ Bit_165 ^ Bit_231 ^ Bit_250 ^ Bit_347 ^ Bit_402 ^ Bit_561 ^ Bit_618 ^ Bit_646 ^ Bit_750 ^ Bit_881 ^ Bit_925 ^ Bit_998 ^ Bit_1010 ^ Bit_1088 ^ Bit_1133 ^ Bit_1334 ^ Bit_1335;
				Check_184 <= Bit_10 ^ Bit_69 ^ Bit_108 ^ Bit_164 ^ Bit_229 ^ Bit_283 ^ Bit_459 ^ Bit_499 ^ Bit_535 ^ Bit_597 ^ Bit_670 ^ Bit_716 ^ Bit_885 ^ Bit_957 ^ Bit_993 ^ Bit_1023 ^ Bit_1098 ^ Bit_1114 ^ Bit_1335 ^ Bit_1336;
				Check_185 <= Bit_29 ^ Bit_87 ^ Bit_122 ^ Bit_145 ^ Bit_209 ^ Bit_275 ^ Bit_324 ^ Bit_343 ^ Bit_470 ^ Bit_704 ^ Bit_768 ^ Bit_774 ^ Bit_900 ^ Bit_948 ^ Bit_991 ^ Bit_1043 ^ Bit_1092 ^ Bit_1140 ^ Bit_1336 ^ Bit_1337;
				Check_186 <= Bit_12 ^ Bit_84 ^ Bit_124 ^ Bit_192 ^ Bit_226 ^ Bit_257 ^ Bit_310 ^ Bit_462 ^ Bit_559 ^ Bit_592 ^ Bit_796 ^ Bit_824 ^ Bit_905 ^ Bit_919 ^ Bit_1002 ^ Bit_1021 ^ Bit_1085 ^ Bit_1135 ^ Bit_1337 ^ Bit_1338;
				Check_187 <= Bit_36 ^ Bit_72 ^ Bit_140 ^ Bit_153 ^ Bit_215 ^ Bit_258 ^ Bit_358 ^ Bit_412 ^ Bit_509 ^ Bit_745 ^ Bit_793 ^ Bit_841 ^ Bit_882 ^ Bit_923 ^ Bit_1005 ^ Bit_1044 ^ Bit_1070 ^ Bit_1129 ^ Bit_1338 ^ Bit_1339;
				Check_188 <= Bit_45 ^ Bit_94 ^ Bit_102 ^ Bit_150 ^ Bit_227 ^ Bit_248 ^ Bit_299 ^ Bit_406 ^ Bit_495 ^ Bit_655 ^ Bit_716 ^ Bit_836 ^ Bit_878 ^ Bit_941 ^ Bit_972 ^ Bit_1052 ^ Bit_1071 ^ Bit_1150 ^ Bit_1339 ^ Bit_1340;
				Check_189 <= Bit_40 ^ Bit_67 ^ Bit_132 ^ Bit_166 ^ Bit_232 ^ Bit_251 ^ Bit_348 ^ Bit_403 ^ Bit_562 ^ Bit_619 ^ Bit_647 ^ Bit_751 ^ Bit_882 ^ Bit_926 ^ Bit_999 ^ Bit_1011 ^ Bit_1089 ^ Bit_1134 ^ Bit_1340 ^ Bit_1341;
				Check_190 <= Bit_11 ^ Bit_70 ^ Bit_109 ^ Bit_165 ^ Bit_230 ^ Bit_284 ^ Bit_460 ^ Bit_500 ^ Bit_536 ^ Bit_598 ^ Bit_671 ^ Bit_717 ^ Bit_886 ^ Bit_958 ^ Bit_994 ^ Bit_1024 ^ Bit_1099 ^ Bit_1115 ^ Bit_1341 ^ Bit_1342;
				Check_191 <= Bit_30 ^ Bit_88 ^ Bit_123 ^ Bit_146 ^ Bit_210 ^ Bit_276 ^ Bit_325 ^ Bit_344 ^ Bit_471 ^ Bit_705 ^ Bit_721 ^ Bit_775 ^ Bit_901 ^ Bit_949 ^ Bit_992 ^ Bit_1044 ^ Bit_1093 ^ Bit_1141 ^ Bit_1342 ^ Bit_1343;
				Check_192 <= Bit_13 ^ Bit_85 ^ Bit_125 ^ Bit_145 ^ Bit_227 ^ Bit_258 ^ Bit_311 ^ Bit_463 ^ Bit_560 ^ Bit_593 ^ Bit_797 ^ Bit_825 ^ Bit_906 ^ Bit_920 ^ Bit_1003 ^ Bit_1022 ^ Bit_1086 ^ Bit_1136 ^ Bit_1343 ^ Bit_1344;
				Check_193 <= Bit_37 ^ Bit_73 ^ Bit_141 ^ Bit_154 ^ Bit_216 ^ Bit_259 ^ Bit_359 ^ Bit_413 ^ Bit_510 ^ Bit_746 ^ Bit_794 ^ Bit_842 ^ Bit_883 ^ Bit_924 ^ Bit_1006 ^ Bit_1045 ^ Bit_1071 ^ Bit_1130 ^ Bit_1344 ^ Bit_1345;
				Check_194 <= Bit_46 ^ Bit_95 ^ Bit_103 ^ Bit_151 ^ Bit_228 ^ Bit_249 ^ Bit_300 ^ Bit_407 ^ Bit_496 ^ Bit_656 ^ Bit_717 ^ Bit_837 ^ Bit_879 ^ Bit_942 ^ Bit_973 ^ Bit_1053 ^ Bit_1072 ^ Bit_1151 ^ Bit_1345 ^ Bit_1346;
				Check_195 <= Bit_41 ^ Bit_68 ^ Bit_133 ^ Bit_167 ^ Bit_233 ^ Bit_252 ^ Bit_349 ^ Bit_404 ^ Bit_563 ^ Bit_620 ^ Bit_648 ^ Bit_752 ^ Bit_883 ^ Bit_927 ^ Bit_1000 ^ Bit_1012 ^ Bit_1090 ^ Bit_1135 ^ Bit_1346 ^ Bit_1347;
				Check_196 <= Bit_12 ^ Bit_71 ^ Bit_110 ^ Bit_166 ^ Bit_231 ^ Bit_285 ^ Bit_461 ^ Bit_501 ^ Bit_537 ^ Bit_599 ^ Bit_672 ^ Bit_718 ^ Bit_887 ^ Bit_959 ^ Bit_995 ^ Bit_1025 ^ Bit_1100 ^ Bit_1116 ^ Bit_1347 ^ Bit_1348;
				Check_197 <= Bit_31 ^ Bit_89 ^ Bit_124 ^ Bit_147 ^ Bit_211 ^ Bit_277 ^ Bit_326 ^ Bit_345 ^ Bit_472 ^ Bit_706 ^ Bit_722 ^ Bit_776 ^ Bit_902 ^ Bit_950 ^ Bit_993 ^ Bit_1045 ^ Bit_1094 ^ Bit_1142 ^ Bit_1348 ^ Bit_1349;
				Check_198 <= Bit_14 ^ Bit_86 ^ Bit_126 ^ Bit_146 ^ Bit_228 ^ Bit_259 ^ Bit_312 ^ Bit_464 ^ Bit_561 ^ Bit_594 ^ Bit_798 ^ Bit_826 ^ Bit_907 ^ Bit_921 ^ Bit_1004 ^ Bit_1023 ^ Bit_1087 ^ Bit_1137 ^ Bit_1349 ^ Bit_1350;
				Check_199 <= Bit_38 ^ Bit_74 ^ Bit_142 ^ Bit_155 ^ Bit_217 ^ Bit_260 ^ Bit_360 ^ Bit_414 ^ Bit_511 ^ Bit_747 ^ Bit_795 ^ Bit_843 ^ Bit_884 ^ Bit_925 ^ Bit_1007 ^ Bit_1046 ^ Bit_1072 ^ Bit_1131 ^ Bit_1350 ^ Bit_1351;
				Check_200 <= Bit_47 ^ Bit_96 ^ Bit_104 ^ Bit_152 ^ Bit_229 ^ Bit_250 ^ Bit_301 ^ Bit_408 ^ Bit_497 ^ Bit_657 ^ Bit_718 ^ Bit_838 ^ Bit_880 ^ Bit_943 ^ Bit_974 ^ Bit_1054 ^ Bit_1073 ^ Bit_1152 ^ Bit_1351 ^ Bit_1352;
				Check_201 <= Bit_42 ^ Bit_69 ^ Bit_134 ^ Bit_168 ^ Bit_234 ^ Bit_253 ^ Bit_350 ^ Bit_405 ^ Bit_564 ^ Bit_621 ^ Bit_649 ^ Bit_753 ^ Bit_884 ^ Bit_928 ^ Bit_1001 ^ Bit_1013 ^ Bit_1091 ^ Bit_1136 ^ Bit_1352 ^ Bit_1353;
				Check_202 <= Bit_13 ^ Bit_72 ^ Bit_111 ^ Bit_167 ^ Bit_232 ^ Bit_286 ^ Bit_462 ^ Bit_502 ^ Bit_538 ^ Bit_600 ^ Bit_625 ^ Bit_719 ^ Bit_888 ^ Bit_960 ^ Bit_996 ^ Bit_1026 ^ Bit_1101 ^ Bit_1117 ^ Bit_1353 ^ Bit_1354;
				Check_203 <= Bit_32 ^ Bit_90 ^ Bit_125 ^ Bit_148 ^ Bit_212 ^ Bit_278 ^ Bit_327 ^ Bit_346 ^ Bit_473 ^ Bit_707 ^ Bit_723 ^ Bit_777 ^ Bit_903 ^ Bit_951 ^ Bit_994 ^ Bit_1046 ^ Bit_1095 ^ Bit_1143 ^ Bit_1354 ^ Bit_1355;
				Check_204 <= Bit_15 ^ Bit_87 ^ Bit_127 ^ Bit_147 ^ Bit_229 ^ Bit_260 ^ Bit_313 ^ Bit_465 ^ Bit_562 ^ Bit_595 ^ Bit_799 ^ Bit_827 ^ Bit_908 ^ Bit_922 ^ Bit_1005 ^ Bit_1024 ^ Bit_1088 ^ Bit_1138 ^ Bit_1355 ^ Bit_1356;
				Check_205 <= Bit_39 ^ Bit_75 ^ Bit_143 ^ Bit_156 ^ Bit_218 ^ Bit_261 ^ Bit_361 ^ Bit_415 ^ Bit_512 ^ Bit_748 ^ Bit_796 ^ Bit_844 ^ Bit_885 ^ Bit_926 ^ Bit_1008 ^ Bit_1047 ^ Bit_1073 ^ Bit_1132 ^ Bit_1356 ^ Bit_1357;
				Check_206 <= Bit_48 ^ Bit_49 ^ Bit_105 ^ Bit_153 ^ Bit_230 ^ Bit_251 ^ Bit_302 ^ Bit_409 ^ Bit_498 ^ Bit_658 ^ Bit_719 ^ Bit_839 ^ Bit_881 ^ Bit_944 ^ Bit_975 ^ Bit_1055 ^ Bit_1074 ^ Bit_1105 ^ Bit_1357 ^ Bit_1358;
				Check_207 <= Bit_43 ^ Bit_70 ^ Bit_135 ^ Bit_169 ^ Bit_235 ^ Bit_254 ^ Bit_351 ^ Bit_406 ^ Bit_565 ^ Bit_622 ^ Bit_650 ^ Bit_754 ^ Bit_885 ^ Bit_929 ^ Bit_1002 ^ Bit_1014 ^ Bit_1092 ^ Bit_1137 ^ Bit_1358 ^ Bit_1359;
				Check_208 <= Bit_14 ^ Bit_73 ^ Bit_112 ^ Bit_168 ^ Bit_233 ^ Bit_287 ^ Bit_463 ^ Bit_503 ^ Bit_539 ^ Bit_601 ^ Bit_626 ^ Bit_720 ^ Bit_889 ^ Bit_913 ^ Bit_997 ^ Bit_1027 ^ Bit_1102 ^ Bit_1118 ^ Bit_1359 ^ Bit_1360;
				Check_209 <= Bit_33 ^ Bit_91 ^ Bit_126 ^ Bit_149 ^ Bit_213 ^ Bit_279 ^ Bit_328 ^ Bit_347 ^ Bit_474 ^ Bit_708 ^ Bit_724 ^ Bit_778 ^ Bit_904 ^ Bit_952 ^ Bit_995 ^ Bit_1047 ^ Bit_1096 ^ Bit_1144 ^ Bit_1360 ^ Bit_1361;
				Check_210 <= Bit_16 ^ Bit_88 ^ Bit_128 ^ Bit_148 ^ Bit_230 ^ Bit_261 ^ Bit_314 ^ Bit_466 ^ Bit_563 ^ Bit_596 ^ Bit_800 ^ Bit_828 ^ Bit_909 ^ Bit_923 ^ Bit_1006 ^ Bit_1025 ^ Bit_1089 ^ Bit_1139 ^ Bit_1361 ^ Bit_1362;
				Check_211 <= Bit_40 ^ Bit_76 ^ Bit_144 ^ Bit_157 ^ Bit_219 ^ Bit_262 ^ Bit_362 ^ Bit_416 ^ Bit_513 ^ Bit_749 ^ Bit_797 ^ Bit_845 ^ Bit_886 ^ Bit_927 ^ Bit_961 ^ Bit_1048 ^ Bit_1074 ^ Bit_1133 ^ Bit_1362 ^ Bit_1363;
				Check_212 <= Bit_1 ^ Bit_50 ^ Bit_106 ^ Bit_154 ^ Bit_231 ^ Bit_252 ^ Bit_303 ^ Bit_410 ^ Bit_499 ^ Bit_659 ^ Bit_720 ^ Bit_840 ^ Bit_882 ^ Bit_945 ^ Bit_976 ^ Bit_1056 ^ Bit_1075 ^ Bit_1106 ^ Bit_1363 ^ Bit_1364;
				Check_213 <= Bit_44 ^ Bit_71 ^ Bit_136 ^ Bit_170 ^ Bit_236 ^ Bit_255 ^ Bit_352 ^ Bit_407 ^ Bit_566 ^ Bit_623 ^ Bit_651 ^ Bit_755 ^ Bit_886 ^ Bit_930 ^ Bit_1003 ^ Bit_1015 ^ Bit_1093 ^ Bit_1138 ^ Bit_1364 ^ Bit_1365;
				Check_214 <= Bit_15 ^ Bit_74 ^ Bit_113 ^ Bit_169 ^ Bit_234 ^ Bit_288 ^ Bit_464 ^ Bit_504 ^ Bit_540 ^ Bit_602 ^ Bit_627 ^ Bit_673 ^ Bit_890 ^ Bit_914 ^ Bit_998 ^ Bit_1028 ^ Bit_1103 ^ Bit_1119 ^ Bit_1365 ^ Bit_1366;
				Check_215 <= Bit_34 ^ Bit_92 ^ Bit_127 ^ Bit_150 ^ Bit_214 ^ Bit_280 ^ Bit_329 ^ Bit_348 ^ Bit_475 ^ Bit_709 ^ Bit_725 ^ Bit_779 ^ Bit_905 ^ Bit_953 ^ Bit_996 ^ Bit_1048 ^ Bit_1097 ^ Bit_1145 ^ Bit_1366 ^ Bit_1367;
				Check_216 <= Bit_17 ^ Bit_89 ^ Bit_129 ^ Bit_149 ^ Bit_231 ^ Bit_262 ^ Bit_315 ^ Bit_467 ^ Bit_564 ^ Bit_597 ^ Bit_801 ^ Bit_829 ^ Bit_910 ^ Bit_924 ^ Bit_1007 ^ Bit_1026 ^ Bit_1090 ^ Bit_1140 ^ Bit_1367 ^ Bit_1368;
				Check_217 <= Bit_41 ^ Bit_77 ^ Bit_97 ^ Bit_158 ^ Bit_220 ^ Bit_263 ^ Bit_363 ^ Bit_417 ^ Bit_514 ^ Bit_750 ^ Bit_798 ^ Bit_846 ^ Bit_887 ^ Bit_928 ^ Bit_962 ^ Bit_1049 ^ Bit_1075 ^ Bit_1134 ^ Bit_1368 ^ Bit_1369;
				Check_218 <= Bit_2 ^ Bit_51 ^ Bit_107 ^ Bit_155 ^ Bit_232 ^ Bit_253 ^ Bit_304 ^ Bit_411 ^ Bit_500 ^ Bit_660 ^ Bit_673 ^ Bit_841 ^ Bit_883 ^ Bit_946 ^ Bit_977 ^ Bit_1009 ^ Bit_1076 ^ Bit_1107 ^ Bit_1369 ^ Bit_1370;
				Check_219 <= Bit_45 ^ Bit_72 ^ Bit_137 ^ Bit_171 ^ Bit_237 ^ Bit_256 ^ Bit_353 ^ Bit_408 ^ Bit_567 ^ Bit_624 ^ Bit_652 ^ Bit_756 ^ Bit_887 ^ Bit_931 ^ Bit_1004 ^ Bit_1016 ^ Bit_1094 ^ Bit_1139 ^ Bit_1370 ^ Bit_1371;
				Check_220 <= Bit_16 ^ Bit_75 ^ Bit_114 ^ Bit_170 ^ Bit_235 ^ Bit_241 ^ Bit_465 ^ Bit_505 ^ Bit_541 ^ Bit_603 ^ Bit_628 ^ Bit_674 ^ Bit_891 ^ Bit_915 ^ Bit_999 ^ Bit_1029 ^ Bit_1104 ^ Bit_1120 ^ Bit_1371 ^ Bit_1372;
				Check_221 <= Bit_35 ^ Bit_93 ^ Bit_128 ^ Bit_151 ^ Bit_215 ^ Bit_281 ^ Bit_330 ^ Bit_349 ^ Bit_476 ^ Bit_710 ^ Bit_726 ^ Bit_780 ^ Bit_906 ^ Bit_954 ^ Bit_997 ^ Bit_1049 ^ Bit_1098 ^ Bit_1146 ^ Bit_1372 ^ Bit_1373;
				Check_222 <= Bit_18 ^ Bit_90 ^ Bit_130 ^ Bit_150 ^ Bit_232 ^ Bit_263 ^ Bit_316 ^ Bit_468 ^ Bit_565 ^ Bit_598 ^ Bit_802 ^ Bit_830 ^ Bit_911 ^ Bit_925 ^ Bit_1008 ^ Bit_1027 ^ Bit_1091 ^ Bit_1141 ^ Bit_1373 ^ Bit_1374;
				Check_223 <= Bit_42 ^ Bit_78 ^ Bit_98 ^ Bit_159 ^ Bit_221 ^ Bit_264 ^ Bit_364 ^ Bit_418 ^ Bit_515 ^ Bit_751 ^ Bit_799 ^ Bit_847 ^ Bit_888 ^ Bit_929 ^ Bit_963 ^ Bit_1050 ^ Bit_1076 ^ Bit_1135 ^ Bit_1374 ^ Bit_1375;
				Check_224 <= Bit_3 ^ Bit_52 ^ Bit_108 ^ Bit_156 ^ Bit_233 ^ Bit_254 ^ Bit_305 ^ Bit_412 ^ Bit_501 ^ Bit_661 ^ Bit_674 ^ Bit_842 ^ Bit_884 ^ Bit_947 ^ Bit_978 ^ Bit_1010 ^ Bit_1077 ^ Bit_1108 ^ Bit_1375 ^ Bit_1376;
				Check_225 <= Bit_46 ^ Bit_73 ^ Bit_138 ^ Bit_172 ^ Bit_238 ^ Bit_257 ^ Bit_354 ^ Bit_409 ^ Bit_568 ^ Bit_577 ^ Bit_653 ^ Bit_757 ^ Bit_888 ^ Bit_932 ^ Bit_1005 ^ Bit_1017 ^ Bit_1095 ^ Bit_1140 ^ Bit_1376 ^ Bit_1377;
				Check_226 <= Bit_17 ^ Bit_76 ^ Bit_115 ^ Bit_171 ^ Bit_236 ^ Bit_242 ^ Bit_466 ^ Bit_506 ^ Bit_542 ^ Bit_604 ^ Bit_629 ^ Bit_675 ^ Bit_892 ^ Bit_916 ^ Bit_1000 ^ Bit_1030 ^ Bit_1057 ^ Bit_1121 ^ Bit_1377 ^ Bit_1378;
				Check_227 <= Bit_36 ^ Bit_94 ^ Bit_129 ^ Bit_152 ^ Bit_216 ^ Bit_282 ^ Bit_331 ^ Bit_350 ^ Bit_477 ^ Bit_711 ^ Bit_727 ^ Bit_781 ^ Bit_907 ^ Bit_955 ^ Bit_998 ^ Bit_1050 ^ Bit_1099 ^ Bit_1147 ^ Bit_1378 ^ Bit_1379;
				Check_228 <= Bit_19 ^ Bit_91 ^ Bit_131 ^ Bit_151 ^ Bit_233 ^ Bit_264 ^ Bit_317 ^ Bit_469 ^ Bit_566 ^ Bit_599 ^ Bit_803 ^ Bit_831 ^ Bit_912 ^ Bit_926 ^ Bit_961 ^ Bit_1028 ^ Bit_1092 ^ Bit_1142 ^ Bit_1379 ^ Bit_1380;
				Check_229 <= Bit_43 ^ Bit_79 ^ Bit_99 ^ Bit_160 ^ Bit_222 ^ Bit_265 ^ Bit_365 ^ Bit_419 ^ Bit_516 ^ Bit_752 ^ Bit_800 ^ Bit_848 ^ Bit_889 ^ Bit_930 ^ Bit_964 ^ Bit_1051 ^ Bit_1077 ^ Bit_1136 ^ Bit_1380 ^ Bit_1381;
				Check_230 <= Bit_4 ^ Bit_53 ^ Bit_109 ^ Bit_157 ^ Bit_234 ^ Bit_255 ^ Bit_306 ^ Bit_413 ^ Bit_502 ^ Bit_662 ^ Bit_675 ^ Bit_843 ^ Bit_885 ^ Bit_948 ^ Bit_979 ^ Bit_1011 ^ Bit_1078 ^ Bit_1109 ^ Bit_1381 ^ Bit_1382;
				Check_231 <= Bit_47 ^ Bit_74 ^ Bit_139 ^ Bit_173 ^ Bit_239 ^ Bit_258 ^ Bit_355 ^ Bit_410 ^ Bit_569 ^ Bit_578 ^ Bit_654 ^ Bit_758 ^ Bit_889 ^ Bit_933 ^ Bit_1006 ^ Bit_1018 ^ Bit_1096 ^ Bit_1141 ^ Bit_1382 ^ Bit_1383;
				Check_232 <= Bit_18 ^ Bit_77 ^ Bit_116 ^ Bit_172 ^ Bit_237 ^ Bit_243 ^ Bit_467 ^ Bit_507 ^ Bit_543 ^ Bit_605 ^ Bit_630 ^ Bit_676 ^ Bit_893 ^ Bit_917 ^ Bit_1001 ^ Bit_1031 ^ Bit_1058 ^ Bit_1122 ^ Bit_1383 ^ Bit_1384;
				Check_233 <= Bit_37 ^ Bit_95 ^ Bit_130 ^ Bit_153 ^ Bit_217 ^ Bit_283 ^ Bit_332 ^ Bit_351 ^ Bit_478 ^ Bit_712 ^ Bit_728 ^ Bit_782 ^ Bit_908 ^ Bit_956 ^ Bit_999 ^ Bit_1051 ^ Bit_1100 ^ Bit_1148 ^ Bit_1384 ^ Bit_1385;
				Check_234 <= Bit_20 ^ Bit_92 ^ Bit_132 ^ Bit_152 ^ Bit_234 ^ Bit_265 ^ Bit_318 ^ Bit_470 ^ Bit_567 ^ Bit_600 ^ Bit_804 ^ Bit_832 ^ Bit_865 ^ Bit_927 ^ Bit_962 ^ Bit_1029 ^ Bit_1093 ^ Bit_1143 ^ Bit_1385 ^ Bit_1386;
				Check_235 <= Bit_44 ^ Bit_80 ^ Bit_100 ^ Bit_161 ^ Bit_223 ^ Bit_266 ^ Bit_366 ^ Bit_420 ^ Bit_517 ^ Bit_753 ^ Bit_801 ^ Bit_849 ^ Bit_890 ^ Bit_931 ^ Bit_965 ^ Bit_1052 ^ Bit_1078 ^ Bit_1137 ^ Bit_1386 ^ Bit_1387;
				Check_236 <= Bit_5 ^ Bit_54 ^ Bit_110 ^ Bit_158 ^ Bit_235 ^ Bit_256 ^ Bit_307 ^ Bit_414 ^ Bit_503 ^ Bit_663 ^ Bit_676 ^ Bit_844 ^ Bit_886 ^ Bit_949 ^ Bit_980 ^ Bit_1012 ^ Bit_1079 ^ Bit_1110 ^ Bit_1387 ^ Bit_1388;
				Check_237 <= Bit_48 ^ Bit_75 ^ Bit_140 ^ Bit_174 ^ Bit_240 ^ Bit_259 ^ Bit_356 ^ Bit_411 ^ Bit_570 ^ Bit_579 ^ Bit_655 ^ Bit_759 ^ Bit_890 ^ Bit_934 ^ Bit_1007 ^ Bit_1019 ^ Bit_1097 ^ Bit_1142 ^ Bit_1388 ^ Bit_1389;
				Check_238 <= Bit_19 ^ Bit_78 ^ Bit_117 ^ Bit_173 ^ Bit_238 ^ Bit_244 ^ Bit_468 ^ Bit_508 ^ Bit_544 ^ Bit_606 ^ Bit_631 ^ Bit_677 ^ Bit_894 ^ Bit_918 ^ Bit_1002 ^ Bit_1032 ^ Bit_1059 ^ Bit_1123 ^ Bit_1389 ^ Bit_1390;
				Check_239 <= Bit_38 ^ Bit_96 ^ Bit_131 ^ Bit_154 ^ Bit_218 ^ Bit_284 ^ Bit_333 ^ Bit_352 ^ Bit_479 ^ Bit_713 ^ Bit_729 ^ Bit_783 ^ Bit_909 ^ Bit_957 ^ Bit_1000 ^ Bit_1052 ^ Bit_1101 ^ Bit_1149 ^ Bit_1390 ^ Bit_1391;
				Check_240 <= Bit_21 ^ Bit_93 ^ Bit_133 ^ Bit_153 ^ Bit_235 ^ Bit_266 ^ Bit_319 ^ Bit_471 ^ Bit_568 ^ Bit_601 ^ Bit_805 ^ Bit_833 ^ Bit_866 ^ Bit_928 ^ Bit_963 ^ Bit_1030 ^ Bit_1094 ^ Bit_1144 ^ Bit_1391 ^ Bit_1392;
				Check_241 <= Bit_45 ^ Bit_81 ^ Bit_101 ^ Bit_162 ^ Bit_224 ^ Bit_267 ^ Bit_367 ^ Bit_421 ^ Bit_518 ^ Bit_754 ^ Bit_802 ^ Bit_850 ^ Bit_891 ^ Bit_932 ^ Bit_966 ^ Bit_1053 ^ Bit_1079 ^ Bit_1138 ^ Bit_1392 ^ Bit_1393;
				Check_242 <= Bit_6 ^ Bit_55 ^ Bit_111 ^ Bit_159 ^ Bit_236 ^ Bit_257 ^ Bit_308 ^ Bit_415 ^ Bit_504 ^ Bit_664 ^ Bit_677 ^ Bit_845 ^ Bit_887 ^ Bit_950 ^ Bit_981 ^ Bit_1013 ^ Bit_1080 ^ Bit_1111 ^ Bit_1393 ^ Bit_1394;
				Check_243 <= Bit_1 ^ Bit_76 ^ Bit_141 ^ Bit_175 ^ Bit_193 ^ Bit_260 ^ Bit_357 ^ Bit_412 ^ Bit_571 ^ Bit_580 ^ Bit_656 ^ Bit_760 ^ Bit_891 ^ Bit_935 ^ Bit_1008 ^ Bit_1020 ^ Bit_1098 ^ Bit_1143 ^ Bit_1394 ^ Bit_1395;
				Check_244 <= Bit_20 ^ Bit_79 ^ Bit_118 ^ Bit_174 ^ Bit_239 ^ Bit_245 ^ Bit_469 ^ Bit_509 ^ Bit_545 ^ Bit_607 ^ Bit_632 ^ Bit_678 ^ Bit_895 ^ Bit_919 ^ Bit_1003 ^ Bit_1033 ^ Bit_1060 ^ Bit_1124 ^ Bit_1395 ^ Bit_1396;
				Check_245 <= Bit_39 ^ Bit_49 ^ Bit_132 ^ Bit_155 ^ Bit_219 ^ Bit_285 ^ Bit_334 ^ Bit_353 ^ Bit_480 ^ Bit_714 ^ Bit_730 ^ Bit_784 ^ Bit_910 ^ Bit_958 ^ Bit_1001 ^ Bit_1053 ^ Bit_1102 ^ Bit_1150 ^ Bit_1396 ^ Bit_1397;
				Check_246 <= Bit_22 ^ Bit_94 ^ Bit_134 ^ Bit_154 ^ Bit_236 ^ Bit_267 ^ Bit_320 ^ Bit_472 ^ Bit_569 ^ Bit_602 ^ Bit_806 ^ Bit_834 ^ Bit_867 ^ Bit_929 ^ Bit_964 ^ Bit_1031 ^ Bit_1095 ^ Bit_1145 ^ Bit_1397 ^ Bit_1398;
				Check_247 <= Bit_46 ^ Bit_82 ^ Bit_102 ^ Bit_163 ^ Bit_225 ^ Bit_268 ^ Bit_368 ^ Bit_422 ^ Bit_519 ^ Bit_755 ^ Bit_803 ^ Bit_851 ^ Bit_892 ^ Bit_933 ^ Bit_967 ^ Bit_1054 ^ Bit_1080 ^ Bit_1139 ^ Bit_1398 ^ Bit_1399;
				Check_248 <= Bit_7 ^ Bit_56 ^ Bit_112 ^ Bit_160 ^ Bit_237 ^ Bit_258 ^ Bit_309 ^ Bit_416 ^ Bit_505 ^ Bit_665 ^ Bit_678 ^ Bit_846 ^ Bit_888 ^ Bit_951 ^ Bit_982 ^ Bit_1014 ^ Bit_1081 ^ Bit_1112 ^ Bit_1399 ^ Bit_1400;
				Check_249 <= Bit_2 ^ Bit_77 ^ Bit_142 ^ Bit_176 ^ Bit_194 ^ Bit_261 ^ Bit_358 ^ Bit_413 ^ Bit_572 ^ Bit_581 ^ Bit_657 ^ Bit_761 ^ Bit_892 ^ Bit_936 ^ Bit_961 ^ Bit_1021 ^ Bit_1099 ^ Bit_1144 ^ Bit_1400 ^ Bit_1401;
				Check_250 <= Bit_21 ^ Bit_80 ^ Bit_119 ^ Bit_175 ^ Bit_240 ^ Bit_246 ^ Bit_470 ^ Bit_510 ^ Bit_546 ^ Bit_608 ^ Bit_633 ^ Bit_679 ^ Bit_896 ^ Bit_920 ^ Bit_1004 ^ Bit_1034 ^ Bit_1061 ^ Bit_1125 ^ Bit_1401 ^ Bit_1402;
				Check_251 <= Bit_40 ^ Bit_50 ^ Bit_133 ^ Bit_156 ^ Bit_220 ^ Bit_286 ^ Bit_335 ^ Bit_354 ^ Bit_433 ^ Bit_715 ^ Bit_731 ^ Bit_785 ^ Bit_911 ^ Bit_959 ^ Bit_1002 ^ Bit_1054 ^ Bit_1103 ^ Bit_1151 ^ Bit_1402 ^ Bit_1403;
				Check_252 <= Bit_23 ^ Bit_95 ^ Bit_135 ^ Bit_155 ^ Bit_237 ^ Bit_268 ^ Bit_321 ^ Bit_473 ^ Bit_570 ^ Bit_603 ^ Bit_807 ^ Bit_835 ^ Bit_868 ^ Bit_930 ^ Bit_965 ^ Bit_1032 ^ Bit_1096 ^ Bit_1146 ^ Bit_1403 ^ Bit_1404;
				Check_253 <= Bit_47 ^ Bit_83 ^ Bit_103 ^ Bit_164 ^ Bit_226 ^ Bit_269 ^ Bit_369 ^ Bit_423 ^ Bit_520 ^ Bit_756 ^ Bit_804 ^ Bit_852 ^ Bit_893 ^ Bit_934 ^ Bit_968 ^ Bit_1055 ^ Bit_1081 ^ Bit_1140 ^ Bit_1404 ^ Bit_1405;
				Check_254 <= Bit_8 ^ Bit_57 ^ Bit_113 ^ Bit_161 ^ Bit_238 ^ Bit_259 ^ Bit_310 ^ Bit_417 ^ Bit_506 ^ Bit_666 ^ Bit_679 ^ Bit_847 ^ Bit_889 ^ Bit_952 ^ Bit_983 ^ Bit_1015 ^ Bit_1082 ^ Bit_1113 ^ Bit_1405 ^ Bit_1406;
				Check_255 <= Bit_3 ^ Bit_78 ^ Bit_143 ^ Bit_177 ^ Bit_195 ^ Bit_262 ^ Bit_359 ^ Bit_414 ^ Bit_573 ^ Bit_582 ^ Bit_658 ^ Bit_762 ^ Bit_893 ^ Bit_937 ^ Bit_962 ^ Bit_1022 ^ Bit_1100 ^ Bit_1145 ^ Bit_1406 ^ Bit_1407;
				Check_256 <= Bit_22 ^ Bit_81 ^ Bit_120 ^ Bit_176 ^ Bit_193 ^ Bit_247 ^ Bit_471 ^ Bit_511 ^ Bit_547 ^ Bit_609 ^ Bit_634 ^ Bit_680 ^ Bit_897 ^ Bit_921 ^ Bit_1005 ^ Bit_1035 ^ Bit_1062 ^ Bit_1126 ^ Bit_1407 ^ Bit_1408;
				Check_257 <= Bit_41 ^ Bit_51 ^ Bit_134 ^ Bit_157 ^ Bit_221 ^ Bit_287 ^ Bit_336 ^ Bit_355 ^ Bit_434 ^ Bit_716 ^ Bit_732 ^ Bit_786 ^ Bit_912 ^ Bit_960 ^ Bit_1003 ^ Bit_1055 ^ Bit_1104 ^ Bit_1152 ^ Bit_1408 ^ Bit_1409;
				Check_258 <= Bit_24 ^ Bit_96 ^ Bit_136 ^ Bit_156 ^ Bit_238 ^ Bit_269 ^ Bit_322 ^ Bit_474 ^ Bit_571 ^ Bit_604 ^ Bit_808 ^ Bit_836 ^ Bit_869 ^ Bit_931 ^ Bit_966 ^ Bit_1033 ^ Bit_1097 ^ Bit_1147 ^ Bit_1409 ^ Bit_1410;
				Check_259 <= Bit_48 ^ Bit_84 ^ Bit_104 ^ Bit_165 ^ Bit_227 ^ Bit_270 ^ Bit_370 ^ Bit_424 ^ Bit_521 ^ Bit_757 ^ Bit_805 ^ Bit_853 ^ Bit_894 ^ Bit_935 ^ Bit_969 ^ Bit_1056 ^ Bit_1082 ^ Bit_1141 ^ Bit_1410 ^ Bit_1411;
				Check_260 <= Bit_9 ^ Bit_58 ^ Bit_114 ^ Bit_162 ^ Bit_239 ^ Bit_260 ^ Bit_311 ^ Bit_418 ^ Bit_507 ^ Bit_667 ^ Bit_680 ^ Bit_848 ^ Bit_890 ^ Bit_953 ^ Bit_984 ^ Bit_1016 ^ Bit_1083 ^ Bit_1114 ^ Bit_1411 ^ Bit_1412;
				Check_261 <= Bit_4 ^ Bit_79 ^ Bit_144 ^ Bit_178 ^ Bit_196 ^ Bit_263 ^ Bit_360 ^ Bit_415 ^ Bit_574 ^ Bit_583 ^ Bit_659 ^ Bit_763 ^ Bit_894 ^ Bit_938 ^ Bit_963 ^ Bit_1023 ^ Bit_1101 ^ Bit_1146 ^ Bit_1412 ^ Bit_1413;
				Check_262 <= Bit_23 ^ Bit_82 ^ Bit_121 ^ Bit_177 ^ Bit_194 ^ Bit_248 ^ Bit_472 ^ Bit_512 ^ Bit_548 ^ Bit_610 ^ Bit_635 ^ Bit_681 ^ Bit_898 ^ Bit_922 ^ Bit_1006 ^ Bit_1036 ^ Bit_1063 ^ Bit_1127 ^ Bit_1413 ^ Bit_1414;
				Check_263 <= Bit_42 ^ Bit_52 ^ Bit_135 ^ Bit_158 ^ Bit_222 ^ Bit_288 ^ Bit_289 ^ Bit_356 ^ Bit_435 ^ Bit_717 ^ Bit_733 ^ Bit_787 ^ Bit_865 ^ Bit_913 ^ Bit_1004 ^ Bit_1056 ^ Bit_1057 ^ Bit_1105 ^ Bit_1414 ^ Bit_1415;
				Check_264 <= Bit_25 ^ Bit_49 ^ Bit_137 ^ Bit_157 ^ Bit_239 ^ Bit_270 ^ Bit_323 ^ Bit_475 ^ Bit_572 ^ Bit_605 ^ Bit_809 ^ Bit_837 ^ Bit_870 ^ Bit_932 ^ Bit_967 ^ Bit_1034 ^ Bit_1098 ^ Bit_1148 ^ Bit_1415 ^ Bit_1416;
				Check_265 <= Bit_1 ^ Bit_85 ^ Bit_105 ^ Bit_166 ^ Bit_228 ^ Bit_271 ^ Bit_371 ^ Bit_425 ^ Bit_522 ^ Bit_758 ^ Bit_806 ^ Bit_854 ^ Bit_895 ^ Bit_936 ^ Bit_970 ^ Bit_1009 ^ Bit_1083 ^ Bit_1142 ^ Bit_1416 ^ Bit_1417;
				Check_266 <= Bit_10 ^ Bit_59 ^ Bit_115 ^ Bit_163 ^ Bit_240 ^ Bit_261 ^ Bit_312 ^ Bit_419 ^ Bit_508 ^ Bit_668 ^ Bit_681 ^ Bit_849 ^ Bit_891 ^ Bit_954 ^ Bit_985 ^ Bit_1017 ^ Bit_1084 ^ Bit_1115 ^ Bit_1417 ^ Bit_1418;
				Check_267 <= Bit_5 ^ Bit_80 ^ Bit_97 ^ Bit_179 ^ Bit_197 ^ Bit_264 ^ Bit_361 ^ Bit_416 ^ Bit_575 ^ Bit_584 ^ Bit_660 ^ Bit_764 ^ Bit_895 ^ Bit_939 ^ Bit_964 ^ Bit_1024 ^ Bit_1102 ^ Bit_1147 ^ Bit_1418 ^ Bit_1419;
				Check_268 <= Bit_24 ^ Bit_83 ^ Bit_122 ^ Bit_178 ^ Bit_195 ^ Bit_249 ^ Bit_473 ^ Bit_513 ^ Bit_549 ^ Bit_611 ^ Bit_636 ^ Bit_682 ^ Bit_899 ^ Bit_923 ^ Bit_1007 ^ Bit_1037 ^ Bit_1064 ^ Bit_1128 ^ Bit_1419 ^ Bit_1420;
				Check_269 <= Bit_43 ^ Bit_53 ^ Bit_136 ^ Bit_159 ^ Bit_223 ^ Bit_241 ^ Bit_290 ^ Bit_357 ^ Bit_436 ^ Bit_718 ^ Bit_734 ^ Bit_788 ^ Bit_866 ^ Bit_914 ^ Bit_1005 ^ Bit_1009 ^ Bit_1058 ^ Bit_1106 ^ Bit_1420 ^ Bit_1421;
				Check_270 <= Bit_26 ^ Bit_50 ^ Bit_138 ^ Bit_158 ^ Bit_240 ^ Bit_271 ^ Bit_324 ^ Bit_476 ^ Bit_573 ^ Bit_606 ^ Bit_810 ^ Bit_838 ^ Bit_871 ^ Bit_933 ^ Bit_968 ^ Bit_1035 ^ Bit_1099 ^ Bit_1149 ^ Bit_1421 ^ Bit_1422;
				Check_271 <= Bit_2 ^ Bit_86 ^ Bit_106 ^ Bit_167 ^ Bit_229 ^ Bit_272 ^ Bit_372 ^ Bit_426 ^ Bit_523 ^ Bit_759 ^ Bit_807 ^ Bit_855 ^ Bit_896 ^ Bit_937 ^ Bit_971 ^ Bit_1010 ^ Bit_1084 ^ Bit_1143 ^ Bit_1422 ^ Bit_1423;
				Check_272 <= Bit_11 ^ Bit_60 ^ Bit_116 ^ Bit_164 ^ Bit_193 ^ Bit_262 ^ Bit_313 ^ Bit_420 ^ Bit_509 ^ Bit_669 ^ Bit_682 ^ Bit_850 ^ Bit_892 ^ Bit_955 ^ Bit_986 ^ Bit_1018 ^ Bit_1085 ^ Bit_1116 ^ Bit_1423 ^ Bit_1424;
				Check_273 <= Bit_6 ^ Bit_81 ^ Bit_98 ^ Bit_180 ^ Bit_198 ^ Bit_265 ^ Bit_362 ^ Bit_417 ^ Bit_576 ^ Bit_585 ^ Bit_661 ^ Bit_765 ^ Bit_896 ^ Bit_940 ^ Bit_965 ^ Bit_1025 ^ Bit_1103 ^ Bit_1148 ^ Bit_1424 ^ Bit_1425;
				Check_274 <= Bit_25 ^ Bit_84 ^ Bit_123 ^ Bit_179 ^ Bit_196 ^ Bit_250 ^ Bit_474 ^ Bit_514 ^ Bit_550 ^ Bit_612 ^ Bit_637 ^ Bit_683 ^ Bit_900 ^ Bit_924 ^ Bit_1008 ^ Bit_1038 ^ Bit_1065 ^ Bit_1129 ^ Bit_1425 ^ Bit_1426;
				Check_275 <= Bit_44 ^ Bit_54 ^ Bit_137 ^ Bit_160 ^ Bit_224 ^ Bit_242 ^ Bit_291 ^ Bit_358 ^ Bit_437 ^ Bit_719 ^ Bit_735 ^ Bit_789 ^ Bit_867 ^ Bit_915 ^ Bit_1006 ^ Bit_1010 ^ Bit_1059 ^ Bit_1107 ^ Bit_1426 ^ Bit_1427;
				Check_276 <= Bit_27 ^ Bit_51 ^ Bit_139 ^ Bit_159 ^ Bit_193 ^ Bit_272 ^ Bit_325 ^ Bit_477 ^ Bit_574 ^ Bit_607 ^ Bit_811 ^ Bit_839 ^ Bit_872 ^ Bit_934 ^ Bit_969 ^ Bit_1036 ^ Bit_1100 ^ Bit_1150 ^ Bit_1427 ^ Bit_1428;
				Check_277 <= Bit_3 ^ Bit_87 ^ Bit_107 ^ Bit_168 ^ Bit_230 ^ Bit_273 ^ Bit_373 ^ Bit_427 ^ Bit_524 ^ Bit_760 ^ Bit_808 ^ Bit_856 ^ Bit_897 ^ Bit_938 ^ Bit_972 ^ Bit_1011 ^ Bit_1085 ^ Bit_1144 ^ Bit_1428 ^ Bit_1429;
				Check_278 <= Bit_12 ^ Bit_61 ^ Bit_117 ^ Bit_165 ^ Bit_194 ^ Bit_263 ^ Bit_314 ^ Bit_421 ^ Bit_510 ^ Bit_670 ^ Bit_683 ^ Bit_851 ^ Bit_893 ^ Bit_956 ^ Bit_987 ^ Bit_1019 ^ Bit_1086 ^ Bit_1117 ^ Bit_1429 ^ Bit_1430;
				Check_279 <= Bit_7 ^ Bit_82 ^ Bit_99 ^ Bit_181 ^ Bit_199 ^ Bit_266 ^ Bit_363 ^ Bit_418 ^ Bit_529 ^ Bit_586 ^ Bit_662 ^ Bit_766 ^ Bit_897 ^ Bit_941 ^ Bit_966 ^ Bit_1026 ^ Bit_1104 ^ Bit_1149 ^ Bit_1430 ^ Bit_1431;
				Check_280 <= Bit_26 ^ Bit_85 ^ Bit_124 ^ Bit_180 ^ Bit_197 ^ Bit_251 ^ Bit_475 ^ Bit_515 ^ Bit_551 ^ Bit_613 ^ Bit_638 ^ Bit_684 ^ Bit_901 ^ Bit_925 ^ Bit_961 ^ Bit_1039 ^ Bit_1066 ^ Bit_1130 ^ Bit_1431 ^ Bit_1432;
				Check_281 <= Bit_45 ^ Bit_55 ^ Bit_138 ^ Bit_161 ^ Bit_225 ^ Bit_243 ^ Bit_292 ^ Bit_359 ^ Bit_438 ^ Bit_720 ^ Bit_736 ^ Bit_790 ^ Bit_868 ^ Bit_916 ^ Bit_1007 ^ Bit_1011 ^ Bit_1060 ^ Bit_1108 ^ Bit_1432 ^ Bit_1433;
				Check_282 <= Bit_28 ^ Bit_52 ^ Bit_140 ^ Bit_160 ^ Bit_194 ^ Bit_273 ^ Bit_326 ^ Bit_478 ^ Bit_575 ^ Bit_608 ^ Bit_812 ^ Bit_840 ^ Bit_873 ^ Bit_935 ^ Bit_970 ^ Bit_1037 ^ Bit_1101 ^ Bit_1151 ^ Bit_1433 ^ Bit_1434;
				Check_283 <= Bit_4 ^ Bit_88 ^ Bit_108 ^ Bit_169 ^ Bit_231 ^ Bit_274 ^ Bit_374 ^ Bit_428 ^ Bit_525 ^ Bit_761 ^ Bit_809 ^ Bit_857 ^ Bit_898 ^ Bit_939 ^ Bit_973 ^ Bit_1012 ^ Bit_1086 ^ Bit_1145 ^ Bit_1434 ^ Bit_1435;
				Check_284 <= Bit_13 ^ Bit_62 ^ Bit_118 ^ Bit_166 ^ Bit_195 ^ Bit_264 ^ Bit_315 ^ Bit_422 ^ Bit_511 ^ Bit_671 ^ Bit_684 ^ Bit_852 ^ Bit_894 ^ Bit_957 ^ Bit_988 ^ Bit_1020 ^ Bit_1087 ^ Bit_1118 ^ Bit_1435 ^ Bit_1436;
				Check_285 <= Bit_8 ^ Bit_83 ^ Bit_100 ^ Bit_182 ^ Bit_200 ^ Bit_267 ^ Bit_364 ^ Bit_419 ^ Bit_530 ^ Bit_587 ^ Bit_663 ^ Bit_767 ^ Bit_898 ^ Bit_942 ^ Bit_967 ^ Bit_1027 ^ Bit_1057 ^ Bit_1150 ^ Bit_1436 ^ Bit_1437;
				Check_286 <= Bit_27 ^ Bit_86 ^ Bit_125 ^ Bit_181 ^ Bit_198 ^ Bit_252 ^ Bit_476 ^ Bit_516 ^ Bit_552 ^ Bit_614 ^ Bit_639 ^ Bit_685 ^ Bit_902 ^ Bit_926 ^ Bit_962 ^ Bit_1040 ^ Bit_1067 ^ Bit_1131 ^ Bit_1437 ^ Bit_1438;
				Check_287 <= Bit_46 ^ Bit_56 ^ Bit_139 ^ Bit_162 ^ Bit_226 ^ Bit_244 ^ Bit_293 ^ Bit_360 ^ Bit_439 ^ Bit_673 ^ Bit_737 ^ Bit_791 ^ Bit_869 ^ Bit_917 ^ Bit_1008 ^ Bit_1012 ^ Bit_1061 ^ Bit_1109 ^ Bit_1438 ^ Bit_1439;
				Check_288 <= Bit_29 ^ Bit_53 ^ Bit_141 ^ Bit_161 ^ Bit_195 ^ Bit_274 ^ Bit_327 ^ Bit_479 ^ Bit_576 ^ Bit_609 ^ Bit_813 ^ Bit_841 ^ Bit_874 ^ Bit_936 ^ Bit_971 ^ Bit_1038 ^ Bit_1102 ^ Bit_1152 ^ Bit_1439 ^ Bit_1440;
				cnt <= cnt + 1;
			end
			else if (cnt == 8'd16) begin
				Check_Sum <= Check_1 | Check_2 | Check_3 | Check_4 | Check_5 | Check_6 | Check_7 | Check_8 | Check_9 | Check_10 | Check_11 | Check_12 | Check_13 | Check_14 | Check_15 | Check_16 | Check_17 | Check_18 | Check_19 | Check_20 | Check_21 | Check_22 | Check_23 | Check_24 | Check_25 | Check_26 | Check_27 | Check_28 | Check_29 | Check_30 | Check_31 | Check_32 | Check_33 | Check_34 | Check_35 | Check_36 | Check_37 | Check_38 | Check_39 | Check_40 | Check_41 | Check_42 | Check_43 | Check_44 | Check_45 | Check_46 | Check_47 | Check_48 | Check_49 | Check_50 | Check_51 | Check_52 | Check_53 | Check_54 | Check_55 | Check_56 | Check_57 | Check_58 | Check_59 | Check_60 | Check_61 | Check_62 | Check_63 | Check_64 | Check_65 | Check_66 | Check_67 | Check_68 | Check_69 | Check_70 | Check_71 | Check_72 | Check_73 | Check_74 | Check_75 | Check_76 | Check_77 | Check_78 | Check_79 | Check_80 | Check_81 | Check_82 | Check_83 | Check_84 | Check_85 | Check_86 | Check_87 | Check_88 | Check_89 | Check_90 | Check_91 | Check_92 | Check_93 | Check_94 | Check_95 | Check_96 | Check_97 | Check_98 | Check_99 | Check_100 | Check_101 | Check_102 | Check_103 | Check_104 | Check_105 | Check_106 | Check_107 | Check_108 | Check_109 | Check_110 | Check_111 | Check_112 | Check_113 | Check_114 | Check_115 | Check_116 | Check_117 | Check_118 | Check_119 | Check_120 | Check_121 | Check_122 | Check_123 | Check_124 | Check_125 | Check_126 | Check_127 | Check_128 | Check_129 | Check_130 | Check_131 | Check_132 | Check_133 | Check_134 | Check_135 | Check_136 | Check_137 | Check_138 | Check_139 | Check_140 | Check_141 | Check_142 | Check_143 | Check_144 | Check_145 | Check_146 | Check_147 | Check_148 | Check_149 | Check_150 | Check_151 | Check_152 | Check_153 | Check_154 | Check_155 | Check_156 | Check_157 | Check_158 | Check_159 | Check_160 | Check_161 | Check_162 | Check_163 | Check_164 | Check_165 | Check_166 | Check_167 | Check_168 | Check_169 | Check_170 | Check_171 | Check_172 | Check_173 | Check_174 | Check_175 | Check_176 | Check_177 | Check_178 | Check_179 | Check_180 | Check_181 | Check_182 | Check_183 | Check_184 | Check_185 | Check_186 | Check_187 | Check_188 | Check_189 | Check_190 | Check_191 | Check_192 | Check_193 | Check_194 | Check_195 | Check_196 | Check_197 | Check_198 | Check_199 | Check_200 | Check_201 | Check_202 | Check_203 | Check_204 | Check_205 | Check_206 | Check_207 | Check_208 | Check_209 | Check_210 | Check_211 | Check_212 | Check_213 | Check_214 | Check_215 | Check_216 | Check_217 | Check_218 | Check_219 | Check_220 | Check_221 | Check_222 | Check_223 | Check_224 | Check_225 | Check_226 | Check_227 | Check_228 | Check_229 | Check_230 | Check_231 | Check_232 | Check_233 | Check_234 | Check_235 | Check_236 | Check_237 | Check_238 | Check_239 | Check_240 | Check_241 | Check_242 | Check_243 | Check_244 | Check_245 | Check_246 | Check_247 | Check_248 | Check_249 | Check_250 | Check_251 | Check_252 | Check_253 | Check_254 | Check_255 | Check_256 | Check_257 | Check_258 | Check_259 | Check_260 | Check_261 | Check_262 | Check_263 | Check_264 | Check_265 | Check_266 | Check_267 | Check_268 | Check_269 | Check_270 | Check_271 | Check_272 | Check_273 | Check_274 | Check_275 | Check_276 | Check_277 | Check_278 | Check_279 | Check_280 | Check_281 | Check_282 | Check_283 | Check_284 | Check_285 | Check_286 | Check_287 | Check_288;
				cnt <= cnt + 1;
			end
			else if (cnt == 8'd17) begin
				if (Check_Sum == 0 || iter == 5'd30) begin
					cnt <= cnt + 1;
					out_valid <= 1;
				end
				else begin
					out_valid <= 0;
					cnt <= 2;
					iter <= iter + 1;
				end
			end
		end
	end
end
assign Bit_1 = V_1[quan_width-1];
assign Bit_2 = V_2[quan_width-1];
assign Bit_3 = V_3[quan_width-1];
assign Bit_4 = V_4[quan_width-1];
assign Bit_5 = V_5[quan_width-1];
assign Bit_6 = V_6[quan_width-1];
assign Bit_7 = V_7[quan_width-1];
assign Bit_8 = V_8[quan_width-1];
assign Bit_9 = V_9[quan_width-1];
assign Bit_10 = V_10[quan_width-1];
assign Bit_11 = V_11[quan_width-1];
assign Bit_12 = V_12[quan_width-1];
assign Bit_13 = V_13[quan_width-1];
assign Bit_14 = V_14[quan_width-1];
assign Bit_15 = V_15[quan_width-1];
assign Bit_16 = V_16[quan_width-1];
assign Bit_17 = V_17[quan_width-1];
assign Bit_18 = V_18[quan_width-1];
assign Bit_19 = V_19[quan_width-1];
assign Bit_20 = V_20[quan_width-1];
assign Bit_21 = V_21[quan_width-1];
assign Bit_22 = V_22[quan_width-1];
assign Bit_23 = V_23[quan_width-1];
assign Bit_24 = V_24[quan_width-1];
assign Bit_25 = V_25[quan_width-1];
assign Bit_26 = V_26[quan_width-1];
assign Bit_27 = V_27[quan_width-1];
assign Bit_28 = V_28[quan_width-1];
assign Bit_29 = V_29[quan_width-1];
assign Bit_30 = V_30[quan_width-1];
assign Bit_31 = V_31[quan_width-1];
assign Bit_32 = V_32[quan_width-1];
assign Bit_33 = V_33[quan_width-1];
assign Bit_34 = V_34[quan_width-1];
assign Bit_35 = V_35[quan_width-1];
assign Bit_36 = V_36[quan_width-1];
assign Bit_37 = V_37[quan_width-1];
assign Bit_38 = V_38[quan_width-1];
assign Bit_39 = V_39[quan_width-1];
assign Bit_40 = V_40[quan_width-1];
assign Bit_41 = V_41[quan_width-1];
assign Bit_42 = V_42[quan_width-1];
assign Bit_43 = V_43[quan_width-1];
assign Bit_44 = V_44[quan_width-1];
assign Bit_45 = V_45[quan_width-1];
assign Bit_46 = V_46[quan_width-1];
assign Bit_47 = V_47[quan_width-1];
assign Bit_48 = V_48[quan_width-1];
assign Bit_49 = V_49[quan_width-1];
assign Bit_50 = V_50[quan_width-1];
assign Bit_51 = V_51[quan_width-1];
assign Bit_52 = V_52[quan_width-1];
assign Bit_53 = V_53[quan_width-1];
assign Bit_54 = V_54[quan_width-1];
assign Bit_55 = V_55[quan_width-1];
assign Bit_56 = V_56[quan_width-1];
assign Bit_57 = V_57[quan_width-1];
assign Bit_58 = V_58[quan_width-1];
assign Bit_59 = V_59[quan_width-1];
assign Bit_60 = V_60[quan_width-1];
assign Bit_61 = V_61[quan_width-1];
assign Bit_62 = V_62[quan_width-1];
assign Bit_63 = V_63[quan_width-1];
assign Bit_64 = V_64[quan_width-1];
assign Bit_65 = V_65[quan_width-1];
assign Bit_66 = V_66[quan_width-1];
assign Bit_67 = V_67[quan_width-1];
assign Bit_68 = V_68[quan_width-1];
assign Bit_69 = V_69[quan_width-1];
assign Bit_70 = V_70[quan_width-1];
assign Bit_71 = V_71[quan_width-1];
assign Bit_72 = V_72[quan_width-1];
assign Bit_73 = V_73[quan_width-1];
assign Bit_74 = V_74[quan_width-1];
assign Bit_75 = V_75[quan_width-1];
assign Bit_76 = V_76[quan_width-1];
assign Bit_77 = V_77[quan_width-1];
assign Bit_78 = V_78[quan_width-1];
assign Bit_79 = V_79[quan_width-1];
assign Bit_80 = V_80[quan_width-1];
assign Bit_81 = V_81[quan_width-1];
assign Bit_82 = V_82[quan_width-1];
assign Bit_83 = V_83[quan_width-1];
assign Bit_84 = V_84[quan_width-1];
assign Bit_85 = V_85[quan_width-1];
assign Bit_86 = V_86[quan_width-1];
assign Bit_87 = V_87[quan_width-1];
assign Bit_88 = V_88[quan_width-1];
assign Bit_89 = V_89[quan_width-1];
assign Bit_90 = V_90[quan_width-1];
assign Bit_91 = V_91[quan_width-1];
assign Bit_92 = V_92[quan_width-1];
assign Bit_93 = V_93[quan_width-1];
assign Bit_94 = V_94[quan_width-1];
assign Bit_95 = V_95[quan_width-1];
assign Bit_96 = V_96[quan_width-1];
assign Bit_97 = V_97[quan_width-1];
assign Bit_98 = V_98[quan_width-1];
assign Bit_99 = V_99[quan_width-1];
assign Bit_100 = V_100[quan_width-1];
assign Bit_101 = V_101[quan_width-1];
assign Bit_102 = V_102[quan_width-1];
assign Bit_103 = V_103[quan_width-1];
assign Bit_104 = V_104[quan_width-1];
assign Bit_105 = V_105[quan_width-1];
assign Bit_106 = V_106[quan_width-1];
assign Bit_107 = V_107[quan_width-1];
assign Bit_108 = V_108[quan_width-1];
assign Bit_109 = V_109[quan_width-1];
assign Bit_110 = V_110[quan_width-1];
assign Bit_111 = V_111[quan_width-1];
assign Bit_112 = V_112[quan_width-1];
assign Bit_113 = V_113[quan_width-1];
assign Bit_114 = V_114[quan_width-1];
assign Bit_115 = V_115[quan_width-1];
assign Bit_116 = V_116[quan_width-1];
assign Bit_117 = V_117[quan_width-1];
assign Bit_118 = V_118[quan_width-1];
assign Bit_119 = V_119[quan_width-1];
assign Bit_120 = V_120[quan_width-1];
assign Bit_121 = V_121[quan_width-1];
assign Bit_122 = V_122[quan_width-1];
assign Bit_123 = V_123[quan_width-1];
assign Bit_124 = V_124[quan_width-1];
assign Bit_125 = V_125[quan_width-1];
assign Bit_126 = V_126[quan_width-1];
assign Bit_127 = V_127[quan_width-1];
assign Bit_128 = V_128[quan_width-1];
assign Bit_129 = V_129[quan_width-1];
assign Bit_130 = V_130[quan_width-1];
assign Bit_131 = V_131[quan_width-1];
assign Bit_132 = V_132[quan_width-1];
assign Bit_133 = V_133[quan_width-1];
assign Bit_134 = V_134[quan_width-1];
assign Bit_135 = V_135[quan_width-1];
assign Bit_136 = V_136[quan_width-1];
assign Bit_137 = V_137[quan_width-1];
assign Bit_138 = V_138[quan_width-1];
assign Bit_139 = V_139[quan_width-1];
assign Bit_140 = V_140[quan_width-1];
assign Bit_141 = V_141[quan_width-1];
assign Bit_142 = V_142[quan_width-1];
assign Bit_143 = V_143[quan_width-1];
assign Bit_144 = V_144[quan_width-1];
assign Bit_145 = V_145[quan_width-1];
assign Bit_146 = V_146[quan_width-1];
assign Bit_147 = V_147[quan_width-1];
assign Bit_148 = V_148[quan_width-1];
assign Bit_149 = V_149[quan_width-1];
assign Bit_150 = V_150[quan_width-1];
assign Bit_151 = V_151[quan_width-1];
assign Bit_152 = V_152[quan_width-1];
assign Bit_153 = V_153[quan_width-1];
assign Bit_154 = V_154[quan_width-1];
assign Bit_155 = V_155[quan_width-1];
assign Bit_156 = V_156[quan_width-1];
assign Bit_157 = V_157[quan_width-1];
assign Bit_158 = V_158[quan_width-1];
assign Bit_159 = V_159[quan_width-1];
assign Bit_160 = V_160[quan_width-1];
assign Bit_161 = V_161[quan_width-1];
assign Bit_162 = V_162[quan_width-1];
assign Bit_163 = V_163[quan_width-1];
assign Bit_164 = V_164[quan_width-1];
assign Bit_165 = V_165[quan_width-1];
assign Bit_166 = V_166[quan_width-1];
assign Bit_167 = V_167[quan_width-1];
assign Bit_168 = V_168[quan_width-1];
assign Bit_169 = V_169[quan_width-1];
assign Bit_170 = V_170[quan_width-1];
assign Bit_171 = V_171[quan_width-1];
assign Bit_172 = V_172[quan_width-1];
assign Bit_173 = V_173[quan_width-1];
assign Bit_174 = V_174[quan_width-1];
assign Bit_175 = V_175[quan_width-1];
assign Bit_176 = V_176[quan_width-1];
assign Bit_177 = V_177[quan_width-1];
assign Bit_178 = V_178[quan_width-1];
assign Bit_179 = V_179[quan_width-1];
assign Bit_180 = V_180[quan_width-1];
assign Bit_181 = V_181[quan_width-1];
assign Bit_182 = V_182[quan_width-1];
assign Bit_183 = V_183[quan_width-1];
assign Bit_184 = V_184[quan_width-1];
assign Bit_185 = V_185[quan_width-1];
assign Bit_186 = V_186[quan_width-1];
assign Bit_187 = V_187[quan_width-1];
assign Bit_188 = V_188[quan_width-1];
assign Bit_189 = V_189[quan_width-1];
assign Bit_190 = V_190[quan_width-1];
assign Bit_191 = V_191[quan_width-1];
assign Bit_192 = V_192[quan_width-1];
assign Bit_193 = V_193[quan_width-1];
assign Bit_194 = V_194[quan_width-1];
assign Bit_195 = V_195[quan_width-1];
assign Bit_196 = V_196[quan_width-1];
assign Bit_197 = V_197[quan_width-1];
assign Bit_198 = V_198[quan_width-1];
assign Bit_199 = V_199[quan_width-1];
assign Bit_200 = V_200[quan_width-1];
assign Bit_201 = V_201[quan_width-1];
assign Bit_202 = V_202[quan_width-1];
assign Bit_203 = V_203[quan_width-1];
assign Bit_204 = V_204[quan_width-1];
assign Bit_205 = V_205[quan_width-1];
assign Bit_206 = V_206[quan_width-1];
assign Bit_207 = V_207[quan_width-1];
assign Bit_208 = V_208[quan_width-1];
assign Bit_209 = V_209[quan_width-1];
assign Bit_210 = V_210[quan_width-1];
assign Bit_211 = V_211[quan_width-1];
assign Bit_212 = V_212[quan_width-1];
assign Bit_213 = V_213[quan_width-1];
assign Bit_214 = V_214[quan_width-1];
assign Bit_215 = V_215[quan_width-1];
assign Bit_216 = V_216[quan_width-1];
assign Bit_217 = V_217[quan_width-1];
assign Bit_218 = V_218[quan_width-1];
assign Bit_219 = V_219[quan_width-1];
assign Bit_220 = V_220[quan_width-1];
assign Bit_221 = V_221[quan_width-1];
assign Bit_222 = V_222[quan_width-1];
assign Bit_223 = V_223[quan_width-1];
assign Bit_224 = V_224[quan_width-1];
assign Bit_225 = V_225[quan_width-1];
assign Bit_226 = V_226[quan_width-1];
assign Bit_227 = V_227[quan_width-1];
assign Bit_228 = V_228[quan_width-1];
assign Bit_229 = V_229[quan_width-1];
assign Bit_230 = V_230[quan_width-1];
assign Bit_231 = V_231[quan_width-1];
assign Bit_232 = V_232[quan_width-1];
assign Bit_233 = V_233[quan_width-1];
assign Bit_234 = V_234[quan_width-1];
assign Bit_235 = V_235[quan_width-1];
assign Bit_236 = V_236[quan_width-1];
assign Bit_237 = V_237[quan_width-1];
assign Bit_238 = V_238[quan_width-1];
assign Bit_239 = V_239[quan_width-1];
assign Bit_240 = V_240[quan_width-1];
assign Bit_241 = V_241[quan_width-1];
assign Bit_242 = V_242[quan_width-1];
assign Bit_243 = V_243[quan_width-1];
assign Bit_244 = V_244[quan_width-1];
assign Bit_245 = V_245[quan_width-1];
assign Bit_246 = V_246[quan_width-1];
assign Bit_247 = V_247[quan_width-1];
assign Bit_248 = V_248[quan_width-1];
assign Bit_249 = V_249[quan_width-1];
assign Bit_250 = V_250[quan_width-1];
assign Bit_251 = V_251[quan_width-1];
assign Bit_252 = V_252[quan_width-1];
assign Bit_253 = V_253[quan_width-1];
assign Bit_254 = V_254[quan_width-1];
assign Bit_255 = V_255[quan_width-1];
assign Bit_256 = V_256[quan_width-1];
assign Bit_257 = V_257[quan_width-1];
assign Bit_258 = V_258[quan_width-1];
assign Bit_259 = V_259[quan_width-1];
assign Bit_260 = V_260[quan_width-1];
assign Bit_261 = V_261[quan_width-1];
assign Bit_262 = V_262[quan_width-1];
assign Bit_263 = V_263[quan_width-1];
assign Bit_264 = V_264[quan_width-1];
assign Bit_265 = V_265[quan_width-1];
assign Bit_266 = V_266[quan_width-1];
assign Bit_267 = V_267[quan_width-1];
assign Bit_268 = V_268[quan_width-1];
assign Bit_269 = V_269[quan_width-1];
assign Bit_270 = V_270[quan_width-1];
assign Bit_271 = V_271[quan_width-1];
assign Bit_272 = V_272[quan_width-1];
assign Bit_273 = V_273[quan_width-1];
assign Bit_274 = V_274[quan_width-1];
assign Bit_275 = V_275[quan_width-1];
assign Bit_276 = V_276[quan_width-1];
assign Bit_277 = V_277[quan_width-1];
assign Bit_278 = V_278[quan_width-1];
assign Bit_279 = V_279[quan_width-1];
assign Bit_280 = V_280[quan_width-1];
assign Bit_281 = V_281[quan_width-1];
assign Bit_282 = V_282[quan_width-1];
assign Bit_283 = V_283[quan_width-1];
assign Bit_284 = V_284[quan_width-1];
assign Bit_285 = V_285[quan_width-1];
assign Bit_286 = V_286[quan_width-1];
assign Bit_287 = V_287[quan_width-1];
assign Bit_288 = V_288[quan_width-1];
assign Bit_289 = V_289[quan_width-1];
assign Bit_290 = V_290[quan_width-1];
assign Bit_291 = V_291[quan_width-1];
assign Bit_292 = V_292[quan_width-1];
assign Bit_293 = V_293[quan_width-1];
assign Bit_294 = V_294[quan_width-1];
assign Bit_295 = V_295[quan_width-1];
assign Bit_296 = V_296[quan_width-1];
assign Bit_297 = V_297[quan_width-1];
assign Bit_298 = V_298[quan_width-1];
assign Bit_299 = V_299[quan_width-1];
assign Bit_300 = V_300[quan_width-1];
assign Bit_301 = V_301[quan_width-1];
assign Bit_302 = V_302[quan_width-1];
assign Bit_303 = V_303[quan_width-1];
assign Bit_304 = V_304[quan_width-1];
assign Bit_305 = V_305[quan_width-1];
assign Bit_306 = V_306[quan_width-1];
assign Bit_307 = V_307[quan_width-1];
assign Bit_308 = V_308[quan_width-1];
assign Bit_309 = V_309[quan_width-1];
assign Bit_310 = V_310[quan_width-1];
assign Bit_311 = V_311[quan_width-1];
assign Bit_312 = V_312[quan_width-1];
assign Bit_313 = V_313[quan_width-1];
assign Bit_314 = V_314[quan_width-1];
assign Bit_315 = V_315[quan_width-1];
assign Bit_316 = V_316[quan_width-1];
assign Bit_317 = V_317[quan_width-1];
assign Bit_318 = V_318[quan_width-1];
assign Bit_319 = V_319[quan_width-1];
assign Bit_320 = V_320[quan_width-1];
assign Bit_321 = V_321[quan_width-1];
assign Bit_322 = V_322[quan_width-1];
assign Bit_323 = V_323[quan_width-1];
assign Bit_324 = V_324[quan_width-1];
assign Bit_325 = V_325[quan_width-1];
assign Bit_326 = V_326[quan_width-1];
assign Bit_327 = V_327[quan_width-1];
assign Bit_328 = V_328[quan_width-1];
assign Bit_329 = V_329[quan_width-1];
assign Bit_330 = V_330[quan_width-1];
assign Bit_331 = V_331[quan_width-1];
assign Bit_332 = V_332[quan_width-1];
assign Bit_333 = V_333[quan_width-1];
assign Bit_334 = V_334[quan_width-1];
assign Bit_335 = V_335[quan_width-1];
assign Bit_336 = V_336[quan_width-1];
assign Bit_337 = V_337[quan_width-1];
assign Bit_338 = V_338[quan_width-1];
assign Bit_339 = V_339[quan_width-1];
assign Bit_340 = V_340[quan_width-1];
assign Bit_341 = V_341[quan_width-1];
assign Bit_342 = V_342[quan_width-1];
assign Bit_343 = V_343[quan_width-1];
assign Bit_344 = V_344[quan_width-1];
assign Bit_345 = V_345[quan_width-1];
assign Bit_346 = V_346[quan_width-1];
assign Bit_347 = V_347[quan_width-1];
assign Bit_348 = V_348[quan_width-1];
assign Bit_349 = V_349[quan_width-1];
assign Bit_350 = V_350[quan_width-1];
assign Bit_351 = V_351[quan_width-1];
assign Bit_352 = V_352[quan_width-1];
assign Bit_353 = V_353[quan_width-1];
assign Bit_354 = V_354[quan_width-1];
assign Bit_355 = V_355[quan_width-1];
assign Bit_356 = V_356[quan_width-1];
assign Bit_357 = V_357[quan_width-1];
assign Bit_358 = V_358[quan_width-1];
assign Bit_359 = V_359[quan_width-1];
assign Bit_360 = V_360[quan_width-1];
assign Bit_361 = V_361[quan_width-1];
assign Bit_362 = V_362[quan_width-1];
assign Bit_363 = V_363[quan_width-1];
assign Bit_364 = V_364[quan_width-1];
assign Bit_365 = V_365[quan_width-1];
assign Bit_366 = V_366[quan_width-1];
assign Bit_367 = V_367[quan_width-1];
assign Bit_368 = V_368[quan_width-1];
assign Bit_369 = V_369[quan_width-1];
assign Bit_370 = V_370[quan_width-1];
assign Bit_371 = V_371[quan_width-1];
assign Bit_372 = V_372[quan_width-1];
assign Bit_373 = V_373[quan_width-1];
assign Bit_374 = V_374[quan_width-1];
assign Bit_375 = V_375[quan_width-1];
assign Bit_376 = V_376[quan_width-1];
assign Bit_377 = V_377[quan_width-1];
assign Bit_378 = V_378[quan_width-1];
assign Bit_379 = V_379[quan_width-1];
assign Bit_380 = V_380[quan_width-1];
assign Bit_381 = V_381[quan_width-1];
assign Bit_382 = V_382[quan_width-1];
assign Bit_383 = V_383[quan_width-1];
assign Bit_384 = V_384[quan_width-1];
assign Bit_385 = V_385[quan_width-1];
assign Bit_386 = V_386[quan_width-1];
assign Bit_387 = V_387[quan_width-1];
assign Bit_388 = V_388[quan_width-1];
assign Bit_389 = V_389[quan_width-1];
assign Bit_390 = V_390[quan_width-1];
assign Bit_391 = V_391[quan_width-1];
assign Bit_392 = V_392[quan_width-1];
assign Bit_393 = V_393[quan_width-1];
assign Bit_394 = V_394[quan_width-1];
assign Bit_395 = V_395[quan_width-1];
assign Bit_396 = V_396[quan_width-1];
assign Bit_397 = V_397[quan_width-1];
assign Bit_398 = V_398[quan_width-1];
assign Bit_399 = V_399[quan_width-1];
assign Bit_400 = V_400[quan_width-1];
assign Bit_401 = V_401[quan_width-1];
assign Bit_402 = V_402[quan_width-1];
assign Bit_403 = V_403[quan_width-1];
assign Bit_404 = V_404[quan_width-1];
assign Bit_405 = V_405[quan_width-1];
assign Bit_406 = V_406[quan_width-1];
assign Bit_407 = V_407[quan_width-1];
assign Bit_408 = V_408[quan_width-1];
assign Bit_409 = V_409[quan_width-1];
assign Bit_410 = V_410[quan_width-1];
assign Bit_411 = V_411[quan_width-1];
assign Bit_412 = V_412[quan_width-1];
assign Bit_413 = V_413[quan_width-1];
assign Bit_414 = V_414[quan_width-1];
assign Bit_415 = V_415[quan_width-1];
assign Bit_416 = V_416[quan_width-1];
assign Bit_417 = V_417[quan_width-1];
assign Bit_418 = V_418[quan_width-1];
assign Bit_419 = V_419[quan_width-1];
assign Bit_420 = V_420[quan_width-1];
assign Bit_421 = V_421[quan_width-1];
assign Bit_422 = V_422[quan_width-1];
assign Bit_423 = V_423[quan_width-1];
assign Bit_424 = V_424[quan_width-1];
assign Bit_425 = V_425[quan_width-1];
assign Bit_426 = V_426[quan_width-1];
assign Bit_427 = V_427[quan_width-1];
assign Bit_428 = V_428[quan_width-1];
assign Bit_429 = V_429[quan_width-1];
assign Bit_430 = V_430[quan_width-1];
assign Bit_431 = V_431[quan_width-1];
assign Bit_432 = V_432[quan_width-1];
assign Bit_433 = V_433[quan_width-1];
assign Bit_434 = V_434[quan_width-1];
assign Bit_435 = V_435[quan_width-1];
assign Bit_436 = V_436[quan_width-1];
assign Bit_437 = V_437[quan_width-1];
assign Bit_438 = V_438[quan_width-1];
assign Bit_439 = V_439[quan_width-1];
assign Bit_440 = V_440[quan_width-1];
assign Bit_441 = V_441[quan_width-1];
assign Bit_442 = V_442[quan_width-1];
assign Bit_443 = V_443[quan_width-1];
assign Bit_444 = V_444[quan_width-1];
assign Bit_445 = V_445[quan_width-1];
assign Bit_446 = V_446[quan_width-1];
assign Bit_447 = V_447[quan_width-1];
assign Bit_448 = V_448[quan_width-1];
assign Bit_449 = V_449[quan_width-1];
assign Bit_450 = V_450[quan_width-1];
assign Bit_451 = V_451[quan_width-1];
assign Bit_452 = V_452[quan_width-1];
assign Bit_453 = V_453[quan_width-1];
assign Bit_454 = V_454[quan_width-1];
assign Bit_455 = V_455[quan_width-1];
assign Bit_456 = V_456[quan_width-1];
assign Bit_457 = V_457[quan_width-1];
assign Bit_458 = V_458[quan_width-1];
assign Bit_459 = V_459[quan_width-1];
assign Bit_460 = V_460[quan_width-1];
assign Bit_461 = V_461[quan_width-1];
assign Bit_462 = V_462[quan_width-1];
assign Bit_463 = V_463[quan_width-1];
assign Bit_464 = V_464[quan_width-1];
assign Bit_465 = V_465[quan_width-1];
assign Bit_466 = V_466[quan_width-1];
assign Bit_467 = V_467[quan_width-1];
assign Bit_468 = V_468[quan_width-1];
assign Bit_469 = V_469[quan_width-1];
assign Bit_470 = V_470[quan_width-1];
assign Bit_471 = V_471[quan_width-1];
assign Bit_472 = V_472[quan_width-1];
assign Bit_473 = V_473[quan_width-1];
assign Bit_474 = V_474[quan_width-1];
assign Bit_475 = V_475[quan_width-1];
assign Bit_476 = V_476[quan_width-1];
assign Bit_477 = V_477[quan_width-1];
assign Bit_478 = V_478[quan_width-1];
assign Bit_479 = V_479[quan_width-1];
assign Bit_480 = V_480[quan_width-1];
assign Bit_481 = V_481[quan_width-1];
assign Bit_482 = V_482[quan_width-1];
assign Bit_483 = V_483[quan_width-1];
assign Bit_484 = V_484[quan_width-1];
assign Bit_485 = V_485[quan_width-1];
assign Bit_486 = V_486[quan_width-1];
assign Bit_487 = V_487[quan_width-1];
assign Bit_488 = V_488[quan_width-1];
assign Bit_489 = V_489[quan_width-1];
assign Bit_490 = V_490[quan_width-1];
assign Bit_491 = V_491[quan_width-1];
assign Bit_492 = V_492[quan_width-1];
assign Bit_493 = V_493[quan_width-1];
assign Bit_494 = V_494[quan_width-1];
assign Bit_495 = V_495[quan_width-1];
assign Bit_496 = V_496[quan_width-1];
assign Bit_497 = V_497[quan_width-1];
assign Bit_498 = V_498[quan_width-1];
assign Bit_499 = V_499[quan_width-1];
assign Bit_500 = V_500[quan_width-1];
assign Bit_501 = V_501[quan_width-1];
assign Bit_502 = V_502[quan_width-1];
assign Bit_503 = V_503[quan_width-1];
assign Bit_504 = V_504[quan_width-1];
assign Bit_505 = V_505[quan_width-1];
assign Bit_506 = V_506[quan_width-1];
assign Bit_507 = V_507[quan_width-1];
assign Bit_508 = V_508[quan_width-1];
assign Bit_509 = V_509[quan_width-1];
assign Bit_510 = V_510[quan_width-1];
assign Bit_511 = V_511[quan_width-1];
assign Bit_512 = V_512[quan_width-1];
assign Bit_513 = V_513[quan_width-1];
assign Bit_514 = V_514[quan_width-1];
assign Bit_515 = V_515[quan_width-1];
assign Bit_516 = V_516[quan_width-1];
assign Bit_517 = V_517[quan_width-1];
assign Bit_518 = V_518[quan_width-1];
assign Bit_519 = V_519[quan_width-1];
assign Bit_520 = V_520[quan_width-1];
assign Bit_521 = V_521[quan_width-1];
assign Bit_522 = V_522[quan_width-1];
assign Bit_523 = V_523[quan_width-1];
assign Bit_524 = V_524[quan_width-1];
assign Bit_525 = V_525[quan_width-1];
assign Bit_526 = V_526[quan_width-1];
assign Bit_527 = V_527[quan_width-1];
assign Bit_528 = V_528[quan_width-1];
assign Bit_529 = V_529[quan_width-1];
assign Bit_530 = V_530[quan_width-1];
assign Bit_531 = V_531[quan_width-1];
assign Bit_532 = V_532[quan_width-1];
assign Bit_533 = V_533[quan_width-1];
assign Bit_534 = V_534[quan_width-1];
assign Bit_535 = V_535[quan_width-1];
assign Bit_536 = V_536[quan_width-1];
assign Bit_537 = V_537[quan_width-1];
assign Bit_538 = V_538[quan_width-1];
assign Bit_539 = V_539[quan_width-1];
assign Bit_540 = V_540[quan_width-1];
assign Bit_541 = V_541[quan_width-1];
assign Bit_542 = V_542[quan_width-1];
assign Bit_543 = V_543[quan_width-1];
assign Bit_544 = V_544[quan_width-1];
assign Bit_545 = V_545[quan_width-1];
assign Bit_546 = V_546[quan_width-1];
assign Bit_547 = V_547[quan_width-1];
assign Bit_548 = V_548[quan_width-1];
assign Bit_549 = V_549[quan_width-1];
assign Bit_550 = V_550[quan_width-1];
assign Bit_551 = V_551[quan_width-1];
assign Bit_552 = V_552[quan_width-1];
assign Bit_553 = V_553[quan_width-1];
assign Bit_554 = V_554[quan_width-1];
assign Bit_555 = V_555[quan_width-1];
assign Bit_556 = V_556[quan_width-1];
assign Bit_557 = V_557[quan_width-1];
assign Bit_558 = V_558[quan_width-1];
assign Bit_559 = V_559[quan_width-1];
assign Bit_560 = V_560[quan_width-1];
assign Bit_561 = V_561[quan_width-1];
assign Bit_562 = V_562[quan_width-1];
assign Bit_563 = V_563[quan_width-1];
assign Bit_564 = V_564[quan_width-1];
assign Bit_565 = V_565[quan_width-1];
assign Bit_566 = V_566[quan_width-1];
assign Bit_567 = V_567[quan_width-1];
assign Bit_568 = V_568[quan_width-1];
assign Bit_569 = V_569[quan_width-1];
assign Bit_570 = V_570[quan_width-1];
assign Bit_571 = V_571[quan_width-1];
assign Bit_572 = V_572[quan_width-1];
assign Bit_573 = V_573[quan_width-1];
assign Bit_574 = V_574[quan_width-1];
assign Bit_575 = V_575[quan_width-1];
assign Bit_576 = V_576[quan_width-1];
assign Bit_577 = V_577[quan_width-1];
assign Bit_578 = V_578[quan_width-1];
assign Bit_579 = V_579[quan_width-1];
assign Bit_580 = V_580[quan_width-1];
assign Bit_581 = V_581[quan_width-1];
assign Bit_582 = V_582[quan_width-1];
assign Bit_583 = V_583[quan_width-1];
assign Bit_584 = V_584[quan_width-1];
assign Bit_585 = V_585[quan_width-1];
assign Bit_586 = V_586[quan_width-1];
assign Bit_587 = V_587[quan_width-1];
assign Bit_588 = V_588[quan_width-1];
assign Bit_589 = V_589[quan_width-1];
assign Bit_590 = V_590[quan_width-1];
assign Bit_591 = V_591[quan_width-1];
assign Bit_592 = V_592[quan_width-1];
assign Bit_593 = V_593[quan_width-1];
assign Bit_594 = V_594[quan_width-1];
assign Bit_595 = V_595[quan_width-1];
assign Bit_596 = V_596[quan_width-1];
assign Bit_597 = V_597[quan_width-1];
assign Bit_598 = V_598[quan_width-1];
assign Bit_599 = V_599[quan_width-1];
assign Bit_600 = V_600[quan_width-1];
assign Bit_601 = V_601[quan_width-1];
assign Bit_602 = V_602[quan_width-1];
assign Bit_603 = V_603[quan_width-1];
assign Bit_604 = V_604[quan_width-1];
assign Bit_605 = V_605[quan_width-1];
assign Bit_606 = V_606[quan_width-1];
assign Bit_607 = V_607[quan_width-1];
assign Bit_608 = V_608[quan_width-1];
assign Bit_609 = V_609[quan_width-1];
assign Bit_610 = V_610[quan_width-1];
assign Bit_611 = V_611[quan_width-1];
assign Bit_612 = V_612[quan_width-1];
assign Bit_613 = V_613[quan_width-1];
assign Bit_614 = V_614[quan_width-1];
assign Bit_615 = V_615[quan_width-1];
assign Bit_616 = V_616[quan_width-1];
assign Bit_617 = V_617[quan_width-1];
assign Bit_618 = V_618[quan_width-1];
assign Bit_619 = V_619[quan_width-1];
assign Bit_620 = V_620[quan_width-1];
assign Bit_621 = V_621[quan_width-1];
assign Bit_622 = V_622[quan_width-1];
assign Bit_623 = V_623[quan_width-1];
assign Bit_624 = V_624[quan_width-1];
assign Bit_625 = V_625[quan_width-1];
assign Bit_626 = V_626[quan_width-1];
assign Bit_627 = V_627[quan_width-1];
assign Bit_628 = V_628[quan_width-1];
assign Bit_629 = V_629[quan_width-1];
assign Bit_630 = V_630[quan_width-1];
assign Bit_631 = V_631[quan_width-1];
assign Bit_632 = V_632[quan_width-1];
assign Bit_633 = V_633[quan_width-1];
assign Bit_634 = V_634[quan_width-1];
assign Bit_635 = V_635[quan_width-1];
assign Bit_636 = V_636[quan_width-1];
assign Bit_637 = V_637[quan_width-1];
assign Bit_638 = V_638[quan_width-1];
assign Bit_639 = V_639[quan_width-1];
assign Bit_640 = V_640[quan_width-1];
assign Bit_641 = V_641[quan_width-1];
assign Bit_642 = V_642[quan_width-1];
assign Bit_643 = V_643[quan_width-1];
assign Bit_644 = V_644[quan_width-1];
assign Bit_645 = V_645[quan_width-1];
assign Bit_646 = V_646[quan_width-1];
assign Bit_647 = V_647[quan_width-1];
assign Bit_648 = V_648[quan_width-1];
assign Bit_649 = V_649[quan_width-1];
assign Bit_650 = V_650[quan_width-1];
assign Bit_651 = V_651[quan_width-1];
assign Bit_652 = V_652[quan_width-1];
assign Bit_653 = V_653[quan_width-1];
assign Bit_654 = V_654[quan_width-1];
assign Bit_655 = V_655[quan_width-1];
assign Bit_656 = V_656[quan_width-1];
assign Bit_657 = V_657[quan_width-1];
assign Bit_658 = V_658[quan_width-1];
assign Bit_659 = V_659[quan_width-1];
assign Bit_660 = V_660[quan_width-1];
assign Bit_661 = V_661[quan_width-1];
assign Bit_662 = V_662[quan_width-1];
assign Bit_663 = V_663[quan_width-1];
assign Bit_664 = V_664[quan_width-1];
assign Bit_665 = V_665[quan_width-1];
assign Bit_666 = V_666[quan_width-1];
assign Bit_667 = V_667[quan_width-1];
assign Bit_668 = V_668[quan_width-1];
assign Bit_669 = V_669[quan_width-1];
assign Bit_670 = V_670[quan_width-1];
assign Bit_671 = V_671[quan_width-1];
assign Bit_672 = V_672[quan_width-1];
assign Bit_673 = V_673[quan_width-1];
assign Bit_674 = V_674[quan_width-1];
assign Bit_675 = V_675[quan_width-1];
assign Bit_676 = V_676[quan_width-1];
assign Bit_677 = V_677[quan_width-1];
assign Bit_678 = V_678[quan_width-1];
assign Bit_679 = V_679[quan_width-1];
assign Bit_680 = V_680[quan_width-1];
assign Bit_681 = V_681[quan_width-1];
assign Bit_682 = V_682[quan_width-1];
assign Bit_683 = V_683[quan_width-1];
assign Bit_684 = V_684[quan_width-1];
assign Bit_685 = V_685[quan_width-1];
assign Bit_686 = V_686[quan_width-1];
assign Bit_687 = V_687[quan_width-1];
assign Bit_688 = V_688[quan_width-1];
assign Bit_689 = V_689[quan_width-1];
assign Bit_690 = V_690[quan_width-1];
assign Bit_691 = V_691[quan_width-1];
assign Bit_692 = V_692[quan_width-1];
assign Bit_693 = V_693[quan_width-1];
assign Bit_694 = V_694[quan_width-1];
assign Bit_695 = V_695[quan_width-1];
assign Bit_696 = V_696[quan_width-1];
assign Bit_697 = V_697[quan_width-1];
assign Bit_698 = V_698[quan_width-1];
assign Bit_699 = V_699[quan_width-1];
assign Bit_700 = V_700[quan_width-1];
assign Bit_701 = V_701[quan_width-1];
assign Bit_702 = V_702[quan_width-1];
assign Bit_703 = V_703[quan_width-1];
assign Bit_704 = V_704[quan_width-1];
assign Bit_705 = V_705[quan_width-1];
assign Bit_706 = V_706[quan_width-1];
assign Bit_707 = V_707[quan_width-1];
assign Bit_708 = V_708[quan_width-1];
assign Bit_709 = V_709[quan_width-1];
assign Bit_710 = V_710[quan_width-1];
assign Bit_711 = V_711[quan_width-1];
assign Bit_712 = V_712[quan_width-1];
assign Bit_713 = V_713[quan_width-1];
assign Bit_714 = V_714[quan_width-1];
assign Bit_715 = V_715[quan_width-1];
assign Bit_716 = V_716[quan_width-1];
assign Bit_717 = V_717[quan_width-1];
assign Bit_718 = V_718[quan_width-1];
assign Bit_719 = V_719[quan_width-1];
assign Bit_720 = V_720[quan_width-1];
assign Bit_721 = V_721[quan_width-1];
assign Bit_722 = V_722[quan_width-1];
assign Bit_723 = V_723[quan_width-1];
assign Bit_724 = V_724[quan_width-1];
assign Bit_725 = V_725[quan_width-1];
assign Bit_726 = V_726[quan_width-1];
assign Bit_727 = V_727[quan_width-1];
assign Bit_728 = V_728[quan_width-1];
assign Bit_729 = V_729[quan_width-1];
assign Bit_730 = V_730[quan_width-1];
assign Bit_731 = V_731[quan_width-1];
assign Bit_732 = V_732[quan_width-1];
assign Bit_733 = V_733[quan_width-1];
assign Bit_734 = V_734[quan_width-1];
assign Bit_735 = V_735[quan_width-1];
assign Bit_736 = V_736[quan_width-1];
assign Bit_737 = V_737[quan_width-1];
assign Bit_738 = V_738[quan_width-1];
assign Bit_739 = V_739[quan_width-1];
assign Bit_740 = V_740[quan_width-1];
assign Bit_741 = V_741[quan_width-1];
assign Bit_742 = V_742[quan_width-1];
assign Bit_743 = V_743[quan_width-1];
assign Bit_744 = V_744[quan_width-1];
assign Bit_745 = V_745[quan_width-1];
assign Bit_746 = V_746[quan_width-1];
assign Bit_747 = V_747[quan_width-1];
assign Bit_748 = V_748[quan_width-1];
assign Bit_749 = V_749[quan_width-1];
assign Bit_750 = V_750[quan_width-1];
assign Bit_751 = V_751[quan_width-1];
assign Bit_752 = V_752[quan_width-1];
assign Bit_753 = V_753[quan_width-1];
assign Bit_754 = V_754[quan_width-1];
assign Bit_755 = V_755[quan_width-1];
assign Bit_756 = V_756[quan_width-1];
assign Bit_757 = V_757[quan_width-1];
assign Bit_758 = V_758[quan_width-1];
assign Bit_759 = V_759[quan_width-1];
assign Bit_760 = V_760[quan_width-1];
assign Bit_761 = V_761[quan_width-1];
assign Bit_762 = V_762[quan_width-1];
assign Bit_763 = V_763[quan_width-1];
assign Bit_764 = V_764[quan_width-1];
assign Bit_765 = V_765[quan_width-1];
assign Bit_766 = V_766[quan_width-1];
assign Bit_767 = V_767[quan_width-1];
assign Bit_768 = V_768[quan_width-1];
assign Bit_769 = V_769[quan_width-1];
assign Bit_770 = V_770[quan_width-1];
assign Bit_771 = V_771[quan_width-1];
assign Bit_772 = V_772[quan_width-1];
assign Bit_773 = V_773[quan_width-1];
assign Bit_774 = V_774[quan_width-1];
assign Bit_775 = V_775[quan_width-1];
assign Bit_776 = V_776[quan_width-1];
assign Bit_777 = V_777[quan_width-1];
assign Bit_778 = V_778[quan_width-1];
assign Bit_779 = V_779[quan_width-1];
assign Bit_780 = V_780[quan_width-1];
assign Bit_781 = V_781[quan_width-1];
assign Bit_782 = V_782[quan_width-1];
assign Bit_783 = V_783[quan_width-1];
assign Bit_784 = V_784[quan_width-1];
assign Bit_785 = V_785[quan_width-1];
assign Bit_786 = V_786[quan_width-1];
assign Bit_787 = V_787[quan_width-1];
assign Bit_788 = V_788[quan_width-1];
assign Bit_789 = V_789[quan_width-1];
assign Bit_790 = V_790[quan_width-1];
assign Bit_791 = V_791[quan_width-1];
assign Bit_792 = V_792[quan_width-1];
assign Bit_793 = V_793[quan_width-1];
assign Bit_794 = V_794[quan_width-1];
assign Bit_795 = V_795[quan_width-1];
assign Bit_796 = V_796[quan_width-1];
assign Bit_797 = V_797[quan_width-1];
assign Bit_798 = V_798[quan_width-1];
assign Bit_799 = V_799[quan_width-1];
assign Bit_800 = V_800[quan_width-1];
assign Bit_801 = V_801[quan_width-1];
assign Bit_802 = V_802[quan_width-1];
assign Bit_803 = V_803[quan_width-1];
assign Bit_804 = V_804[quan_width-1];
assign Bit_805 = V_805[quan_width-1];
assign Bit_806 = V_806[quan_width-1];
assign Bit_807 = V_807[quan_width-1];
assign Bit_808 = V_808[quan_width-1];
assign Bit_809 = V_809[quan_width-1];
assign Bit_810 = V_810[quan_width-1];
assign Bit_811 = V_811[quan_width-1];
assign Bit_812 = V_812[quan_width-1];
assign Bit_813 = V_813[quan_width-1];
assign Bit_814 = V_814[quan_width-1];
assign Bit_815 = V_815[quan_width-1];
assign Bit_816 = V_816[quan_width-1];
assign Bit_817 = V_817[quan_width-1];
assign Bit_818 = V_818[quan_width-1];
assign Bit_819 = V_819[quan_width-1];
assign Bit_820 = V_820[quan_width-1];
assign Bit_821 = V_821[quan_width-1];
assign Bit_822 = V_822[quan_width-1];
assign Bit_823 = V_823[quan_width-1];
assign Bit_824 = V_824[quan_width-1];
assign Bit_825 = V_825[quan_width-1];
assign Bit_826 = V_826[quan_width-1];
assign Bit_827 = V_827[quan_width-1];
assign Bit_828 = V_828[quan_width-1];
assign Bit_829 = V_829[quan_width-1];
assign Bit_830 = V_830[quan_width-1];
assign Bit_831 = V_831[quan_width-1];
assign Bit_832 = V_832[quan_width-1];
assign Bit_833 = V_833[quan_width-1];
assign Bit_834 = V_834[quan_width-1];
assign Bit_835 = V_835[quan_width-1];
assign Bit_836 = V_836[quan_width-1];
assign Bit_837 = V_837[quan_width-1];
assign Bit_838 = V_838[quan_width-1];
assign Bit_839 = V_839[quan_width-1];
assign Bit_840 = V_840[quan_width-1];
assign Bit_841 = V_841[quan_width-1];
assign Bit_842 = V_842[quan_width-1];
assign Bit_843 = V_843[quan_width-1];
assign Bit_844 = V_844[quan_width-1];
assign Bit_845 = V_845[quan_width-1];
assign Bit_846 = V_846[quan_width-1];
assign Bit_847 = V_847[quan_width-1];
assign Bit_848 = V_848[quan_width-1];
assign Bit_849 = V_849[quan_width-1];
assign Bit_850 = V_850[quan_width-1];
assign Bit_851 = V_851[quan_width-1];
assign Bit_852 = V_852[quan_width-1];
assign Bit_853 = V_853[quan_width-1];
assign Bit_854 = V_854[quan_width-1];
assign Bit_855 = V_855[quan_width-1];
assign Bit_856 = V_856[quan_width-1];
assign Bit_857 = V_857[quan_width-1];
assign Bit_858 = V_858[quan_width-1];
assign Bit_859 = V_859[quan_width-1];
assign Bit_860 = V_860[quan_width-1];
assign Bit_861 = V_861[quan_width-1];
assign Bit_862 = V_862[quan_width-1];
assign Bit_863 = V_863[quan_width-1];
assign Bit_864 = V_864[quan_width-1];
assign Bit_865 = V_865[quan_width-1];
assign Bit_866 = V_866[quan_width-1];
assign Bit_867 = V_867[quan_width-1];
assign Bit_868 = V_868[quan_width-1];
assign Bit_869 = V_869[quan_width-1];
assign Bit_870 = V_870[quan_width-1];
assign Bit_871 = V_871[quan_width-1];
assign Bit_872 = V_872[quan_width-1];
assign Bit_873 = V_873[quan_width-1];
assign Bit_874 = V_874[quan_width-1];
assign Bit_875 = V_875[quan_width-1];
assign Bit_876 = V_876[quan_width-1];
assign Bit_877 = V_877[quan_width-1];
assign Bit_878 = V_878[quan_width-1];
assign Bit_879 = V_879[quan_width-1];
assign Bit_880 = V_880[quan_width-1];
assign Bit_881 = V_881[quan_width-1];
assign Bit_882 = V_882[quan_width-1];
assign Bit_883 = V_883[quan_width-1];
assign Bit_884 = V_884[quan_width-1];
assign Bit_885 = V_885[quan_width-1];
assign Bit_886 = V_886[quan_width-1];
assign Bit_887 = V_887[quan_width-1];
assign Bit_888 = V_888[quan_width-1];
assign Bit_889 = V_889[quan_width-1];
assign Bit_890 = V_890[quan_width-1];
assign Bit_891 = V_891[quan_width-1];
assign Bit_892 = V_892[quan_width-1];
assign Bit_893 = V_893[quan_width-1];
assign Bit_894 = V_894[quan_width-1];
assign Bit_895 = V_895[quan_width-1];
assign Bit_896 = V_896[quan_width-1];
assign Bit_897 = V_897[quan_width-1];
assign Bit_898 = V_898[quan_width-1];
assign Bit_899 = V_899[quan_width-1];
assign Bit_900 = V_900[quan_width-1];
assign Bit_901 = V_901[quan_width-1];
assign Bit_902 = V_902[quan_width-1];
assign Bit_903 = V_903[quan_width-1];
assign Bit_904 = V_904[quan_width-1];
assign Bit_905 = V_905[quan_width-1];
assign Bit_906 = V_906[quan_width-1];
assign Bit_907 = V_907[quan_width-1];
assign Bit_908 = V_908[quan_width-1];
assign Bit_909 = V_909[quan_width-1];
assign Bit_910 = V_910[quan_width-1];
assign Bit_911 = V_911[quan_width-1];
assign Bit_912 = V_912[quan_width-1];
assign Bit_913 = V_913[quan_width-1];
assign Bit_914 = V_914[quan_width-1];
assign Bit_915 = V_915[quan_width-1];
assign Bit_916 = V_916[quan_width-1];
assign Bit_917 = V_917[quan_width-1];
assign Bit_918 = V_918[quan_width-1];
assign Bit_919 = V_919[quan_width-1];
assign Bit_920 = V_920[quan_width-1];
assign Bit_921 = V_921[quan_width-1];
assign Bit_922 = V_922[quan_width-1];
assign Bit_923 = V_923[quan_width-1];
assign Bit_924 = V_924[quan_width-1];
assign Bit_925 = V_925[quan_width-1];
assign Bit_926 = V_926[quan_width-1];
assign Bit_927 = V_927[quan_width-1];
assign Bit_928 = V_928[quan_width-1];
assign Bit_929 = V_929[quan_width-1];
assign Bit_930 = V_930[quan_width-1];
assign Bit_931 = V_931[quan_width-1];
assign Bit_932 = V_932[quan_width-1];
assign Bit_933 = V_933[quan_width-1];
assign Bit_934 = V_934[quan_width-1];
assign Bit_935 = V_935[quan_width-1];
assign Bit_936 = V_936[quan_width-1];
assign Bit_937 = V_937[quan_width-1];
assign Bit_938 = V_938[quan_width-1];
assign Bit_939 = V_939[quan_width-1];
assign Bit_940 = V_940[quan_width-1];
assign Bit_941 = V_941[quan_width-1];
assign Bit_942 = V_942[quan_width-1];
assign Bit_943 = V_943[quan_width-1];
assign Bit_944 = V_944[quan_width-1];
assign Bit_945 = V_945[quan_width-1];
assign Bit_946 = V_946[quan_width-1];
assign Bit_947 = V_947[quan_width-1];
assign Bit_948 = V_948[quan_width-1];
assign Bit_949 = V_949[quan_width-1];
assign Bit_950 = V_950[quan_width-1];
assign Bit_951 = V_951[quan_width-1];
assign Bit_952 = V_952[quan_width-1];
assign Bit_953 = V_953[quan_width-1];
assign Bit_954 = V_954[quan_width-1];
assign Bit_955 = V_955[quan_width-1];
assign Bit_956 = V_956[quan_width-1];
assign Bit_957 = V_957[quan_width-1];
assign Bit_958 = V_958[quan_width-1];
assign Bit_959 = V_959[quan_width-1];
assign Bit_960 = V_960[quan_width-1];
assign Bit_961 = V_961[quan_width-1];
assign Bit_962 = V_962[quan_width-1];
assign Bit_963 = V_963[quan_width-1];
assign Bit_964 = V_964[quan_width-1];
assign Bit_965 = V_965[quan_width-1];
assign Bit_966 = V_966[quan_width-1];
assign Bit_967 = V_967[quan_width-1];
assign Bit_968 = V_968[quan_width-1];
assign Bit_969 = V_969[quan_width-1];
assign Bit_970 = V_970[quan_width-1];
assign Bit_971 = V_971[quan_width-1];
assign Bit_972 = V_972[quan_width-1];
assign Bit_973 = V_973[quan_width-1];
assign Bit_974 = V_974[quan_width-1];
assign Bit_975 = V_975[quan_width-1];
assign Bit_976 = V_976[quan_width-1];
assign Bit_977 = V_977[quan_width-1];
assign Bit_978 = V_978[quan_width-1];
assign Bit_979 = V_979[quan_width-1];
assign Bit_980 = V_980[quan_width-1];
assign Bit_981 = V_981[quan_width-1];
assign Bit_982 = V_982[quan_width-1];
assign Bit_983 = V_983[quan_width-1];
assign Bit_984 = V_984[quan_width-1];
assign Bit_985 = V_985[quan_width-1];
assign Bit_986 = V_986[quan_width-1];
assign Bit_987 = V_987[quan_width-1];
assign Bit_988 = V_988[quan_width-1];
assign Bit_989 = V_989[quan_width-1];
assign Bit_990 = V_990[quan_width-1];
assign Bit_991 = V_991[quan_width-1];
assign Bit_992 = V_992[quan_width-1];
assign Bit_993 = V_993[quan_width-1];
assign Bit_994 = V_994[quan_width-1];
assign Bit_995 = V_995[quan_width-1];
assign Bit_996 = V_996[quan_width-1];
assign Bit_997 = V_997[quan_width-1];
assign Bit_998 = V_998[quan_width-1];
assign Bit_999 = V_999[quan_width-1];
assign Bit_1000 = V_1000[quan_width-1];
assign Bit_1001 = V_1001[quan_width-1];
assign Bit_1002 = V_1002[quan_width-1];
assign Bit_1003 = V_1003[quan_width-1];
assign Bit_1004 = V_1004[quan_width-1];
assign Bit_1005 = V_1005[quan_width-1];
assign Bit_1006 = V_1006[quan_width-1];
assign Bit_1007 = V_1007[quan_width-1];
assign Bit_1008 = V_1008[quan_width-1];
assign Bit_1009 = V_1009[quan_width-1];
assign Bit_1010 = V_1010[quan_width-1];
assign Bit_1011 = V_1011[quan_width-1];
assign Bit_1012 = V_1012[quan_width-1];
assign Bit_1013 = V_1013[quan_width-1];
assign Bit_1014 = V_1014[quan_width-1];
assign Bit_1015 = V_1015[quan_width-1];
assign Bit_1016 = V_1016[quan_width-1];
assign Bit_1017 = V_1017[quan_width-1];
assign Bit_1018 = V_1018[quan_width-1];
assign Bit_1019 = V_1019[quan_width-1];
assign Bit_1020 = V_1020[quan_width-1];
assign Bit_1021 = V_1021[quan_width-1];
assign Bit_1022 = V_1022[quan_width-1];
assign Bit_1023 = V_1023[quan_width-1];
assign Bit_1024 = V_1024[quan_width-1];
assign Bit_1025 = V_1025[quan_width-1];
assign Bit_1026 = V_1026[quan_width-1];
assign Bit_1027 = V_1027[quan_width-1];
assign Bit_1028 = V_1028[quan_width-1];
assign Bit_1029 = V_1029[quan_width-1];
assign Bit_1030 = V_1030[quan_width-1];
assign Bit_1031 = V_1031[quan_width-1];
assign Bit_1032 = V_1032[quan_width-1];
assign Bit_1033 = V_1033[quan_width-1];
assign Bit_1034 = V_1034[quan_width-1];
assign Bit_1035 = V_1035[quan_width-1];
assign Bit_1036 = V_1036[quan_width-1];
assign Bit_1037 = V_1037[quan_width-1];
assign Bit_1038 = V_1038[quan_width-1];
assign Bit_1039 = V_1039[quan_width-1];
assign Bit_1040 = V_1040[quan_width-1];
assign Bit_1041 = V_1041[quan_width-1];
assign Bit_1042 = V_1042[quan_width-1];
assign Bit_1043 = V_1043[quan_width-1];
assign Bit_1044 = V_1044[quan_width-1];
assign Bit_1045 = V_1045[quan_width-1];
assign Bit_1046 = V_1046[quan_width-1];
assign Bit_1047 = V_1047[quan_width-1];
assign Bit_1048 = V_1048[quan_width-1];
assign Bit_1049 = V_1049[quan_width-1];
assign Bit_1050 = V_1050[quan_width-1];
assign Bit_1051 = V_1051[quan_width-1];
assign Bit_1052 = V_1052[quan_width-1];
assign Bit_1053 = V_1053[quan_width-1];
assign Bit_1054 = V_1054[quan_width-1];
assign Bit_1055 = V_1055[quan_width-1];
assign Bit_1056 = V_1056[quan_width-1];
assign Bit_1057 = V_1057[quan_width-1];
assign Bit_1058 = V_1058[quan_width-1];
assign Bit_1059 = V_1059[quan_width-1];
assign Bit_1060 = V_1060[quan_width-1];
assign Bit_1061 = V_1061[quan_width-1];
assign Bit_1062 = V_1062[quan_width-1];
assign Bit_1063 = V_1063[quan_width-1];
assign Bit_1064 = V_1064[quan_width-1];
assign Bit_1065 = V_1065[quan_width-1];
assign Bit_1066 = V_1066[quan_width-1];
assign Bit_1067 = V_1067[quan_width-1];
assign Bit_1068 = V_1068[quan_width-1];
assign Bit_1069 = V_1069[quan_width-1];
assign Bit_1070 = V_1070[quan_width-1];
assign Bit_1071 = V_1071[quan_width-1];
assign Bit_1072 = V_1072[quan_width-1];
assign Bit_1073 = V_1073[quan_width-1];
assign Bit_1074 = V_1074[quan_width-1];
assign Bit_1075 = V_1075[quan_width-1];
assign Bit_1076 = V_1076[quan_width-1];
assign Bit_1077 = V_1077[quan_width-1];
assign Bit_1078 = V_1078[quan_width-1];
assign Bit_1079 = V_1079[quan_width-1];
assign Bit_1080 = V_1080[quan_width-1];
assign Bit_1081 = V_1081[quan_width-1];
assign Bit_1082 = V_1082[quan_width-1];
assign Bit_1083 = V_1083[quan_width-1];
assign Bit_1084 = V_1084[quan_width-1];
assign Bit_1085 = V_1085[quan_width-1];
assign Bit_1086 = V_1086[quan_width-1];
assign Bit_1087 = V_1087[quan_width-1];
assign Bit_1088 = V_1088[quan_width-1];
assign Bit_1089 = V_1089[quan_width-1];
assign Bit_1090 = V_1090[quan_width-1];
assign Bit_1091 = V_1091[quan_width-1];
assign Bit_1092 = V_1092[quan_width-1];
assign Bit_1093 = V_1093[quan_width-1];
assign Bit_1094 = V_1094[quan_width-1];
assign Bit_1095 = V_1095[quan_width-1];
assign Bit_1096 = V_1096[quan_width-1];
assign Bit_1097 = V_1097[quan_width-1];
assign Bit_1098 = V_1098[quan_width-1];
assign Bit_1099 = V_1099[quan_width-1];
assign Bit_1100 = V_1100[quan_width-1];
assign Bit_1101 = V_1101[quan_width-1];
assign Bit_1102 = V_1102[quan_width-1];
assign Bit_1103 = V_1103[quan_width-1];
assign Bit_1104 = V_1104[quan_width-1];
assign Bit_1105 = V_1105[quan_width-1];
assign Bit_1106 = V_1106[quan_width-1];
assign Bit_1107 = V_1107[quan_width-1];
assign Bit_1108 = V_1108[quan_width-1];
assign Bit_1109 = V_1109[quan_width-1];
assign Bit_1110 = V_1110[quan_width-1];
assign Bit_1111 = V_1111[quan_width-1];
assign Bit_1112 = V_1112[quan_width-1];
assign Bit_1113 = V_1113[quan_width-1];
assign Bit_1114 = V_1114[quan_width-1];
assign Bit_1115 = V_1115[quan_width-1];
assign Bit_1116 = V_1116[quan_width-1];
assign Bit_1117 = V_1117[quan_width-1];
assign Bit_1118 = V_1118[quan_width-1];
assign Bit_1119 = V_1119[quan_width-1];
assign Bit_1120 = V_1120[quan_width-1];
assign Bit_1121 = V_1121[quan_width-1];
assign Bit_1122 = V_1122[quan_width-1];
assign Bit_1123 = V_1123[quan_width-1];
assign Bit_1124 = V_1124[quan_width-1];
assign Bit_1125 = V_1125[quan_width-1];
assign Bit_1126 = V_1126[quan_width-1];
assign Bit_1127 = V_1127[quan_width-1];
assign Bit_1128 = V_1128[quan_width-1];
assign Bit_1129 = V_1129[quan_width-1];
assign Bit_1130 = V_1130[quan_width-1];
assign Bit_1131 = V_1131[quan_width-1];
assign Bit_1132 = V_1132[quan_width-1];
assign Bit_1133 = V_1133[quan_width-1];
assign Bit_1134 = V_1134[quan_width-1];
assign Bit_1135 = V_1135[quan_width-1];
assign Bit_1136 = V_1136[quan_width-1];
assign Bit_1137 = V_1137[quan_width-1];
assign Bit_1138 = V_1138[quan_width-1];
assign Bit_1139 = V_1139[quan_width-1];
assign Bit_1140 = V_1140[quan_width-1];
assign Bit_1141 = V_1141[quan_width-1];
assign Bit_1142 = V_1142[quan_width-1];
assign Bit_1143 = V_1143[quan_width-1];
assign Bit_1144 = V_1144[quan_width-1];
assign Bit_1145 = V_1145[quan_width-1];
assign Bit_1146 = V_1146[quan_width-1];
assign Bit_1147 = V_1147[quan_width-1];
assign Bit_1148 = V_1148[quan_width-1];
assign Bit_1149 = V_1149[quan_width-1];
assign Bit_1150 = V_1150[quan_width-1];
assign Bit_1151 = V_1151[quan_width-1];
assign Bit_1152 = V_1152[quan_width-1];
assign Bit_1153 = V_1153[quan_width-1];
assign Bit_1154 = V_1154[quan_width-1];
assign Bit_1155 = V_1155[quan_width-1];
assign Bit_1156 = V_1156[quan_width-1];
assign Bit_1157 = V_1157[quan_width-1];
assign Bit_1158 = V_1158[quan_width-1];
assign Bit_1159 = V_1159[quan_width-1];
assign Bit_1160 = V_1160[quan_width-1];
assign Bit_1161 = V_1161[quan_width-1];
assign Bit_1162 = V_1162[quan_width-1];
assign Bit_1163 = V_1163[quan_width-1];
assign Bit_1164 = V_1164[quan_width-1];
assign Bit_1165 = V_1165[quan_width-1];
assign Bit_1166 = V_1166[quan_width-1];
assign Bit_1167 = V_1167[quan_width-1];
assign Bit_1168 = V_1168[quan_width-1];
assign Bit_1169 = V_1169[quan_width-1];
assign Bit_1170 = V_1170[quan_width-1];
assign Bit_1171 = V_1171[quan_width-1];
assign Bit_1172 = V_1172[quan_width-1];
assign Bit_1173 = V_1173[quan_width-1];
assign Bit_1174 = V_1174[quan_width-1];
assign Bit_1175 = V_1175[quan_width-1];
assign Bit_1176 = V_1176[quan_width-1];
assign Bit_1177 = V_1177[quan_width-1];
assign Bit_1178 = V_1178[quan_width-1];
assign Bit_1179 = V_1179[quan_width-1];
assign Bit_1180 = V_1180[quan_width-1];
assign Bit_1181 = V_1181[quan_width-1];
assign Bit_1182 = V_1182[quan_width-1];
assign Bit_1183 = V_1183[quan_width-1];
assign Bit_1184 = V_1184[quan_width-1];
assign Bit_1185 = V_1185[quan_width-1];
assign Bit_1186 = V_1186[quan_width-1];
assign Bit_1187 = V_1187[quan_width-1];
assign Bit_1188 = V_1188[quan_width-1];
assign Bit_1189 = V_1189[quan_width-1];
assign Bit_1190 = V_1190[quan_width-1];
assign Bit_1191 = V_1191[quan_width-1];
assign Bit_1192 = V_1192[quan_width-1];
assign Bit_1193 = V_1193[quan_width-1];
assign Bit_1194 = V_1194[quan_width-1];
assign Bit_1195 = V_1195[quan_width-1];
assign Bit_1196 = V_1196[quan_width-1];
assign Bit_1197 = V_1197[quan_width-1];
assign Bit_1198 = V_1198[quan_width-1];
assign Bit_1199 = V_1199[quan_width-1];
assign Bit_1200 = V_1200[quan_width-1];
assign Bit_1201 = V_1201[quan_width-1];
assign Bit_1202 = V_1202[quan_width-1];
assign Bit_1203 = V_1203[quan_width-1];
assign Bit_1204 = V_1204[quan_width-1];
assign Bit_1205 = V_1205[quan_width-1];
assign Bit_1206 = V_1206[quan_width-1];
assign Bit_1207 = V_1207[quan_width-1];
assign Bit_1208 = V_1208[quan_width-1];
assign Bit_1209 = V_1209[quan_width-1];
assign Bit_1210 = V_1210[quan_width-1];
assign Bit_1211 = V_1211[quan_width-1];
assign Bit_1212 = V_1212[quan_width-1];
assign Bit_1213 = V_1213[quan_width-1];
assign Bit_1214 = V_1214[quan_width-1];
assign Bit_1215 = V_1215[quan_width-1];
assign Bit_1216 = V_1216[quan_width-1];
assign Bit_1217 = V_1217[quan_width-1];
assign Bit_1218 = V_1218[quan_width-1];
assign Bit_1219 = V_1219[quan_width-1];
assign Bit_1220 = V_1220[quan_width-1];
assign Bit_1221 = V_1221[quan_width-1];
assign Bit_1222 = V_1222[quan_width-1];
assign Bit_1223 = V_1223[quan_width-1];
assign Bit_1224 = V_1224[quan_width-1];
assign Bit_1225 = V_1225[quan_width-1];
assign Bit_1226 = V_1226[quan_width-1];
assign Bit_1227 = V_1227[quan_width-1];
assign Bit_1228 = V_1228[quan_width-1];
assign Bit_1229 = V_1229[quan_width-1];
assign Bit_1230 = V_1230[quan_width-1];
assign Bit_1231 = V_1231[quan_width-1];
assign Bit_1232 = V_1232[quan_width-1];
assign Bit_1233 = V_1233[quan_width-1];
assign Bit_1234 = V_1234[quan_width-1];
assign Bit_1235 = V_1235[quan_width-1];
assign Bit_1236 = V_1236[quan_width-1];
assign Bit_1237 = V_1237[quan_width-1];
assign Bit_1238 = V_1238[quan_width-1];
assign Bit_1239 = V_1239[quan_width-1];
assign Bit_1240 = V_1240[quan_width-1];
assign Bit_1241 = V_1241[quan_width-1];
assign Bit_1242 = V_1242[quan_width-1];
assign Bit_1243 = V_1243[quan_width-1];
assign Bit_1244 = V_1244[quan_width-1];
assign Bit_1245 = V_1245[quan_width-1];
assign Bit_1246 = V_1246[quan_width-1];
assign Bit_1247 = V_1247[quan_width-1];
assign Bit_1248 = V_1248[quan_width-1];
assign Bit_1249 = V_1249[quan_width-1];
assign Bit_1250 = V_1250[quan_width-1];
assign Bit_1251 = V_1251[quan_width-1];
assign Bit_1252 = V_1252[quan_width-1];
assign Bit_1253 = V_1253[quan_width-1];
assign Bit_1254 = V_1254[quan_width-1];
assign Bit_1255 = V_1255[quan_width-1];
assign Bit_1256 = V_1256[quan_width-1];
assign Bit_1257 = V_1257[quan_width-1];
assign Bit_1258 = V_1258[quan_width-1];
assign Bit_1259 = V_1259[quan_width-1];
assign Bit_1260 = V_1260[quan_width-1];
assign Bit_1261 = V_1261[quan_width-1];
assign Bit_1262 = V_1262[quan_width-1];
assign Bit_1263 = V_1263[quan_width-1];
assign Bit_1264 = V_1264[quan_width-1];
assign Bit_1265 = V_1265[quan_width-1];
assign Bit_1266 = V_1266[quan_width-1];
assign Bit_1267 = V_1267[quan_width-1];
assign Bit_1268 = V_1268[quan_width-1];
assign Bit_1269 = V_1269[quan_width-1];
assign Bit_1270 = V_1270[quan_width-1];
assign Bit_1271 = V_1271[quan_width-1];
assign Bit_1272 = V_1272[quan_width-1];
assign Bit_1273 = V_1273[quan_width-1];
assign Bit_1274 = V_1274[quan_width-1];
assign Bit_1275 = V_1275[quan_width-1];
assign Bit_1276 = V_1276[quan_width-1];
assign Bit_1277 = V_1277[quan_width-1];
assign Bit_1278 = V_1278[quan_width-1];
assign Bit_1279 = V_1279[quan_width-1];
assign Bit_1280 = V_1280[quan_width-1];
assign Bit_1281 = V_1281[quan_width-1];
assign Bit_1282 = V_1282[quan_width-1];
assign Bit_1283 = V_1283[quan_width-1];
assign Bit_1284 = V_1284[quan_width-1];
assign Bit_1285 = V_1285[quan_width-1];
assign Bit_1286 = V_1286[quan_width-1];
assign Bit_1287 = V_1287[quan_width-1];
assign Bit_1288 = V_1288[quan_width-1];
assign Bit_1289 = V_1289[quan_width-1];
assign Bit_1290 = V_1290[quan_width-1];
assign Bit_1291 = V_1291[quan_width-1];
assign Bit_1292 = V_1292[quan_width-1];
assign Bit_1293 = V_1293[quan_width-1];
assign Bit_1294 = V_1294[quan_width-1];
assign Bit_1295 = V_1295[quan_width-1];
assign Bit_1296 = V_1296[quan_width-1];
assign Bit_1297 = V_1297[quan_width-1];
assign Bit_1298 = V_1298[quan_width-1];
assign Bit_1299 = V_1299[quan_width-1];
assign Bit_1300 = V_1300[quan_width-1];
assign Bit_1301 = V_1301[quan_width-1];
assign Bit_1302 = V_1302[quan_width-1];
assign Bit_1303 = V_1303[quan_width-1];
assign Bit_1304 = V_1304[quan_width-1];
assign Bit_1305 = V_1305[quan_width-1];
assign Bit_1306 = V_1306[quan_width-1];
assign Bit_1307 = V_1307[quan_width-1];
assign Bit_1308 = V_1308[quan_width-1];
assign Bit_1309 = V_1309[quan_width-1];
assign Bit_1310 = V_1310[quan_width-1];
assign Bit_1311 = V_1311[quan_width-1];
assign Bit_1312 = V_1312[quan_width-1];
assign Bit_1313 = V_1313[quan_width-1];
assign Bit_1314 = V_1314[quan_width-1];
assign Bit_1315 = V_1315[quan_width-1];
assign Bit_1316 = V_1316[quan_width-1];
assign Bit_1317 = V_1317[quan_width-1];
assign Bit_1318 = V_1318[quan_width-1];
assign Bit_1319 = V_1319[quan_width-1];
assign Bit_1320 = V_1320[quan_width-1];
assign Bit_1321 = V_1321[quan_width-1];
assign Bit_1322 = V_1322[quan_width-1];
assign Bit_1323 = V_1323[quan_width-1];
assign Bit_1324 = V_1324[quan_width-1];
assign Bit_1325 = V_1325[quan_width-1];
assign Bit_1326 = V_1326[quan_width-1];
assign Bit_1327 = V_1327[quan_width-1];
assign Bit_1328 = V_1328[quan_width-1];
assign Bit_1329 = V_1329[quan_width-1];
assign Bit_1330 = V_1330[quan_width-1];
assign Bit_1331 = V_1331[quan_width-1];
assign Bit_1332 = V_1332[quan_width-1];
assign Bit_1333 = V_1333[quan_width-1];
assign Bit_1334 = V_1334[quan_width-1];
assign Bit_1335 = V_1335[quan_width-1];
assign Bit_1336 = V_1336[quan_width-1];
assign Bit_1337 = V_1337[quan_width-1];
assign Bit_1338 = V_1338[quan_width-1];
assign Bit_1339 = V_1339[quan_width-1];
assign Bit_1340 = V_1340[quan_width-1];
assign Bit_1341 = V_1341[quan_width-1];
assign Bit_1342 = V_1342[quan_width-1];
assign Bit_1343 = V_1343[quan_width-1];
assign Bit_1344 = V_1344[quan_width-1];
assign Bit_1345 = V_1345[quan_width-1];
assign Bit_1346 = V_1346[quan_width-1];
assign Bit_1347 = V_1347[quan_width-1];
assign Bit_1348 = V_1348[quan_width-1];
assign Bit_1349 = V_1349[quan_width-1];
assign Bit_1350 = V_1350[quan_width-1];
assign Bit_1351 = V_1351[quan_width-1];
assign Bit_1352 = V_1352[quan_width-1];
assign Bit_1353 = V_1353[quan_width-1];
assign Bit_1354 = V_1354[quan_width-1];
assign Bit_1355 = V_1355[quan_width-1];
assign Bit_1356 = V_1356[quan_width-1];
assign Bit_1357 = V_1357[quan_width-1];
assign Bit_1358 = V_1358[quan_width-1];
assign Bit_1359 = V_1359[quan_width-1];
assign Bit_1360 = V_1360[quan_width-1];
assign Bit_1361 = V_1361[quan_width-1];
assign Bit_1362 = V_1362[quan_width-1];
assign Bit_1363 = V_1363[quan_width-1];
assign Bit_1364 = V_1364[quan_width-1];
assign Bit_1365 = V_1365[quan_width-1];
assign Bit_1366 = V_1366[quan_width-1];
assign Bit_1367 = V_1367[quan_width-1];
assign Bit_1368 = V_1368[quan_width-1];
assign Bit_1369 = V_1369[quan_width-1];
assign Bit_1370 = V_1370[quan_width-1];
assign Bit_1371 = V_1371[quan_width-1];
assign Bit_1372 = V_1372[quan_width-1];
assign Bit_1373 = V_1373[quan_width-1];
assign Bit_1374 = V_1374[quan_width-1];
assign Bit_1375 = V_1375[quan_width-1];
assign Bit_1376 = V_1376[quan_width-1];
assign Bit_1377 = V_1377[quan_width-1];
assign Bit_1378 = V_1378[quan_width-1];
assign Bit_1379 = V_1379[quan_width-1];
assign Bit_1380 = V_1380[quan_width-1];
assign Bit_1381 = V_1381[quan_width-1];
assign Bit_1382 = V_1382[quan_width-1];
assign Bit_1383 = V_1383[quan_width-1];
assign Bit_1384 = V_1384[quan_width-1];
assign Bit_1385 = V_1385[quan_width-1];
assign Bit_1386 = V_1386[quan_width-1];
assign Bit_1387 = V_1387[quan_width-1];
assign Bit_1388 = V_1388[quan_width-1];
assign Bit_1389 = V_1389[quan_width-1];
assign Bit_1390 = V_1390[quan_width-1];
assign Bit_1391 = V_1391[quan_width-1];
assign Bit_1392 = V_1392[quan_width-1];
assign Bit_1393 = V_1393[quan_width-1];
assign Bit_1394 = V_1394[quan_width-1];
assign Bit_1395 = V_1395[quan_width-1];
assign Bit_1396 = V_1396[quan_width-1];
assign Bit_1397 = V_1397[quan_width-1];
assign Bit_1398 = V_1398[quan_width-1];
assign Bit_1399 = V_1399[quan_width-1];
assign Bit_1400 = V_1400[quan_width-1];
assign Bit_1401 = V_1401[quan_width-1];
assign Bit_1402 = V_1402[quan_width-1];
assign Bit_1403 = V_1403[quan_width-1];
assign Bit_1404 = V_1404[quan_width-1];
assign Bit_1405 = V_1405[quan_width-1];
assign Bit_1406 = V_1406[quan_width-1];
assign Bit_1407 = V_1407[quan_width-1];
assign Bit_1408 = V_1408[quan_width-1];
assign Bit_1409 = V_1409[quan_width-1];
assign Bit_1410 = V_1410[quan_width-1];
assign Bit_1411 = V_1411[quan_width-1];
assign Bit_1412 = V_1412[quan_width-1];
assign Bit_1413 = V_1413[quan_width-1];
assign Bit_1414 = V_1414[quan_width-1];
assign Bit_1415 = V_1415[quan_width-1];
assign Bit_1416 = V_1416[quan_width-1];
assign Bit_1417 = V_1417[quan_width-1];
assign Bit_1418 = V_1418[quan_width-1];
assign Bit_1419 = V_1419[quan_width-1];
assign Bit_1420 = V_1420[quan_width-1];
assign Bit_1421 = V_1421[quan_width-1];
assign Bit_1422 = V_1422[quan_width-1];
assign Bit_1423 = V_1423[quan_width-1];
assign Bit_1424 = V_1424[quan_width-1];
assign Bit_1425 = V_1425[quan_width-1];
assign Bit_1426 = V_1426[quan_width-1];
assign Bit_1427 = V_1427[quan_width-1];
assign Bit_1428 = V_1428[quan_width-1];
assign Bit_1429 = V_1429[quan_width-1];
assign Bit_1430 = V_1430[quan_width-1];
assign Bit_1431 = V_1431[quan_width-1];
assign Bit_1432 = V_1432[quan_width-1];
assign Bit_1433 = V_1433[quan_width-1];
assign Bit_1434 = V_1434[quan_width-1];
assign Bit_1435 = V_1435[quan_width-1];
assign Bit_1436 = V_1436[quan_width-1];
assign Bit_1437 = V_1437[quan_width-1];
assign Bit_1438 = V_1438[quan_width-1];
assign Bit_1439 = V_1439[quan_width-1];
assign Bit_1440 = V_1440[quan_width-1];

CNU_19 #(quan_width) CNU1 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_5_1),
	.V2C_2 (V2C_89_1),
	.V2C_3 (V2C_109_1),
	.V2C_4 (V2C_170_1),
	.V2C_5 (V2C_232_1),
	.V2C_6 (V2C_275_1),
	.V2C_7 (V2C_375_1),
	.V2C_8 (V2C_429_1),
	.V2C_9 (V2C_526_1),
	.V2C_10 (V2C_762_1),
	.V2C_11 (V2C_810_1),
	.V2C_12 (V2C_858_1),
	.V2C_13 (V2C_899_1),
	.V2C_14 (V2C_940_1),
	.V2C_15 (V2C_974_1),
	.V2C_16 (V2C_1013_1),
	.V2C_17 (V2C_1087_1),
	.V2C_18 (V2C_1146_1),
	.V2C_19 (V2C_1153_1),
	.C2V_1 (C2V_1_5),
	.C2V_2 (C2V_1_89),
	.C2V_3 (C2V_1_109),
	.C2V_4 (C2V_1_170),
	.C2V_5 (C2V_1_232),
	.C2V_6 (C2V_1_275),
	.C2V_7 (C2V_1_375),
	.C2V_8 (C2V_1_429),
	.C2V_9 (C2V_1_526),
	.C2V_10 (C2V_1_762),
	.C2V_11 (C2V_1_810),
	.C2V_12 (C2V_1_858),
	.C2V_13 (C2V_1_899),
	.C2V_14 (C2V_1_940),
	.C2V_15 (C2V_1_974),
	.C2V_16 (C2V_1_1013),
	.C2V_17 (C2V_1_1087),
	.C2V_18 (C2V_1_1146),
	.C2V_19 (C2V_1_1153),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU2 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_14_2),
	.V2C_2 (V2C_63_2),
	.V2C_3 (V2C_119_2),
	.V2C_4 (V2C_167_2),
	.V2C_5 (V2C_196_2),
	.V2C_6 (V2C_265_2),
	.V2C_7 (V2C_316_2),
	.V2C_8 (V2C_423_2),
	.V2C_9 (V2C_512_2),
	.V2C_10 (V2C_672_2),
	.V2C_11 (V2C_685_2),
	.V2C_12 (V2C_853_2),
	.V2C_13 (V2C_895_2),
	.V2C_14 (V2C_958_2),
	.V2C_15 (V2C_989_2),
	.V2C_16 (V2C_1021_2),
	.V2C_17 (V2C_1088_2),
	.V2C_18 (V2C_1119_2),
	.V2C_19 (V2C_1153_2),
	.V2C_20 (V2C_1154_2),
	.C2V_1 (C2V_2_14),
	.C2V_2 (C2V_2_63),
	.C2V_3 (C2V_2_119),
	.C2V_4 (C2V_2_167),
	.C2V_5 (C2V_2_196),
	.C2V_6 (C2V_2_265),
	.C2V_7 (C2V_2_316),
	.C2V_8 (C2V_2_423),
	.C2V_9 (C2V_2_512),
	.C2V_10 (C2V_2_672),
	.C2V_11 (C2V_2_685),
	.C2V_12 (C2V_2_853),
	.C2V_13 (C2V_2_895),
	.C2V_14 (C2V_2_958),
	.C2V_15 (C2V_2_989),
	.C2V_16 (C2V_2_1021),
	.C2V_17 (C2V_2_1088),
	.C2V_18 (C2V_2_1119),
	.C2V_19 (C2V_2_1153),
	.C2V_20 (C2V_2_1154),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU3 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_9_3),
	.V2C_2 (V2C_84_3),
	.V2C_3 (V2C_101_3),
	.V2C_4 (V2C_183_3),
	.V2C_5 (V2C_201_3),
	.V2C_6 (V2C_268_3),
	.V2C_7 (V2C_365_3),
	.V2C_8 (V2C_420_3),
	.V2C_9 (V2C_531_3),
	.V2C_10 (V2C_588_3),
	.V2C_11 (V2C_664_3),
	.V2C_12 (V2C_768_3),
	.V2C_13 (V2C_899_3),
	.V2C_14 (V2C_943_3),
	.V2C_15 (V2C_968_3),
	.V2C_16 (V2C_1028_3),
	.V2C_17 (V2C_1058_3),
	.V2C_18 (V2C_1151_3),
	.V2C_19 (V2C_1154_3),
	.V2C_20 (V2C_1155_3),
	.C2V_1 (C2V_3_9),
	.C2V_2 (C2V_3_84),
	.C2V_3 (C2V_3_101),
	.C2V_4 (C2V_3_183),
	.C2V_5 (C2V_3_201),
	.C2V_6 (C2V_3_268),
	.C2V_7 (C2V_3_365),
	.C2V_8 (C2V_3_420),
	.C2V_9 (C2V_3_531),
	.C2V_10 (C2V_3_588),
	.C2V_11 (C2V_3_664),
	.C2V_12 (C2V_3_768),
	.C2V_13 (C2V_3_899),
	.C2V_14 (C2V_3_943),
	.C2V_15 (C2V_3_968),
	.C2V_16 (C2V_3_1028),
	.C2V_17 (C2V_3_1058),
	.C2V_18 (C2V_3_1151),
	.C2V_19 (C2V_3_1154),
	.C2V_20 (C2V_3_1155),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU4 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_28_4),
	.V2C_2 (V2C_87_4),
	.V2C_3 (V2C_126_4),
	.V2C_4 (V2C_182_4),
	.V2C_5 (V2C_199_4),
	.V2C_6 (V2C_253_4),
	.V2C_7 (V2C_477_4),
	.V2C_8 (V2C_517_4),
	.V2C_9 (V2C_553_4),
	.V2C_10 (V2C_615_4),
	.V2C_11 (V2C_640_4),
	.V2C_12 (V2C_686_4),
	.V2C_13 (V2C_903_4),
	.V2C_14 (V2C_927_4),
	.V2C_15 (V2C_963_4),
	.V2C_16 (V2C_1041_4),
	.V2C_17 (V2C_1068_4),
	.V2C_18 (V2C_1132_4),
	.V2C_19 (V2C_1155_4),
	.V2C_20 (V2C_1156_4),
	.C2V_1 (C2V_4_28),
	.C2V_2 (C2V_4_87),
	.C2V_3 (C2V_4_126),
	.C2V_4 (C2V_4_182),
	.C2V_5 (C2V_4_199),
	.C2V_6 (C2V_4_253),
	.C2V_7 (C2V_4_477),
	.C2V_8 (C2V_4_517),
	.C2V_9 (C2V_4_553),
	.C2V_10 (C2V_4_615),
	.C2V_11 (C2V_4_640),
	.C2V_12 (C2V_4_686),
	.C2V_13 (C2V_4_903),
	.C2V_14 (C2V_4_927),
	.C2V_15 (C2V_4_963),
	.C2V_16 (C2V_4_1041),
	.C2V_17 (C2V_4_1068),
	.C2V_18 (C2V_4_1132),
	.C2V_19 (C2V_4_1155),
	.C2V_20 (C2V_4_1156),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU5 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_47_5),
	.V2C_2 (V2C_57_5),
	.V2C_3 (V2C_140_5),
	.V2C_4 (V2C_163_5),
	.V2C_5 (V2C_227_5),
	.V2C_6 (V2C_245_5),
	.V2C_7 (V2C_294_5),
	.V2C_8 (V2C_361_5),
	.V2C_9 (V2C_440_5),
	.V2C_10 (V2C_674_5),
	.V2C_11 (V2C_738_5),
	.V2C_12 (V2C_792_5),
	.V2C_13 (V2C_870_5),
	.V2C_14 (V2C_918_5),
	.V2C_15 (V2C_961_5),
	.V2C_16 (V2C_1013_5),
	.V2C_17 (V2C_1062_5),
	.V2C_18 (V2C_1110_5),
	.V2C_19 (V2C_1156_5),
	.V2C_20 (V2C_1157_5),
	.C2V_1 (C2V_5_47),
	.C2V_2 (C2V_5_57),
	.C2V_3 (C2V_5_140),
	.C2V_4 (C2V_5_163),
	.C2V_5 (C2V_5_227),
	.C2V_6 (C2V_5_245),
	.C2V_7 (C2V_5_294),
	.C2V_8 (C2V_5_361),
	.C2V_9 (C2V_5_440),
	.C2V_10 (C2V_5_674),
	.C2V_11 (C2V_5_738),
	.C2V_12 (C2V_5_792),
	.C2V_13 (C2V_5_870),
	.C2V_14 (C2V_5_918),
	.C2V_15 (C2V_5_961),
	.C2V_16 (C2V_5_1013),
	.C2V_17 (C2V_5_1062),
	.C2V_18 (C2V_5_1110),
	.C2V_19 (C2V_5_1156),
	.C2V_20 (C2V_5_1157),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU6 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_30_6),
	.V2C_2 (V2C_54_6),
	.V2C_3 (V2C_142_6),
	.V2C_4 (V2C_162_6),
	.V2C_5 (V2C_196_6),
	.V2C_6 (V2C_275_6),
	.V2C_7 (V2C_328_6),
	.V2C_8 (V2C_480_6),
	.V2C_9 (V2C_529_6),
	.V2C_10 (V2C_610_6),
	.V2C_11 (V2C_814_6),
	.V2C_12 (V2C_842_6),
	.V2C_13 (V2C_875_6),
	.V2C_14 (V2C_937_6),
	.V2C_15 (V2C_972_6),
	.V2C_16 (V2C_1039_6),
	.V2C_17 (V2C_1103_6),
	.V2C_18 (V2C_1105_6),
	.V2C_19 (V2C_1157_6),
	.V2C_20 (V2C_1158_6),
	.C2V_1 (C2V_6_30),
	.C2V_2 (C2V_6_54),
	.C2V_3 (C2V_6_142),
	.C2V_4 (C2V_6_162),
	.C2V_5 (C2V_6_196),
	.C2V_6 (C2V_6_275),
	.C2V_7 (C2V_6_328),
	.C2V_8 (C2V_6_480),
	.C2V_9 (C2V_6_529),
	.C2V_10 (C2V_6_610),
	.C2V_11 (C2V_6_814),
	.C2V_12 (C2V_6_842),
	.C2V_13 (C2V_6_875),
	.C2V_14 (C2V_6_937),
	.C2V_15 (C2V_6_972),
	.C2V_16 (C2V_6_1039),
	.C2V_17 (C2V_6_1103),
	.C2V_18 (C2V_6_1105),
	.C2V_19 (C2V_6_1157),
	.C2V_20 (C2V_6_1158),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU7 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_6_7),
	.V2C_2 (V2C_90_7),
	.V2C_3 (V2C_110_7),
	.V2C_4 (V2C_171_7),
	.V2C_5 (V2C_233_7),
	.V2C_6 (V2C_276_7),
	.V2C_7 (V2C_376_7),
	.V2C_8 (V2C_430_7),
	.V2C_9 (V2C_527_7),
	.V2C_10 (V2C_763_7),
	.V2C_11 (V2C_811_7),
	.V2C_12 (V2C_859_7),
	.V2C_13 (V2C_900_7),
	.V2C_14 (V2C_941_7),
	.V2C_15 (V2C_975_7),
	.V2C_16 (V2C_1014_7),
	.V2C_17 (V2C_1088_7),
	.V2C_18 (V2C_1147_7),
	.V2C_19 (V2C_1158_7),
	.V2C_20 (V2C_1159_7),
	.C2V_1 (C2V_7_6),
	.C2V_2 (C2V_7_90),
	.C2V_3 (C2V_7_110),
	.C2V_4 (C2V_7_171),
	.C2V_5 (C2V_7_233),
	.C2V_6 (C2V_7_276),
	.C2V_7 (C2V_7_376),
	.C2V_8 (C2V_7_430),
	.C2V_9 (C2V_7_527),
	.C2V_10 (C2V_7_763),
	.C2V_11 (C2V_7_811),
	.C2V_12 (C2V_7_859),
	.C2V_13 (C2V_7_900),
	.C2V_14 (C2V_7_941),
	.C2V_15 (C2V_7_975),
	.C2V_16 (C2V_7_1014),
	.C2V_17 (C2V_7_1088),
	.C2V_18 (C2V_7_1147),
	.C2V_19 (C2V_7_1158),
	.C2V_20 (C2V_7_1159),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU8 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_15_8),
	.V2C_2 (V2C_64_8),
	.V2C_3 (V2C_120_8),
	.V2C_4 (V2C_168_8),
	.V2C_5 (V2C_197_8),
	.V2C_6 (V2C_266_8),
	.V2C_7 (V2C_317_8),
	.V2C_8 (V2C_424_8),
	.V2C_9 (V2C_513_8),
	.V2C_10 (V2C_625_8),
	.V2C_11 (V2C_686_8),
	.V2C_12 (V2C_854_8),
	.V2C_13 (V2C_896_8),
	.V2C_14 (V2C_959_8),
	.V2C_15 (V2C_990_8),
	.V2C_16 (V2C_1022_8),
	.V2C_17 (V2C_1089_8),
	.V2C_18 (V2C_1120_8),
	.V2C_19 (V2C_1159_8),
	.V2C_20 (V2C_1160_8),
	.C2V_1 (C2V_8_15),
	.C2V_2 (C2V_8_64),
	.C2V_3 (C2V_8_120),
	.C2V_4 (C2V_8_168),
	.C2V_5 (C2V_8_197),
	.C2V_6 (C2V_8_266),
	.C2V_7 (C2V_8_317),
	.C2V_8 (C2V_8_424),
	.C2V_9 (C2V_8_513),
	.C2V_10 (C2V_8_625),
	.C2V_11 (C2V_8_686),
	.C2V_12 (C2V_8_854),
	.C2V_13 (C2V_8_896),
	.C2V_14 (C2V_8_959),
	.C2V_15 (C2V_8_990),
	.C2V_16 (C2V_8_1022),
	.C2V_17 (C2V_8_1089),
	.C2V_18 (C2V_8_1120),
	.C2V_19 (C2V_8_1159),
	.C2V_20 (C2V_8_1160),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU9 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_10_9),
	.V2C_2 (V2C_85_9),
	.V2C_3 (V2C_102_9),
	.V2C_4 (V2C_184_9),
	.V2C_5 (V2C_202_9),
	.V2C_6 (V2C_269_9),
	.V2C_7 (V2C_366_9),
	.V2C_8 (V2C_421_9),
	.V2C_9 (V2C_532_9),
	.V2C_10 (V2C_589_9),
	.V2C_11 (V2C_665_9),
	.V2C_12 (V2C_721_9),
	.V2C_13 (V2C_900_9),
	.V2C_14 (V2C_944_9),
	.V2C_15 (V2C_969_9),
	.V2C_16 (V2C_1029_9),
	.V2C_17 (V2C_1059_9),
	.V2C_18 (V2C_1152_9),
	.V2C_19 (V2C_1160_9),
	.V2C_20 (V2C_1161_9),
	.C2V_1 (C2V_9_10),
	.C2V_2 (C2V_9_85),
	.C2V_3 (C2V_9_102),
	.C2V_4 (C2V_9_184),
	.C2V_5 (C2V_9_202),
	.C2V_6 (C2V_9_269),
	.C2V_7 (C2V_9_366),
	.C2V_8 (C2V_9_421),
	.C2V_9 (C2V_9_532),
	.C2V_10 (C2V_9_589),
	.C2V_11 (C2V_9_665),
	.C2V_12 (C2V_9_721),
	.C2V_13 (C2V_9_900),
	.C2V_14 (C2V_9_944),
	.C2V_15 (C2V_9_969),
	.C2V_16 (C2V_9_1029),
	.C2V_17 (C2V_9_1059),
	.C2V_18 (C2V_9_1152),
	.C2V_19 (C2V_9_1160),
	.C2V_20 (C2V_9_1161),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU10 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_29_10),
	.V2C_2 (V2C_88_10),
	.V2C_3 (V2C_127_10),
	.V2C_4 (V2C_183_10),
	.V2C_5 (V2C_200_10),
	.V2C_6 (V2C_254_10),
	.V2C_7 (V2C_478_10),
	.V2C_8 (V2C_518_10),
	.V2C_9 (V2C_554_10),
	.V2C_10 (V2C_616_10),
	.V2C_11 (V2C_641_10),
	.V2C_12 (V2C_687_10),
	.V2C_13 (V2C_904_10),
	.V2C_14 (V2C_928_10),
	.V2C_15 (V2C_964_10),
	.V2C_16 (V2C_1042_10),
	.V2C_17 (V2C_1069_10),
	.V2C_18 (V2C_1133_10),
	.V2C_19 (V2C_1161_10),
	.V2C_20 (V2C_1162_10),
	.C2V_1 (C2V_10_29),
	.C2V_2 (C2V_10_88),
	.C2V_3 (C2V_10_127),
	.C2V_4 (C2V_10_183),
	.C2V_5 (C2V_10_200),
	.C2V_6 (C2V_10_254),
	.C2V_7 (C2V_10_478),
	.C2V_8 (C2V_10_518),
	.C2V_9 (C2V_10_554),
	.C2V_10 (C2V_10_616),
	.C2V_11 (C2V_10_641),
	.C2V_12 (C2V_10_687),
	.C2V_13 (C2V_10_904),
	.C2V_14 (C2V_10_928),
	.C2V_15 (C2V_10_964),
	.C2V_16 (C2V_10_1042),
	.C2V_17 (C2V_10_1069),
	.C2V_18 (C2V_10_1133),
	.C2V_19 (C2V_10_1161),
	.C2V_20 (C2V_10_1162),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU11 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_48_11),
	.V2C_2 (V2C_58_11),
	.V2C_3 (V2C_141_11),
	.V2C_4 (V2C_164_11),
	.V2C_5 (V2C_228_11),
	.V2C_6 (V2C_246_11),
	.V2C_7 (V2C_295_11),
	.V2C_8 (V2C_362_11),
	.V2C_9 (V2C_441_11),
	.V2C_10 (V2C_675_11),
	.V2C_11 (V2C_739_11),
	.V2C_12 (V2C_793_11),
	.V2C_13 (V2C_871_11),
	.V2C_14 (V2C_919_11),
	.V2C_15 (V2C_962_11),
	.V2C_16 (V2C_1014_11),
	.V2C_17 (V2C_1063_11),
	.V2C_18 (V2C_1111_11),
	.V2C_19 (V2C_1162_11),
	.V2C_20 (V2C_1163_11),
	.C2V_1 (C2V_11_48),
	.C2V_2 (C2V_11_58),
	.C2V_3 (C2V_11_141),
	.C2V_4 (C2V_11_164),
	.C2V_5 (C2V_11_228),
	.C2V_6 (C2V_11_246),
	.C2V_7 (C2V_11_295),
	.C2V_8 (C2V_11_362),
	.C2V_9 (C2V_11_441),
	.C2V_10 (C2V_11_675),
	.C2V_11 (C2V_11_739),
	.C2V_12 (C2V_11_793),
	.C2V_13 (C2V_11_871),
	.C2V_14 (C2V_11_919),
	.C2V_15 (C2V_11_962),
	.C2V_16 (C2V_11_1014),
	.C2V_17 (C2V_11_1063),
	.C2V_18 (C2V_11_1111),
	.C2V_19 (C2V_11_1162),
	.C2V_20 (C2V_11_1163),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU12 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_31_12),
	.V2C_2 (V2C_55_12),
	.V2C_3 (V2C_143_12),
	.V2C_4 (V2C_163_12),
	.V2C_5 (V2C_197_12),
	.V2C_6 (V2C_276_12),
	.V2C_7 (V2C_329_12),
	.V2C_8 (V2C_433_12),
	.V2C_9 (V2C_530_12),
	.V2C_10 (V2C_611_12),
	.V2C_11 (V2C_815_12),
	.V2C_12 (V2C_843_12),
	.V2C_13 (V2C_876_12),
	.V2C_14 (V2C_938_12),
	.V2C_15 (V2C_973_12),
	.V2C_16 (V2C_1040_12),
	.V2C_17 (V2C_1104_12),
	.V2C_18 (V2C_1106_12),
	.V2C_19 (V2C_1163_12),
	.V2C_20 (V2C_1164_12),
	.C2V_1 (C2V_12_31),
	.C2V_2 (C2V_12_55),
	.C2V_3 (C2V_12_143),
	.C2V_4 (C2V_12_163),
	.C2V_5 (C2V_12_197),
	.C2V_6 (C2V_12_276),
	.C2V_7 (C2V_12_329),
	.C2V_8 (C2V_12_433),
	.C2V_9 (C2V_12_530),
	.C2V_10 (C2V_12_611),
	.C2V_11 (C2V_12_815),
	.C2V_12 (C2V_12_843),
	.C2V_13 (C2V_12_876),
	.C2V_14 (C2V_12_938),
	.C2V_15 (C2V_12_973),
	.C2V_16 (C2V_12_1040),
	.C2V_17 (C2V_12_1104),
	.C2V_18 (C2V_12_1106),
	.C2V_19 (C2V_12_1163),
	.C2V_20 (C2V_12_1164),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU13 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_7_13),
	.V2C_2 (V2C_91_13),
	.V2C_3 (V2C_111_13),
	.V2C_4 (V2C_172_13),
	.V2C_5 (V2C_234_13),
	.V2C_6 (V2C_277_13),
	.V2C_7 (V2C_377_13),
	.V2C_8 (V2C_431_13),
	.V2C_9 (V2C_528_13),
	.V2C_10 (V2C_764_13),
	.V2C_11 (V2C_812_13),
	.V2C_12 (V2C_860_13),
	.V2C_13 (V2C_901_13),
	.V2C_14 (V2C_942_13),
	.V2C_15 (V2C_976_13),
	.V2C_16 (V2C_1015_13),
	.V2C_17 (V2C_1089_13),
	.V2C_18 (V2C_1148_13),
	.V2C_19 (V2C_1164_13),
	.V2C_20 (V2C_1165_13),
	.C2V_1 (C2V_13_7),
	.C2V_2 (C2V_13_91),
	.C2V_3 (C2V_13_111),
	.C2V_4 (C2V_13_172),
	.C2V_5 (C2V_13_234),
	.C2V_6 (C2V_13_277),
	.C2V_7 (C2V_13_377),
	.C2V_8 (C2V_13_431),
	.C2V_9 (C2V_13_528),
	.C2V_10 (C2V_13_764),
	.C2V_11 (C2V_13_812),
	.C2V_12 (C2V_13_860),
	.C2V_13 (C2V_13_901),
	.C2V_14 (C2V_13_942),
	.C2V_15 (C2V_13_976),
	.C2V_16 (C2V_13_1015),
	.C2V_17 (C2V_13_1089),
	.C2V_18 (C2V_13_1148),
	.C2V_19 (C2V_13_1164),
	.C2V_20 (C2V_13_1165),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU14 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_16_14),
	.V2C_2 (V2C_65_14),
	.V2C_3 (V2C_121_14),
	.V2C_4 (V2C_169_14),
	.V2C_5 (V2C_198_14),
	.V2C_6 (V2C_267_14),
	.V2C_7 (V2C_318_14),
	.V2C_8 (V2C_425_14),
	.V2C_9 (V2C_514_14),
	.V2C_10 (V2C_626_14),
	.V2C_11 (V2C_687_14),
	.V2C_12 (V2C_855_14),
	.V2C_13 (V2C_897_14),
	.V2C_14 (V2C_960_14),
	.V2C_15 (V2C_991_14),
	.V2C_16 (V2C_1023_14),
	.V2C_17 (V2C_1090_14),
	.V2C_18 (V2C_1121_14),
	.V2C_19 (V2C_1165_14),
	.V2C_20 (V2C_1166_14),
	.C2V_1 (C2V_14_16),
	.C2V_2 (C2V_14_65),
	.C2V_3 (C2V_14_121),
	.C2V_4 (C2V_14_169),
	.C2V_5 (C2V_14_198),
	.C2V_6 (C2V_14_267),
	.C2V_7 (C2V_14_318),
	.C2V_8 (C2V_14_425),
	.C2V_9 (C2V_14_514),
	.C2V_10 (C2V_14_626),
	.C2V_11 (C2V_14_687),
	.C2V_12 (C2V_14_855),
	.C2V_13 (C2V_14_897),
	.C2V_14 (C2V_14_960),
	.C2V_15 (C2V_14_991),
	.C2V_16 (C2V_14_1023),
	.C2V_17 (C2V_14_1090),
	.C2V_18 (C2V_14_1121),
	.C2V_19 (C2V_14_1165),
	.C2V_20 (C2V_14_1166),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU15 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_11_15),
	.V2C_2 (V2C_86_15),
	.V2C_3 (V2C_103_15),
	.V2C_4 (V2C_185_15),
	.V2C_5 (V2C_203_15),
	.V2C_6 (V2C_270_15),
	.V2C_7 (V2C_367_15),
	.V2C_8 (V2C_422_15),
	.V2C_9 (V2C_533_15),
	.V2C_10 (V2C_590_15),
	.V2C_11 (V2C_666_15),
	.V2C_12 (V2C_722_15),
	.V2C_13 (V2C_901_15),
	.V2C_14 (V2C_945_15),
	.V2C_15 (V2C_970_15),
	.V2C_16 (V2C_1030_15),
	.V2C_17 (V2C_1060_15),
	.V2C_18 (V2C_1105_15),
	.V2C_19 (V2C_1166_15),
	.V2C_20 (V2C_1167_15),
	.C2V_1 (C2V_15_11),
	.C2V_2 (C2V_15_86),
	.C2V_3 (C2V_15_103),
	.C2V_4 (C2V_15_185),
	.C2V_5 (C2V_15_203),
	.C2V_6 (C2V_15_270),
	.C2V_7 (C2V_15_367),
	.C2V_8 (C2V_15_422),
	.C2V_9 (C2V_15_533),
	.C2V_10 (C2V_15_590),
	.C2V_11 (C2V_15_666),
	.C2V_12 (C2V_15_722),
	.C2V_13 (C2V_15_901),
	.C2V_14 (C2V_15_945),
	.C2V_15 (C2V_15_970),
	.C2V_16 (C2V_15_1030),
	.C2V_17 (C2V_15_1060),
	.C2V_18 (C2V_15_1105),
	.C2V_19 (C2V_15_1166),
	.C2V_20 (C2V_15_1167),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU16 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_30_16),
	.V2C_2 (V2C_89_16),
	.V2C_3 (V2C_128_16),
	.V2C_4 (V2C_184_16),
	.V2C_5 (V2C_201_16),
	.V2C_6 (V2C_255_16),
	.V2C_7 (V2C_479_16),
	.V2C_8 (V2C_519_16),
	.V2C_9 (V2C_555_16),
	.V2C_10 (V2C_617_16),
	.V2C_11 (V2C_642_16),
	.V2C_12 (V2C_688_16),
	.V2C_13 (V2C_905_16),
	.V2C_14 (V2C_929_16),
	.V2C_15 (V2C_965_16),
	.V2C_16 (V2C_1043_16),
	.V2C_17 (V2C_1070_16),
	.V2C_18 (V2C_1134_16),
	.V2C_19 (V2C_1167_16),
	.V2C_20 (V2C_1168_16),
	.C2V_1 (C2V_16_30),
	.C2V_2 (C2V_16_89),
	.C2V_3 (C2V_16_128),
	.C2V_4 (C2V_16_184),
	.C2V_5 (C2V_16_201),
	.C2V_6 (C2V_16_255),
	.C2V_7 (C2V_16_479),
	.C2V_8 (C2V_16_519),
	.C2V_9 (C2V_16_555),
	.C2V_10 (C2V_16_617),
	.C2V_11 (C2V_16_642),
	.C2V_12 (C2V_16_688),
	.C2V_13 (C2V_16_905),
	.C2V_14 (C2V_16_929),
	.C2V_15 (C2V_16_965),
	.C2V_16 (C2V_16_1043),
	.C2V_17 (C2V_16_1070),
	.C2V_18 (C2V_16_1134),
	.C2V_19 (C2V_16_1167),
	.C2V_20 (C2V_16_1168),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU17 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_1_17),
	.V2C_2 (V2C_59_17),
	.V2C_3 (V2C_142_17),
	.V2C_4 (V2C_165_17),
	.V2C_5 (V2C_229_17),
	.V2C_6 (V2C_247_17),
	.V2C_7 (V2C_296_17),
	.V2C_8 (V2C_363_17),
	.V2C_9 (V2C_442_17),
	.V2C_10 (V2C_676_17),
	.V2C_11 (V2C_740_17),
	.V2C_12 (V2C_794_17),
	.V2C_13 (V2C_872_17),
	.V2C_14 (V2C_920_17),
	.V2C_15 (V2C_963_17),
	.V2C_16 (V2C_1015_17),
	.V2C_17 (V2C_1064_17),
	.V2C_18 (V2C_1112_17),
	.V2C_19 (V2C_1168_17),
	.V2C_20 (V2C_1169_17),
	.C2V_1 (C2V_17_1),
	.C2V_2 (C2V_17_59),
	.C2V_3 (C2V_17_142),
	.C2V_4 (C2V_17_165),
	.C2V_5 (C2V_17_229),
	.C2V_6 (C2V_17_247),
	.C2V_7 (C2V_17_296),
	.C2V_8 (C2V_17_363),
	.C2V_9 (C2V_17_442),
	.C2V_10 (C2V_17_676),
	.C2V_11 (C2V_17_740),
	.C2V_12 (C2V_17_794),
	.C2V_13 (C2V_17_872),
	.C2V_14 (C2V_17_920),
	.C2V_15 (C2V_17_963),
	.C2V_16 (C2V_17_1015),
	.C2V_17 (C2V_17_1064),
	.C2V_18 (C2V_17_1112),
	.C2V_19 (C2V_17_1168),
	.C2V_20 (C2V_17_1169),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU18 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_32_18),
	.V2C_2 (V2C_56_18),
	.V2C_3 (V2C_144_18),
	.V2C_4 (V2C_164_18),
	.V2C_5 (V2C_198_18),
	.V2C_6 (V2C_277_18),
	.V2C_7 (V2C_330_18),
	.V2C_8 (V2C_434_18),
	.V2C_9 (V2C_531_18),
	.V2C_10 (V2C_612_18),
	.V2C_11 (V2C_816_18),
	.V2C_12 (V2C_844_18),
	.V2C_13 (V2C_877_18),
	.V2C_14 (V2C_939_18),
	.V2C_15 (V2C_974_18),
	.V2C_16 (V2C_1041_18),
	.V2C_17 (V2C_1057_18),
	.V2C_18 (V2C_1107_18),
	.V2C_19 (V2C_1169_18),
	.V2C_20 (V2C_1170_18),
	.C2V_1 (C2V_18_32),
	.C2V_2 (C2V_18_56),
	.C2V_3 (C2V_18_144),
	.C2V_4 (C2V_18_164),
	.C2V_5 (C2V_18_198),
	.C2V_6 (C2V_18_277),
	.C2V_7 (C2V_18_330),
	.C2V_8 (C2V_18_434),
	.C2V_9 (C2V_18_531),
	.C2V_10 (C2V_18_612),
	.C2V_11 (C2V_18_816),
	.C2V_12 (C2V_18_844),
	.C2V_13 (C2V_18_877),
	.C2V_14 (C2V_18_939),
	.C2V_15 (C2V_18_974),
	.C2V_16 (C2V_18_1041),
	.C2V_17 (C2V_18_1057),
	.C2V_18 (C2V_18_1107),
	.C2V_19 (C2V_18_1169),
	.C2V_20 (C2V_18_1170),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU19 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_8_19),
	.V2C_2 (V2C_92_19),
	.V2C_3 (V2C_112_19),
	.V2C_4 (V2C_173_19),
	.V2C_5 (V2C_235_19),
	.V2C_6 (V2C_278_19),
	.V2C_7 (V2C_378_19),
	.V2C_8 (V2C_432_19),
	.V2C_9 (V2C_481_19),
	.V2C_10 (V2C_765_19),
	.V2C_11 (V2C_813_19),
	.V2C_12 (V2C_861_19),
	.V2C_13 (V2C_902_19),
	.V2C_14 (V2C_943_19),
	.V2C_15 (V2C_977_19),
	.V2C_16 (V2C_1016_19),
	.V2C_17 (V2C_1090_19),
	.V2C_18 (V2C_1149_19),
	.V2C_19 (V2C_1170_19),
	.V2C_20 (V2C_1171_19),
	.C2V_1 (C2V_19_8),
	.C2V_2 (C2V_19_92),
	.C2V_3 (C2V_19_112),
	.C2V_4 (C2V_19_173),
	.C2V_5 (C2V_19_235),
	.C2V_6 (C2V_19_278),
	.C2V_7 (C2V_19_378),
	.C2V_8 (C2V_19_432),
	.C2V_9 (C2V_19_481),
	.C2V_10 (C2V_19_765),
	.C2V_11 (C2V_19_813),
	.C2V_12 (C2V_19_861),
	.C2V_13 (C2V_19_902),
	.C2V_14 (C2V_19_943),
	.C2V_15 (C2V_19_977),
	.C2V_16 (C2V_19_1016),
	.C2V_17 (C2V_19_1090),
	.C2V_18 (C2V_19_1149),
	.C2V_19 (C2V_19_1170),
	.C2V_20 (C2V_19_1171),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU20 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_17_20),
	.V2C_2 (V2C_66_20),
	.V2C_3 (V2C_122_20),
	.V2C_4 (V2C_170_20),
	.V2C_5 (V2C_199_20),
	.V2C_6 (V2C_268_20),
	.V2C_7 (V2C_319_20),
	.V2C_8 (V2C_426_20),
	.V2C_9 (V2C_515_20),
	.V2C_10 (V2C_627_20),
	.V2C_11 (V2C_688_20),
	.V2C_12 (V2C_856_20),
	.V2C_13 (V2C_898_20),
	.V2C_14 (V2C_913_20),
	.V2C_15 (V2C_992_20),
	.V2C_16 (V2C_1024_20),
	.V2C_17 (V2C_1091_20),
	.V2C_18 (V2C_1122_20),
	.V2C_19 (V2C_1171_20),
	.V2C_20 (V2C_1172_20),
	.C2V_1 (C2V_20_17),
	.C2V_2 (C2V_20_66),
	.C2V_3 (C2V_20_122),
	.C2V_4 (C2V_20_170),
	.C2V_5 (C2V_20_199),
	.C2V_6 (C2V_20_268),
	.C2V_7 (C2V_20_319),
	.C2V_8 (C2V_20_426),
	.C2V_9 (C2V_20_515),
	.C2V_10 (C2V_20_627),
	.C2V_11 (C2V_20_688),
	.C2V_12 (C2V_20_856),
	.C2V_13 (C2V_20_898),
	.C2V_14 (C2V_20_913),
	.C2V_15 (C2V_20_992),
	.C2V_16 (C2V_20_1024),
	.C2V_17 (C2V_20_1091),
	.C2V_18 (C2V_20_1122),
	.C2V_19 (C2V_20_1171),
	.C2V_20 (C2V_20_1172),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU21 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_12_21),
	.V2C_2 (V2C_87_21),
	.V2C_3 (V2C_104_21),
	.V2C_4 (V2C_186_21),
	.V2C_5 (V2C_204_21),
	.V2C_6 (V2C_271_21),
	.V2C_7 (V2C_368_21),
	.V2C_8 (V2C_423_21),
	.V2C_9 (V2C_534_21),
	.V2C_10 (V2C_591_21),
	.V2C_11 (V2C_667_21),
	.V2C_12 (V2C_723_21),
	.V2C_13 (V2C_902_21),
	.V2C_14 (V2C_946_21),
	.V2C_15 (V2C_971_21),
	.V2C_16 (V2C_1031_21),
	.V2C_17 (V2C_1061_21),
	.V2C_18 (V2C_1106_21),
	.V2C_19 (V2C_1172_21),
	.V2C_20 (V2C_1173_21),
	.C2V_1 (C2V_21_12),
	.C2V_2 (C2V_21_87),
	.C2V_3 (C2V_21_104),
	.C2V_4 (C2V_21_186),
	.C2V_5 (C2V_21_204),
	.C2V_6 (C2V_21_271),
	.C2V_7 (C2V_21_368),
	.C2V_8 (C2V_21_423),
	.C2V_9 (C2V_21_534),
	.C2V_10 (C2V_21_591),
	.C2V_11 (C2V_21_667),
	.C2V_12 (C2V_21_723),
	.C2V_13 (C2V_21_902),
	.C2V_14 (C2V_21_946),
	.C2V_15 (C2V_21_971),
	.C2V_16 (C2V_21_1031),
	.C2V_17 (C2V_21_1061),
	.C2V_18 (C2V_21_1106),
	.C2V_19 (C2V_21_1172),
	.C2V_20 (C2V_21_1173),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU22 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_31_22),
	.V2C_2 (V2C_90_22),
	.V2C_3 (V2C_129_22),
	.V2C_4 (V2C_185_22),
	.V2C_5 (V2C_202_22),
	.V2C_6 (V2C_256_22),
	.V2C_7 (V2C_480_22),
	.V2C_8 (V2C_520_22),
	.V2C_9 (V2C_556_22),
	.V2C_10 (V2C_618_22),
	.V2C_11 (V2C_643_22),
	.V2C_12 (V2C_689_22),
	.V2C_13 (V2C_906_22),
	.V2C_14 (V2C_930_22),
	.V2C_15 (V2C_966_22),
	.V2C_16 (V2C_1044_22),
	.V2C_17 (V2C_1071_22),
	.V2C_18 (V2C_1135_22),
	.V2C_19 (V2C_1173_22),
	.V2C_20 (V2C_1174_22),
	.C2V_1 (C2V_22_31),
	.C2V_2 (C2V_22_90),
	.C2V_3 (C2V_22_129),
	.C2V_4 (C2V_22_185),
	.C2V_5 (C2V_22_202),
	.C2V_6 (C2V_22_256),
	.C2V_7 (C2V_22_480),
	.C2V_8 (C2V_22_520),
	.C2V_9 (C2V_22_556),
	.C2V_10 (C2V_22_618),
	.C2V_11 (C2V_22_643),
	.C2V_12 (C2V_22_689),
	.C2V_13 (C2V_22_906),
	.C2V_14 (C2V_22_930),
	.C2V_15 (C2V_22_966),
	.C2V_16 (C2V_22_1044),
	.C2V_17 (C2V_22_1071),
	.C2V_18 (C2V_22_1135),
	.C2V_19 (C2V_22_1173),
	.C2V_20 (C2V_22_1174),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU23 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_2_23),
	.V2C_2 (V2C_60_23),
	.V2C_3 (V2C_143_23),
	.V2C_4 (V2C_166_23),
	.V2C_5 (V2C_230_23),
	.V2C_6 (V2C_248_23),
	.V2C_7 (V2C_297_23),
	.V2C_8 (V2C_364_23),
	.V2C_9 (V2C_443_23),
	.V2C_10 (V2C_677_23),
	.V2C_11 (V2C_741_23),
	.V2C_12 (V2C_795_23),
	.V2C_13 (V2C_873_23),
	.V2C_14 (V2C_921_23),
	.V2C_15 (V2C_964_23),
	.V2C_16 (V2C_1016_23),
	.V2C_17 (V2C_1065_23),
	.V2C_18 (V2C_1113_23),
	.V2C_19 (V2C_1174_23),
	.V2C_20 (V2C_1175_23),
	.C2V_1 (C2V_23_2),
	.C2V_2 (C2V_23_60),
	.C2V_3 (C2V_23_143),
	.C2V_4 (C2V_23_166),
	.C2V_5 (C2V_23_230),
	.C2V_6 (C2V_23_248),
	.C2V_7 (C2V_23_297),
	.C2V_8 (C2V_23_364),
	.C2V_9 (C2V_23_443),
	.C2V_10 (C2V_23_677),
	.C2V_11 (C2V_23_741),
	.C2V_12 (C2V_23_795),
	.C2V_13 (C2V_23_873),
	.C2V_14 (C2V_23_921),
	.C2V_15 (C2V_23_964),
	.C2V_16 (C2V_23_1016),
	.C2V_17 (C2V_23_1065),
	.C2V_18 (C2V_23_1113),
	.C2V_19 (C2V_23_1174),
	.C2V_20 (C2V_23_1175),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU24 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_33_24),
	.V2C_2 (V2C_57_24),
	.V2C_3 (V2C_97_24),
	.V2C_4 (V2C_165_24),
	.V2C_5 (V2C_199_24),
	.V2C_6 (V2C_278_24),
	.V2C_7 (V2C_331_24),
	.V2C_8 (V2C_435_24),
	.V2C_9 (V2C_532_24),
	.V2C_10 (V2C_613_24),
	.V2C_11 (V2C_769_24),
	.V2C_12 (V2C_845_24),
	.V2C_13 (V2C_878_24),
	.V2C_14 (V2C_940_24),
	.V2C_15 (V2C_975_24),
	.V2C_16 (V2C_1042_24),
	.V2C_17 (V2C_1058_24),
	.V2C_18 (V2C_1108_24),
	.V2C_19 (V2C_1175_24),
	.V2C_20 (V2C_1176_24),
	.C2V_1 (C2V_24_33),
	.C2V_2 (C2V_24_57),
	.C2V_3 (C2V_24_97),
	.C2V_4 (C2V_24_165),
	.C2V_5 (C2V_24_199),
	.C2V_6 (C2V_24_278),
	.C2V_7 (C2V_24_331),
	.C2V_8 (C2V_24_435),
	.C2V_9 (C2V_24_532),
	.C2V_10 (C2V_24_613),
	.C2V_11 (C2V_24_769),
	.C2V_12 (C2V_24_845),
	.C2V_13 (C2V_24_878),
	.C2V_14 (C2V_24_940),
	.C2V_15 (C2V_24_975),
	.C2V_16 (C2V_24_1042),
	.C2V_17 (C2V_24_1058),
	.C2V_18 (C2V_24_1108),
	.C2V_19 (C2V_24_1175),
	.C2V_20 (C2V_24_1176),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU25 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_9_25),
	.V2C_2 (V2C_93_25),
	.V2C_3 (V2C_113_25),
	.V2C_4 (V2C_174_25),
	.V2C_5 (V2C_236_25),
	.V2C_6 (V2C_279_25),
	.V2C_7 (V2C_379_25),
	.V2C_8 (V2C_385_25),
	.V2C_9 (V2C_482_25),
	.V2C_10 (V2C_766_25),
	.V2C_11 (V2C_814_25),
	.V2C_12 (V2C_862_25),
	.V2C_13 (V2C_903_25),
	.V2C_14 (V2C_944_25),
	.V2C_15 (V2C_978_25),
	.V2C_16 (V2C_1017_25),
	.V2C_17 (V2C_1091_25),
	.V2C_18 (V2C_1150_25),
	.V2C_19 (V2C_1176_25),
	.V2C_20 (V2C_1177_25),
	.C2V_1 (C2V_25_9),
	.C2V_2 (C2V_25_93),
	.C2V_3 (C2V_25_113),
	.C2V_4 (C2V_25_174),
	.C2V_5 (C2V_25_236),
	.C2V_6 (C2V_25_279),
	.C2V_7 (C2V_25_379),
	.C2V_8 (C2V_25_385),
	.C2V_9 (C2V_25_482),
	.C2V_10 (C2V_25_766),
	.C2V_11 (C2V_25_814),
	.C2V_12 (C2V_25_862),
	.C2V_13 (C2V_25_903),
	.C2V_14 (C2V_25_944),
	.C2V_15 (C2V_25_978),
	.C2V_16 (C2V_25_1017),
	.C2V_17 (C2V_25_1091),
	.C2V_18 (C2V_25_1150),
	.C2V_19 (C2V_25_1176),
	.C2V_20 (C2V_25_1177),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU26 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_18_26),
	.V2C_2 (V2C_67_26),
	.V2C_3 (V2C_123_26),
	.V2C_4 (V2C_171_26),
	.V2C_5 (V2C_200_26),
	.V2C_6 (V2C_269_26),
	.V2C_7 (V2C_320_26),
	.V2C_8 (V2C_427_26),
	.V2C_9 (V2C_516_26),
	.V2C_10 (V2C_628_26),
	.V2C_11 (V2C_689_26),
	.V2C_12 (V2C_857_26),
	.V2C_13 (V2C_899_26),
	.V2C_14 (V2C_914_26),
	.V2C_15 (V2C_993_26),
	.V2C_16 (V2C_1025_26),
	.V2C_17 (V2C_1092_26),
	.V2C_18 (V2C_1123_26),
	.V2C_19 (V2C_1177_26),
	.V2C_20 (V2C_1178_26),
	.C2V_1 (C2V_26_18),
	.C2V_2 (C2V_26_67),
	.C2V_3 (C2V_26_123),
	.C2V_4 (C2V_26_171),
	.C2V_5 (C2V_26_200),
	.C2V_6 (C2V_26_269),
	.C2V_7 (C2V_26_320),
	.C2V_8 (C2V_26_427),
	.C2V_9 (C2V_26_516),
	.C2V_10 (C2V_26_628),
	.C2V_11 (C2V_26_689),
	.C2V_12 (C2V_26_857),
	.C2V_13 (C2V_26_899),
	.C2V_14 (C2V_26_914),
	.C2V_15 (C2V_26_993),
	.C2V_16 (C2V_26_1025),
	.C2V_17 (C2V_26_1092),
	.C2V_18 (C2V_26_1123),
	.C2V_19 (C2V_26_1177),
	.C2V_20 (C2V_26_1178),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU27 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_13_27),
	.V2C_2 (V2C_88_27),
	.V2C_3 (V2C_105_27),
	.V2C_4 (V2C_187_27),
	.V2C_5 (V2C_205_27),
	.V2C_6 (V2C_272_27),
	.V2C_7 (V2C_369_27),
	.V2C_8 (V2C_424_27),
	.V2C_9 (V2C_535_27),
	.V2C_10 (V2C_592_27),
	.V2C_11 (V2C_668_27),
	.V2C_12 (V2C_724_27),
	.V2C_13 (V2C_903_27),
	.V2C_14 (V2C_947_27),
	.V2C_15 (V2C_972_27),
	.V2C_16 (V2C_1032_27),
	.V2C_17 (V2C_1062_27),
	.V2C_18 (V2C_1107_27),
	.V2C_19 (V2C_1178_27),
	.V2C_20 (V2C_1179_27),
	.C2V_1 (C2V_27_13),
	.C2V_2 (C2V_27_88),
	.C2V_3 (C2V_27_105),
	.C2V_4 (C2V_27_187),
	.C2V_5 (C2V_27_205),
	.C2V_6 (C2V_27_272),
	.C2V_7 (C2V_27_369),
	.C2V_8 (C2V_27_424),
	.C2V_9 (C2V_27_535),
	.C2V_10 (C2V_27_592),
	.C2V_11 (C2V_27_668),
	.C2V_12 (C2V_27_724),
	.C2V_13 (C2V_27_903),
	.C2V_14 (C2V_27_947),
	.C2V_15 (C2V_27_972),
	.C2V_16 (C2V_27_1032),
	.C2V_17 (C2V_27_1062),
	.C2V_18 (C2V_27_1107),
	.C2V_19 (C2V_27_1178),
	.C2V_20 (C2V_27_1179),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU28 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_32_28),
	.V2C_2 (V2C_91_28),
	.V2C_3 (V2C_130_28),
	.V2C_4 (V2C_186_28),
	.V2C_5 (V2C_203_28),
	.V2C_6 (V2C_257_28),
	.V2C_7 (V2C_433_28),
	.V2C_8 (V2C_521_28),
	.V2C_9 (V2C_557_28),
	.V2C_10 (V2C_619_28),
	.V2C_11 (V2C_644_28),
	.V2C_12 (V2C_690_28),
	.V2C_13 (V2C_907_28),
	.V2C_14 (V2C_931_28),
	.V2C_15 (V2C_967_28),
	.V2C_16 (V2C_1045_28),
	.V2C_17 (V2C_1072_28),
	.V2C_18 (V2C_1136_28),
	.V2C_19 (V2C_1179_28),
	.V2C_20 (V2C_1180_28),
	.C2V_1 (C2V_28_32),
	.C2V_2 (C2V_28_91),
	.C2V_3 (C2V_28_130),
	.C2V_4 (C2V_28_186),
	.C2V_5 (C2V_28_203),
	.C2V_6 (C2V_28_257),
	.C2V_7 (C2V_28_433),
	.C2V_8 (C2V_28_521),
	.C2V_9 (C2V_28_557),
	.C2V_10 (C2V_28_619),
	.C2V_11 (C2V_28_644),
	.C2V_12 (C2V_28_690),
	.C2V_13 (C2V_28_907),
	.C2V_14 (C2V_28_931),
	.C2V_15 (C2V_28_967),
	.C2V_16 (C2V_28_1045),
	.C2V_17 (C2V_28_1072),
	.C2V_18 (C2V_28_1136),
	.C2V_19 (C2V_28_1179),
	.C2V_20 (C2V_28_1180),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU29 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_3_29),
	.V2C_2 (V2C_61_29),
	.V2C_3 (V2C_144_29),
	.V2C_4 (V2C_167_29),
	.V2C_5 (V2C_231_29),
	.V2C_6 (V2C_249_29),
	.V2C_7 (V2C_298_29),
	.V2C_8 (V2C_365_29),
	.V2C_9 (V2C_444_29),
	.V2C_10 (V2C_678_29),
	.V2C_11 (V2C_742_29),
	.V2C_12 (V2C_796_29),
	.V2C_13 (V2C_874_29),
	.V2C_14 (V2C_922_29),
	.V2C_15 (V2C_965_29),
	.V2C_16 (V2C_1017_29),
	.V2C_17 (V2C_1066_29),
	.V2C_18 (V2C_1114_29),
	.V2C_19 (V2C_1180_29),
	.V2C_20 (V2C_1181_29),
	.C2V_1 (C2V_29_3),
	.C2V_2 (C2V_29_61),
	.C2V_3 (C2V_29_144),
	.C2V_4 (C2V_29_167),
	.C2V_5 (C2V_29_231),
	.C2V_6 (C2V_29_249),
	.C2V_7 (C2V_29_298),
	.C2V_8 (C2V_29_365),
	.C2V_9 (C2V_29_444),
	.C2V_10 (C2V_29_678),
	.C2V_11 (C2V_29_742),
	.C2V_12 (C2V_29_796),
	.C2V_13 (C2V_29_874),
	.C2V_14 (C2V_29_922),
	.C2V_15 (C2V_29_965),
	.C2V_16 (C2V_29_1017),
	.C2V_17 (C2V_29_1066),
	.C2V_18 (C2V_29_1114),
	.C2V_19 (C2V_29_1180),
	.C2V_20 (C2V_29_1181),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU30 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_34_30),
	.V2C_2 (V2C_58_30),
	.V2C_3 (V2C_98_30),
	.V2C_4 (V2C_166_30),
	.V2C_5 (V2C_200_30),
	.V2C_6 (V2C_279_30),
	.V2C_7 (V2C_332_30),
	.V2C_8 (V2C_436_30),
	.V2C_9 (V2C_533_30),
	.V2C_10 (V2C_614_30),
	.V2C_11 (V2C_770_30),
	.V2C_12 (V2C_846_30),
	.V2C_13 (V2C_879_30),
	.V2C_14 (V2C_941_30),
	.V2C_15 (V2C_976_30),
	.V2C_16 (V2C_1043_30),
	.V2C_17 (V2C_1059_30),
	.V2C_18 (V2C_1109_30),
	.V2C_19 (V2C_1181_30),
	.V2C_20 (V2C_1182_30),
	.C2V_1 (C2V_30_34),
	.C2V_2 (C2V_30_58),
	.C2V_3 (C2V_30_98),
	.C2V_4 (C2V_30_166),
	.C2V_5 (C2V_30_200),
	.C2V_6 (C2V_30_279),
	.C2V_7 (C2V_30_332),
	.C2V_8 (C2V_30_436),
	.C2V_9 (C2V_30_533),
	.C2V_10 (C2V_30_614),
	.C2V_11 (C2V_30_770),
	.C2V_12 (C2V_30_846),
	.C2V_13 (C2V_30_879),
	.C2V_14 (C2V_30_941),
	.C2V_15 (C2V_30_976),
	.C2V_16 (C2V_30_1043),
	.C2V_17 (C2V_30_1059),
	.C2V_18 (C2V_30_1109),
	.C2V_19 (C2V_30_1181),
	.C2V_20 (C2V_30_1182),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU31 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_10_31),
	.V2C_2 (V2C_94_31),
	.V2C_3 (V2C_114_31),
	.V2C_4 (V2C_175_31),
	.V2C_5 (V2C_237_31),
	.V2C_6 (V2C_280_31),
	.V2C_7 (V2C_380_31),
	.V2C_8 (V2C_386_31),
	.V2C_9 (V2C_483_31),
	.V2C_10 (V2C_767_31),
	.V2C_11 (V2C_815_31),
	.V2C_12 (V2C_863_31),
	.V2C_13 (V2C_904_31),
	.V2C_14 (V2C_945_31),
	.V2C_15 (V2C_979_31),
	.V2C_16 (V2C_1018_31),
	.V2C_17 (V2C_1092_31),
	.V2C_18 (V2C_1151_31),
	.V2C_19 (V2C_1182_31),
	.V2C_20 (V2C_1183_31),
	.C2V_1 (C2V_31_10),
	.C2V_2 (C2V_31_94),
	.C2V_3 (C2V_31_114),
	.C2V_4 (C2V_31_175),
	.C2V_5 (C2V_31_237),
	.C2V_6 (C2V_31_280),
	.C2V_7 (C2V_31_380),
	.C2V_8 (C2V_31_386),
	.C2V_9 (C2V_31_483),
	.C2V_10 (C2V_31_767),
	.C2V_11 (C2V_31_815),
	.C2V_12 (C2V_31_863),
	.C2V_13 (C2V_31_904),
	.C2V_14 (C2V_31_945),
	.C2V_15 (C2V_31_979),
	.C2V_16 (C2V_31_1018),
	.C2V_17 (C2V_31_1092),
	.C2V_18 (C2V_31_1151),
	.C2V_19 (C2V_31_1182),
	.C2V_20 (C2V_31_1183),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU32 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_19_32),
	.V2C_2 (V2C_68_32),
	.V2C_3 (V2C_124_32),
	.V2C_4 (V2C_172_32),
	.V2C_5 (V2C_201_32),
	.V2C_6 (V2C_270_32),
	.V2C_7 (V2C_321_32),
	.V2C_8 (V2C_428_32),
	.V2C_9 (V2C_517_32),
	.V2C_10 (V2C_629_32),
	.V2C_11 (V2C_690_32),
	.V2C_12 (V2C_858_32),
	.V2C_13 (V2C_900_32),
	.V2C_14 (V2C_915_32),
	.V2C_15 (V2C_994_32),
	.V2C_16 (V2C_1026_32),
	.V2C_17 (V2C_1093_32),
	.V2C_18 (V2C_1124_32),
	.V2C_19 (V2C_1183_32),
	.V2C_20 (V2C_1184_32),
	.C2V_1 (C2V_32_19),
	.C2V_2 (C2V_32_68),
	.C2V_3 (C2V_32_124),
	.C2V_4 (C2V_32_172),
	.C2V_5 (C2V_32_201),
	.C2V_6 (C2V_32_270),
	.C2V_7 (C2V_32_321),
	.C2V_8 (C2V_32_428),
	.C2V_9 (C2V_32_517),
	.C2V_10 (C2V_32_629),
	.C2V_11 (C2V_32_690),
	.C2V_12 (C2V_32_858),
	.C2V_13 (C2V_32_900),
	.C2V_14 (C2V_32_915),
	.C2V_15 (C2V_32_994),
	.C2V_16 (C2V_32_1026),
	.C2V_17 (C2V_32_1093),
	.C2V_18 (C2V_32_1124),
	.C2V_19 (C2V_32_1183),
	.C2V_20 (C2V_32_1184),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU33 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_14_33),
	.V2C_2 (V2C_89_33),
	.V2C_3 (V2C_106_33),
	.V2C_4 (V2C_188_33),
	.V2C_5 (V2C_206_33),
	.V2C_6 (V2C_273_33),
	.V2C_7 (V2C_370_33),
	.V2C_8 (V2C_425_33),
	.V2C_9 (V2C_536_33),
	.V2C_10 (V2C_593_33),
	.V2C_11 (V2C_669_33),
	.V2C_12 (V2C_725_33),
	.V2C_13 (V2C_904_33),
	.V2C_14 (V2C_948_33),
	.V2C_15 (V2C_973_33),
	.V2C_16 (V2C_1033_33),
	.V2C_17 (V2C_1063_33),
	.V2C_18 (V2C_1108_33),
	.V2C_19 (V2C_1184_33),
	.V2C_20 (V2C_1185_33),
	.C2V_1 (C2V_33_14),
	.C2V_2 (C2V_33_89),
	.C2V_3 (C2V_33_106),
	.C2V_4 (C2V_33_188),
	.C2V_5 (C2V_33_206),
	.C2V_6 (C2V_33_273),
	.C2V_7 (C2V_33_370),
	.C2V_8 (C2V_33_425),
	.C2V_9 (C2V_33_536),
	.C2V_10 (C2V_33_593),
	.C2V_11 (C2V_33_669),
	.C2V_12 (C2V_33_725),
	.C2V_13 (C2V_33_904),
	.C2V_14 (C2V_33_948),
	.C2V_15 (C2V_33_973),
	.C2V_16 (C2V_33_1033),
	.C2V_17 (C2V_33_1063),
	.C2V_18 (C2V_33_1108),
	.C2V_19 (C2V_33_1184),
	.C2V_20 (C2V_33_1185),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU34 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_33_34),
	.V2C_2 (V2C_92_34),
	.V2C_3 (V2C_131_34),
	.V2C_4 (V2C_187_34),
	.V2C_5 (V2C_204_34),
	.V2C_6 (V2C_258_34),
	.V2C_7 (V2C_434_34),
	.V2C_8 (V2C_522_34),
	.V2C_9 (V2C_558_34),
	.V2C_10 (V2C_620_34),
	.V2C_11 (V2C_645_34),
	.V2C_12 (V2C_691_34),
	.V2C_13 (V2C_908_34),
	.V2C_14 (V2C_932_34),
	.V2C_15 (V2C_968_34),
	.V2C_16 (V2C_1046_34),
	.V2C_17 (V2C_1073_34),
	.V2C_18 (V2C_1137_34),
	.V2C_19 (V2C_1185_34),
	.V2C_20 (V2C_1186_34),
	.C2V_1 (C2V_34_33),
	.C2V_2 (C2V_34_92),
	.C2V_3 (C2V_34_131),
	.C2V_4 (C2V_34_187),
	.C2V_5 (C2V_34_204),
	.C2V_6 (C2V_34_258),
	.C2V_7 (C2V_34_434),
	.C2V_8 (C2V_34_522),
	.C2V_9 (C2V_34_558),
	.C2V_10 (C2V_34_620),
	.C2V_11 (C2V_34_645),
	.C2V_12 (C2V_34_691),
	.C2V_13 (C2V_34_908),
	.C2V_14 (C2V_34_932),
	.C2V_15 (C2V_34_968),
	.C2V_16 (C2V_34_1046),
	.C2V_17 (C2V_34_1073),
	.C2V_18 (C2V_34_1137),
	.C2V_19 (C2V_34_1185),
	.C2V_20 (C2V_34_1186),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU35 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_4_35),
	.V2C_2 (V2C_62_35),
	.V2C_3 (V2C_97_35),
	.V2C_4 (V2C_168_35),
	.V2C_5 (V2C_232_35),
	.V2C_6 (V2C_250_35),
	.V2C_7 (V2C_299_35),
	.V2C_8 (V2C_366_35),
	.V2C_9 (V2C_445_35),
	.V2C_10 (V2C_679_35),
	.V2C_11 (V2C_743_35),
	.V2C_12 (V2C_797_35),
	.V2C_13 (V2C_875_35),
	.V2C_14 (V2C_923_35),
	.V2C_15 (V2C_966_35),
	.V2C_16 (V2C_1018_35),
	.V2C_17 (V2C_1067_35),
	.V2C_18 (V2C_1115_35),
	.V2C_19 (V2C_1186_35),
	.V2C_20 (V2C_1187_35),
	.C2V_1 (C2V_35_4),
	.C2V_2 (C2V_35_62),
	.C2V_3 (C2V_35_97),
	.C2V_4 (C2V_35_168),
	.C2V_5 (C2V_35_232),
	.C2V_6 (C2V_35_250),
	.C2V_7 (C2V_35_299),
	.C2V_8 (C2V_35_366),
	.C2V_9 (C2V_35_445),
	.C2V_10 (C2V_35_679),
	.C2V_11 (C2V_35_743),
	.C2V_12 (C2V_35_797),
	.C2V_13 (C2V_35_875),
	.C2V_14 (C2V_35_923),
	.C2V_15 (C2V_35_966),
	.C2V_16 (C2V_35_1018),
	.C2V_17 (C2V_35_1067),
	.C2V_18 (C2V_35_1115),
	.C2V_19 (C2V_35_1186),
	.C2V_20 (C2V_35_1187),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU36 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_35_36),
	.V2C_2 (V2C_59_36),
	.V2C_3 (V2C_99_36),
	.V2C_4 (V2C_167_36),
	.V2C_5 (V2C_201_36),
	.V2C_6 (V2C_280_36),
	.V2C_7 (V2C_333_36),
	.V2C_8 (V2C_437_36),
	.V2C_9 (V2C_534_36),
	.V2C_10 (V2C_615_36),
	.V2C_11 (V2C_771_36),
	.V2C_12 (V2C_847_36),
	.V2C_13 (V2C_880_36),
	.V2C_14 (V2C_942_36),
	.V2C_15 (V2C_977_36),
	.V2C_16 (V2C_1044_36),
	.V2C_17 (V2C_1060_36),
	.V2C_18 (V2C_1110_36),
	.V2C_19 (V2C_1187_36),
	.V2C_20 (V2C_1188_36),
	.C2V_1 (C2V_36_35),
	.C2V_2 (C2V_36_59),
	.C2V_3 (C2V_36_99),
	.C2V_4 (C2V_36_167),
	.C2V_5 (C2V_36_201),
	.C2V_6 (C2V_36_280),
	.C2V_7 (C2V_36_333),
	.C2V_8 (C2V_36_437),
	.C2V_9 (C2V_36_534),
	.C2V_10 (C2V_36_615),
	.C2V_11 (C2V_36_771),
	.C2V_12 (C2V_36_847),
	.C2V_13 (C2V_36_880),
	.C2V_14 (C2V_36_942),
	.C2V_15 (C2V_36_977),
	.C2V_16 (C2V_36_1044),
	.C2V_17 (C2V_36_1060),
	.C2V_18 (C2V_36_1110),
	.C2V_19 (C2V_36_1187),
	.C2V_20 (C2V_36_1188),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU37 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_11_37),
	.V2C_2 (V2C_95_37),
	.V2C_3 (V2C_115_37),
	.V2C_4 (V2C_176_37),
	.V2C_5 (V2C_238_37),
	.V2C_6 (V2C_281_37),
	.V2C_7 (V2C_381_37),
	.V2C_8 (V2C_387_37),
	.V2C_9 (V2C_484_37),
	.V2C_10 (V2C_768_37),
	.V2C_11 (V2C_816_37),
	.V2C_12 (V2C_864_37),
	.V2C_13 (V2C_905_37),
	.V2C_14 (V2C_946_37),
	.V2C_15 (V2C_980_37),
	.V2C_16 (V2C_1019_37),
	.V2C_17 (V2C_1093_37),
	.V2C_18 (V2C_1152_37),
	.V2C_19 (V2C_1188_37),
	.V2C_20 (V2C_1189_37),
	.C2V_1 (C2V_37_11),
	.C2V_2 (C2V_37_95),
	.C2V_3 (C2V_37_115),
	.C2V_4 (C2V_37_176),
	.C2V_5 (C2V_37_238),
	.C2V_6 (C2V_37_281),
	.C2V_7 (C2V_37_381),
	.C2V_8 (C2V_37_387),
	.C2V_9 (C2V_37_484),
	.C2V_10 (C2V_37_768),
	.C2V_11 (C2V_37_816),
	.C2V_12 (C2V_37_864),
	.C2V_13 (C2V_37_905),
	.C2V_14 (C2V_37_946),
	.C2V_15 (C2V_37_980),
	.C2V_16 (C2V_37_1019),
	.C2V_17 (C2V_37_1093),
	.C2V_18 (C2V_37_1152),
	.C2V_19 (C2V_37_1188),
	.C2V_20 (C2V_37_1189),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU38 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_20_38),
	.V2C_2 (V2C_69_38),
	.V2C_3 (V2C_125_38),
	.V2C_4 (V2C_173_38),
	.V2C_5 (V2C_202_38),
	.V2C_6 (V2C_271_38),
	.V2C_7 (V2C_322_38),
	.V2C_8 (V2C_429_38),
	.V2C_9 (V2C_518_38),
	.V2C_10 (V2C_630_38),
	.V2C_11 (V2C_691_38),
	.V2C_12 (V2C_859_38),
	.V2C_13 (V2C_901_38),
	.V2C_14 (V2C_916_38),
	.V2C_15 (V2C_995_38),
	.V2C_16 (V2C_1027_38),
	.V2C_17 (V2C_1094_38),
	.V2C_18 (V2C_1125_38),
	.V2C_19 (V2C_1189_38),
	.V2C_20 (V2C_1190_38),
	.C2V_1 (C2V_38_20),
	.C2V_2 (C2V_38_69),
	.C2V_3 (C2V_38_125),
	.C2V_4 (C2V_38_173),
	.C2V_5 (C2V_38_202),
	.C2V_6 (C2V_38_271),
	.C2V_7 (C2V_38_322),
	.C2V_8 (C2V_38_429),
	.C2V_9 (C2V_38_518),
	.C2V_10 (C2V_38_630),
	.C2V_11 (C2V_38_691),
	.C2V_12 (C2V_38_859),
	.C2V_13 (C2V_38_901),
	.C2V_14 (C2V_38_916),
	.C2V_15 (C2V_38_995),
	.C2V_16 (C2V_38_1027),
	.C2V_17 (C2V_38_1094),
	.C2V_18 (C2V_38_1125),
	.C2V_19 (C2V_38_1189),
	.C2V_20 (C2V_38_1190),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU39 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_15_39),
	.V2C_2 (V2C_90_39),
	.V2C_3 (V2C_107_39),
	.V2C_4 (V2C_189_39),
	.V2C_5 (V2C_207_39),
	.V2C_6 (V2C_274_39),
	.V2C_7 (V2C_371_39),
	.V2C_8 (V2C_426_39),
	.V2C_9 (V2C_537_39),
	.V2C_10 (V2C_594_39),
	.V2C_11 (V2C_670_39),
	.V2C_12 (V2C_726_39),
	.V2C_13 (V2C_905_39),
	.V2C_14 (V2C_949_39),
	.V2C_15 (V2C_974_39),
	.V2C_16 (V2C_1034_39),
	.V2C_17 (V2C_1064_39),
	.V2C_18 (V2C_1109_39),
	.V2C_19 (V2C_1190_39),
	.V2C_20 (V2C_1191_39),
	.C2V_1 (C2V_39_15),
	.C2V_2 (C2V_39_90),
	.C2V_3 (C2V_39_107),
	.C2V_4 (C2V_39_189),
	.C2V_5 (C2V_39_207),
	.C2V_6 (C2V_39_274),
	.C2V_7 (C2V_39_371),
	.C2V_8 (C2V_39_426),
	.C2V_9 (C2V_39_537),
	.C2V_10 (C2V_39_594),
	.C2V_11 (C2V_39_670),
	.C2V_12 (C2V_39_726),
	.C2V_13 (C2V_39_905),
	.C2V_14 (C2V_39_949),
	.C2V_15 (C2V_39_974),
	.C2V_16 (C2V_39_1034),
	.C2V_17 (C2V_39_1064),
	.C2V_18 (C2V_39_1109),
	.C2V_19 (C2V_39_1190),
	.C2V_20 (C2V_39_1191),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU40 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_34_40),
	.V2C_2 (V2C_93_40),
	.V2C_3 (V2C_132_40),
	.V2C_4 (V2C_188_40),
	.V2C_5 (V2C_205_40),
	.V2C_6 (V2C_259_40),
	.V2C_7 (V2C_435_40),
	.V2C_8 (V2C_523_40),
	.V2C_9 (V2C_559_40),
	.V2C_10 (V2C_621_40),
	.V2C_11 (V2C_646_40),
	.V2C_12 (V2C_692_40),
	.V2C_13 (V2C_909_40),
	.V2C_14 (V2C_933_40),
	.V2C_15 (V2C_969_40),
	.V2C_16 (V2C_1047_40),
	.V2C_17 (V2C_1074_40),
	.V2C_18 (V2C_1138_40),
	.V2C_19 (V2C_1191_40),
	.V2C_20 (V2C_1192_40),
	.C2V_1 (C2V_40_34),
	.C2V_2 (C2V_40_93),
	.C2V_3 (C2V_40_132),
	.C2V_4 (C2V_40_188),
	.C2V_5 (C2V_40_205),
	.C2V_6 (C2V_40_259),
	.C2V_7 (C2V_40_435),
	.C2V_8 (C2V_40_523),
	.C2V_9 (C2V_40_559),
	.C2V_10 (C2V_40_621),
	.C2V_11 (C2V_40_646),
	.C2V_12 (C2V_40_692),
	.C2V_13 (C2V_40_909),
	.C2V_14 (C2V_40_933),
	.C2V_15 (C2V_40_969),
	.C2V_16 (C2V_40_1047),
	.C2V_17 (C2V_40_1074),
	.C2V_18 (C2V_40_1138),
	.C2V_19 (C2V_40_1191),
	.C2V_20 (C2V_40_1192),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU41 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_5_41),
	.V2C_2 (V2C_63_41),
	.V2C_3 (V2C_98_41),
	.V2C_4 (V2C_169_41),
	.V2C_5 (V2C_233_41),
	.V2C_6 (V2C_251_41),
	.V2C_7 (V2C_300_41),
	.V2C_8 (V2C_367_41),
	.V2C_9 (V2C_446_41),
	.V2C_10 (V2C_680_41),
	.V2C_11 (V2C_744_41),
	.V2C_12 (V2C_798_41),
	.V2C_13 (V2C_876_41),
	.V2C_14 (V2C_924_41),
	.V2C_15 (V2C_967_41),
	.V2C_16 (V2C_1019_41),
	.V2C_17 (V2C_1068_41),
	.V2C_18 (V2C_1116_41),
	.V2C_19 (V2C_1192_41),
	.V2C_20 (V2C_1193_41),
	.C2V_1 (C2V_41_5),
	.C2V_2 (C2V_41_63),
	.C2V_3 (C2V_41_98),
	.C2V_4 (C2V_41_169),
	.C2V_5 (C2V_41_233),
	.C2V_6 (C2V_41_251),
	.C2V_7 (C2V_41_300),
	.C2V_8 (C2V_41_367),
	.C2V_9 (C2V_41_446),
	.C2V_10 (C2V_41_680),
	.C2V_11 (C2V_41_744),
	.C2V_12 (C2V_41_798),
	.C2V_13 (C2V_41_876),
	.C2V_14 (C2V_41_924),
	.C2V_15 (C2V_41_967),
	.C2V_16 (C2V_41_1019),
	.C2V_17 (C2V_41_1068),
	.C2V_18 (C2V_41_1116),
	.C2V_19 (C2V_41_1192),
	.C2V_20 (C2V_41_1193),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU42 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_36_42),
	.V2C_2 (V2C_60_42),
	.V2C_3 (V2C_100_42),
	.V2C_4 (V2C_168_42),
	.V2C_5 (V2C_202_42),
	.V2C_6 (V2C_281_42),
	.V2C_7 (V2C_334_42),
	.V2C_8 (V2C_438_42),
	.V2C_9 (V2C_535_42),
	.V2C_10 (V2C_616_42),
	.V2C_11 (V2C_772_42),
	.V2C_12 (V2C_848_42),
	.V2C_13 (V2C_881_42),
	.V2C_14 (V2C_943_42),
	.V2C_15 (V2C_978_42),
	.V2C_16 (V2C_1045_42),
	.V2C_17 (V2C_1061_42),
	.V2C_18 (V2C_1111_42),
	.V2C_19 (V2C_1193_42),
	.V2C_20 (V2C_1194_42),
	.C2V_1 (C2V_42_36),
	.C2V_2 (C2V_42_60),
	.C2V_3 (C2V_42_100),
	.C2V_4 (C2V_42_168),
	.C2V_5 (C2V_42_202),
	.C2V_6 (C2V_42_281),
	.C2V_7 (C2V_42_334),
	.C2V_8 (C2V_42_438),
	.C2V_9 (C2V_42_535),
	.C2V_10 (C2V_42_616),
	.C2V_11 (C2V_42_772),
	.C2V_12 (C2V_42_848),
	.C2V_13 (C2V_42_881),
	.C2V_14 (C2V_42_943),
	.C2V_15 (C2V_42_978),
	.C2V_16 (C2V_42_1045),
	.C2V_17 (C2V_42_1061),
	.C2V_18 (C2V_42_1111),
	.C2V_19 (C2V_42_1193),
	.C2V_20 (C2V_42_1194),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU43 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_12_43),
	.V2C_2 (V2C_96_43),
	.V2C_3 (V2C_116_43),
	.V2C_4 (V2C_177_43),
	.V2C_5 (V2C_239_43),
	.V2C_6 (V2C_282_43),
	.V2C_7 (V2C_382_43),
	.V2C_8 (V2C_388_43),
	.V2C_9 (V2C_485_43),
	.V2C_10 (V2C_721_43),
	.V2C_11 (V2C_769_43),
	.V2C_12 (V2C_817_43),
	.V2C_13 (V2C_906_43),
	.V2C_14 (V2C_947_43),
	.V2C_15 (V2C_981_43),
	.V2C_16 (V2C_1020_43),
	.V2C_17 (V2C_1094_43),
	.V2C_18 (V2C_1105_43),
	.V2C_19 (V2C_1194_43),
	.V2C_20 (V2C_1195_43),
	.C2V_1 (C2V_43_12),
	.C2V_2 (C2V_43_96),
	.C2V_3 (C2V_43_116),
	.C2V_4 (C2V_43_177),
	.C2V_5 (C2V_43_239),
	.C2V_6 (C2V_43_282),
	.C2V_7 (C2V_43_382),
	.C2V_8 (C2V_43_388),
	.C2V_9 (C2V_43_485),
	.C2V_10 (C2V_43_721),
	.C2V_11 (C2V_43_769),
	.C2V_12 (C2V_43_817),
	.C2V_13 (C2V_43_906),
	.C2V_14 (C2V_43_947),
	.C2V_15 (C2V_43_981),
	.C2V_16 (C2V_43_1020),
	.C2V_17 (C2V_43_1094),
	.C2V_18 (C2V_43_1105),
	.C2V_19 (C2V_43_1194),
	.C2V_20 (C2V_43_1195),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU44 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_21_44),
	.V2C_2 (V2C_70_44),
	.V2C_3 (V2C_126_44),
	.V2C_4 (V2C_174_44),
	.V2C_5 (V2C_203_44),
	.V2C_6 (V2C_272_44),
	.V2C_7 (V2C_323_44),
	.V2C_8 (V2C_430_44),
	.V2C_9 (V2C_519_44),
	.V2C_10 (V2C_631_44),
	.V2C_11 (V2C_692_44),
	.V2C_12 (V2C_860_44),
	.V2C_13 (V2C_902_44),
	.V2C_14 (V2C_917_44),
	.V2C_15 (V2C_996_44),
	.V2C_16 (V2C_1028_44),
	.V2C_17 (V2C_1095_44),
	.V2C_18 (V2C_1126_44),
	.V2C_19 (V2C_1195_44),
	.V2C_20 (V2C_1196_44),
	.C2V_1 (C2V_44_21),
	.C2V_2 (C2V_44_70),
	.C2V_3 (C2V_44_126),
	.C2V_4 (C2V_44_174),
	.C2V_5 (C2V_44_203),
	.C2V_6 (C2V_44_272),
	.C2V_7 (C2V_44_323),
	.C2V_8 (C2V_44_430),
	.C2V_9 (C2V_44_519),
	.C2V_10 (C2V_44_631),
	.C2V_11 (C2V_44_692),
	.C2V_12 (C2V_44_860),
	.C2V_13 (C2V_44_902),
	.C2V_14 (C2V_44_917),
	.C2V_15 (C2V_44_996),
	.C2V_16 (C2V_44_1028),
	.C2V_17 (C2V_44_1095),
	.C2V_18 (C2V_44_1126),
	.C2V_19 (C2V_44_1195),
	.C2V_20 (C2V_44_1196),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU45 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_16_45),
	.V2C_2 (V2C_91_45),
	.V2C_3 (V2C_108_45),
	.V2C_4 (V2C_190_45),
	.V2C_5 (V2C_208_45),
	.V2C_6 (V2C_275_45),
	.V2C_7 (V2C_372_45),
	.V2C_8 (V2C_427_45),
	.V2C_9 (V2C_538_45),
	.V2C_10 (V2C_595_45),
	.V2C_11 (V2C_671_45),
	.V2C_12 (V2C_727_45),
	.V2C_13 (V2C_906_45),
	.V2C_14 (V2C_950_45),
	.V2C_15 (V2C_975_45),
	.V2C_16 (V2C_1035_45),
	.V2C_17 (V2C_1065_45),
	.V2C_18 (V2C_1110_45),
	.V2C_19 (V2C_1196_45),
	.V2C_20 (V2C_1197_45),
	.C2V_1 (C2V_45_16),
	.C2V_2 (C2V_45_91),
	.C2V_3 (C2V_45_108),
	.C2V_4 (C2V_45_190),
	.C2V_5 (C2V_45_208),
	.C2V_6 (C2V_45_275),
	.C2V_7 (C2V_45_372),
	.C2V_8 (C2V_45_427),
	.C2V_9 (C2V_45_538),
	.C2V_10 (C2V_45_595),
	.C2V_11 (C2V_45_671),
	.C2V_12 (C2V_45_727),
	.C2V_13 (C2V_45_906),
	.C2V_14 (C2V_45_950),
	.C2V_15 (C2V_45_975),
	.C2V_16 (C2V_45_1035),
	.C2V_17 (C2V_45_1065),
	.C2V_18 (C2V_45_1110),
	.C2V_19 (C2V_45_1196),
	.C2V_20 (C2V_45_1197),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU46 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_35_46),
	.V2C_2 (V2C_94_46),
	.V2C_3 (V2C_133_46),
	.V2C_4 (V2C_189_46),
	.V2C_5 (V2C_206_46),
	.V2C_6 (V2C_260_46),
	.V2C_7 (V2C_436_46),
	.V2C_8 (V2C_524_46),
	.V2C_9 (V2C_560_46),
	.V2C_10 (V2C_622_46),
	.V2C_11 (V2C_647_46),
	.V2C_12 (V2C_693_46),
	.V2C_13 (V2C_910_46),
	.V2C_14 (V2C_934_46),
	.V2C_15 (V2C_970_46),
	.V2C_16 (V2C_1048_46),
	.V2C_17 (V2C_1075_46),
	.V2C_18 (V2C_1139_46),
	.V2C_19 (V2C_1197_46),
	.V2C_20 (V2C_1198_46),
	.C2V_1 (C2V_46_35),
	.C2V_2 (C2V_46_94),
	.C2V_3 (C2V_46_133),
	.C2V_4 (C2V_46_189),
	.C2V_5 (C2V_46_206),
	.C2V_6 (C2V_46_260),
	.C2V_7 (C2V_46_436),
	.C2V_8 (C2V_46_524),
	.C2V_9 (C2V_46_560),
	.C2V_10 (C2V_46_622),
	.C2V_11 (C2V_46_647),
	.C2V_12 (C2V_46_693),
	.C2V_13 (C2V_46_910),
	.C2V_14 (C2V_46_934),
	.C2V_15 (C2V_46_970),
	.C2V_16 (C2V_46_1048),
	.C2V_17 (C2V_46_1075),
	.C2V_18 (C2V_46_1139),
	.C2V_19 (C2V_46_1197),
	.C2V_20 (C2V_46_1198),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU47 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_6_47),
	.V2C_2 (V2C_64_47),
	.V2C_3 (V2C_99_47),
	.V2C_4 (V2C_170_47),
	.V2C_5 (V2C_234_47),
	.V2C_6 (V2C_252_47),
	.V2C_7 (V2C_301_47),
	.V2C_8 (V2C_368_47),
	.V2C_9 (V2C_447_47),
	.V2C_10 (V2C_681_47),
	.V2C_11 (V2C_745_47),
	.V2C_12 (V2C_799_47),
	.V2C_13 (V2C_877_47),
	.V2C_14 (V2C_925_47),
	.V2C_15 (V2C_968_47),
	.V2C_16 (V2C_1020_47),
	.V2C_17 (V2C_1069_47),
	.V2C_18 (V2C_1117_47),
	.V2C_19 (V2C_1198_47),
	.V2C_20 (V2C_1199_47),
	.C2V_1 (C2V_47_6),
	.C2V_2 (C2V_47_64),
	.C2V_3 (C2V_47_99),
	.C2V_4 (C2V_47_170),
	.C2V_5 (C2V_47_234),
	.C2V_6 (C2V_47_252),
	.C2V_7 (C2V_47_301),
	.C2V_8 (C2V_47_368),
	.C2V_9 (C2V_47_447),
	.C2V_10 (C2V_47_681),
	.C2V_11 (C2V_47_745),
	.C2V_12 (C2V_47_799),
	.C2V_13 (C2V_47_877),
	.C2V_14 (C2V_47_925),
	.C2V_15 (C2V_47_968),
	.C2V_16 (C2V_47_1020),
	.C2V_17 (C2V_47_1069),
	.C2V_18 (C2V_47_1117),
	.C2V_19 (C2V_47_1198),
	.C2V_20 (C2V_47_1199),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU48 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_37_48),
	.V2C_2 (V2C_61_48),
	.V2C_3 (V2C_101_48),
	.V2C_4 (V2C_169_48),
	.V2C_5 (V2C_203_48),
	.V2C_6 (V2C_282_48),
	.V2C_7 (V2C_335_48),
	.V2C_8 (V2C_439_48),
	.V2C_9 (V2C_536_48),
	.V2C_10 (V2C_617_48),
	.V2C_11 (V2C_773_48),
	.V2C_12 (V2C_849_48),
	.V2C_13 (V2C_882_48),
	.V2C_14 (V2C_944_48),
	.V2C_15 (V2C_979_48),
	.V2C_16 (V2C_1046_48),
	.V2C_17 (V2C_1062_48),
	.V2C_18 (V2C_1112_48),
	.V2C_19 (V2C_1199_48),
	.V2C_20 (V2C_1200_48),
	.C2V_1 (C2V_48_37),
	.C2V_2 (C2V_48_61),
	.C2V_3 (C2V_48_101),
	.C2V_4 (C2V_48_169),
	.C2V_5 (C2V_48_203),
	.C2V_6 (C2V_48_282),
	.C2V_7 (C2V_48_335),
	.C2V_8 (C2V_48_439),
	.C2V_9 (C2V_48_536),
	.C2V_10 (C2V_48_617),
	.C2V_11 (C2V_48_773),
	.C2V_12 (C2V_48_849),
	.C2V_13 (C2V_48_882),
	.C2V_14 (C2V_48_944),
	.C2V_15 (C2V_48_979),
	.C2V_16 (C2V_48_1046),
	.C2V_17 (C2V_48_1062),
	.C2V_18 (C2V_48_1112),
	.C2V_19 (C2V_48_1199),
	.C2V_20 (C2V_48_1200),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU49 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_13_49),
	.V2C_2 (V2C_49_49),
	.V2C_3 (V2C_117_49),
	.V2C_4 (V2C_178_49),
	.V2C_5 (V2C_240_49),
	.V2C_6 (V2C_283_49),
	.V2C_7 (V2C_383_49),
	.V2C_8 (V2C_389_49),
	.V2C_9 (V2C_486_49),
	.V2C_10 (V2C_722_49),
	.V2C_11 (V2C_770_49),
	.V2C_12 (V2C_818_49),
	.V2C_13 (V2C_907_49),
	.V2C_14 (V2C_948_49),
	.V2C_15 (V2C_982_49),
	.V2C_16 (V2C_1021_49),
	.V2C_17 (V2C_1095_49),
	.V2C_18 (V2C_1106_49),
	.V2C_19 (V2C_1200_49),
	.V2C_20 (V2C_1201_49),
	.C2V_1 (C2V_49_13),
	.C2V_2 (C2V_49_49),
	.C2V_3 (C2V_49_117),
	.C2V_4 (C2V_49_178),
	.C2V_5 (C2V_49_240),
	.C2V_6 (C2V_49_283),
	.C2V_7 (C2V_49_383),
	.C2V_8 (C2V_49_389),
	.C2V_9 (C2V_49_486),
	.C2V_10 (C2V_49_722),
	.C2V_11 (C2V_49_770),
	.C2V_12 (C2V_49_818),
	.C2V_13 (C2V_49_907),
	.C2V_14 (C2V_49_948),
	.C2V_15 (C2V_49_982),
	.C2V_16 (C2V_49_1021),
	.C2V_17 (C2V_49_1095),
	.C2V_18 (C2V_49_1106),
	.C2V_19 (C2V_49_1200),
	.C2V_20 (C2V_49_1201),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU50 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_22_50),
	.V2C_2 (V2C_71_50),
	.V2C_3 (V2C_127_50),
	.V2C_4 (V2C_175_50),
	.V2C_5 (V2C_204_50),
	.V2C_6 (V2C_273_50),
	.V2C_7 (V2C_324_50),
	.V2C_8 (V2C_431_50),
	.V2C_9 (V2C_520_50),
	.V2C_10 (V2C_632_50),
	.V2C_11 (V2C_693_50),
	.V2C_12 (V2C_861_50),
	.V2C_13 (V2C_903_50),
	.V2C_14 (V2C_918_50),
	.V2C_15 (V2C_997_50),
	.V2C_16 (V2C_1029_50),
	.V2C_17 (V2C_1096_50),
	.V2C_18 (V2C_1127_50),
	.V2C_19 (V2C_1201_50),
	.V2C_20 (V2C_1202_50),
	.C2V_1 (C2V_50_22),
	.C2V_2 (C2V_50_71),
	.C2V_3 (C2V_50_127),
	.C2V_4 (C2V_50_175),
	.C2V_5 (C2V_50_204),
	.C2V_6 (C2V_50_273),
	.C2V_7 (C2V_50_324),
	.C2V_8 (C2V_50_431),
	.C2V_9 (C2V_50_520),
	.C2V_10 (C2V_50_632),
	.C2V_11 (C2V_50_693),
	.C2V_12 (C2V_50_861),
	.C2V_13 (C2V_50_903),
	.C2V_14 (C2V_50_918),
	.C2V_15 (C2V_50_997),
	.C2V_16 (C2V_50_1029),
	.C2V_17 (C2V_50_1096),
	.C2V_18 (C2V_50_1127),
	.C2V_19 (C2V_50_1201),
	.C2V_20 (C2V_50_1202),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU51 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_17_51),
	.V2C_2 (V2C_92_51),
	.V2C_3 (V2C_109_51),
	.V2C_4 (V2C_191_51),
	.V2C_5 (V2C_209_51),
	.V2C_6 (V2C_276_51),
	.V2C_7 (V2C_373_51),
	.V2C_8 (V2C_428_51),
	.V2C_9 (V2C_539_51),
	.V2C_10 (V2C_596_51),
	.V2C_11 (V2C_672_51),
	.V2C_12 (V2C_728_51),
	.V2C_13 (V2C_907_51),
	.V2C_14 (V2C_951_51),
	.V2C_15 (V2C_976_51),
	.V2C_16 (V2C_1036_51),
	.V2C_17 (V2C_1066_51),
	.V2C_18 (V2C_1111_51),
	.V2C_19 (V2C_1202_51),
	.V2C_20 (V2C_1203_51),
	.C2V_1 (C2V_51_17),
	.C2V_2 (C2V_51_92),
	.C2V_3 (C2V_51_109),
	.C2V_4 (C2V_51_191),
	.C2V_5 (C2V_51_209),
	.C2V_6 (C2V_51_276),
	.C2V_7 (C2V_51_373),
	.C2V_8 (C2V_51_428),
	.C2V_9 (C2V_51_539),
	.C2V_10 (C2V_51_596),
	.C2V_11 (C2V_51_672),
	.C2V_12 (C2V_51_728),
	.C2V_13 (C2V_51_907),
	.C2V_14 (C2V_51_951),
	.C2V_15 (C2V_51_976),
	.C2V_16 (C2V_51_1036),
	.C2V_17 (C2V_51_1066),
	.C2V_18 (C2V_51_1111),
	.C2V_19 (C2V_51_1202),
	.C2V_20 (C2V_51_1203),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU52 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_36_52),
	.V2C_2 (V2C_95_52),
	.V2C_3 (V2C_134_52),
	.V2C_4 (V2C_190_52),
	.V2C_5 (V2C_207_52),
	.V2C_6 (V2C_261_52),
	.V2C_7 (V2C_437_52),
	.V2C_8 (V2C_525_52),
	.V2C_9 (V2C_561_52),
	.V2C_10 (V2C_623_52),
	.V2C_11 (V2C_648_52),
	.V2C_12 (V2C_694_52),
	.V2C_13 (V2C_911_52),
	.V2C_14 (V2C_935_52),
	.V2C_15 (V2C_971_52),
	.V2C_16 (V2C_1049_52),
	.V2C_17 (V2C_1076_52),
	.V2C_18 (V2C_1140_52),
	.V2C_19 (V2C_1203_52),
	.V2C_20 (V2C_1204_52),
	.C2V_1 (C2V_52_36),
	.C2V_2 (C2V_52_95),
	.C2V_3 (C2V_52_134),
	.C2V_4 (C2V_52_190),
	.C2V_5 (C2V_52_207),
	.C2V_6 (C2V_52_261),
	.C2V_7 (C2V_52_437),
	.C2V_8 (C2V_52_525),
	.C2V_9 (C2V_52_561),
	.C2V_10 (C2V_52_623),
	.C2V_11 (C2V_52_648),
	.C2V_12 (C2V_52_694),
	.C2V_13 (C2V_52_911),
	.C2V_14 (C2V_52_935),
	.C2V_15 (C2V_52_971),
	.C2V_16 (C2V_52_1049),
	.C2V_17 (C2V_52_1076),
	.C2V_18 (C2V_52_1140),
	.C2V_19 (C2V_52_1203),
	.C2V_20 (C2V_52_1204),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU53 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_7_53),
	.V2C_2 (V2C_65_53),
	.V2C_3 (V2C_100_53),
	.V2C_4 (V2C_171_53),
	.V2C_5 (V2C_235_53),
	.V2C_6 (V2C_253_53),
	.V2C_7 (V2C_302_53),
	.V2C_8 (V2C_369_53),
	.V2C_9 (V2C_448_53),
	.V2C_10 (V2C_682_53),
	.V2C_11 (V2C_746_53),
	.V2C_12 (V2C_800_53),
	.V2C_13 (V2C_878_53),
	.V2C_14 (V2C_926_53),
	.V2C_15 (V2C_969_53),
	.V2C_16 (V2C_1021_53),
	.V2C_17 (V2C_1070_53),
	.V2C_18 (V2C_1118_53),
	.V2C_19 (V2C_1204_53),
	.V2C_20 (V2C_1205_53),
	.C2V_1 (C2V_53_7),
	.C2V_2 (C2V_53_65),
	.C2V_3 (C2V_53_100),
	.C2V_4 (C2V_53_171),
	.C2V_5 (C2V_53_235),
	.C2V_6 (C2V_53_253),
	.C2V_7 (C2V_53_302),
	.C2V_8 (C2V_53_369),
	.C2V_9 (C2V_53_448),
	.C2V_10 (C2V_53_682),
	.C2V_11 (C2V_53_746),
	.C2V_12 (C2V_53_800),
	.C2V_13 (C2V_53_878),
	.C2V_14 (C2V_53_926),
	.C2V_15 (C2V_53_969),
	.C2V_16 (C2V_53_1021),
	.C2V_17 (C2V_53_1070),
	.C2V_18 (C2V_53_1118),
	.C2V_19 (C2V_53_1204),
	.C2V_20 (C2V_53_1205),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU54 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_38_54),
	.V2C_2 (V2C_62_54),
	.V2C_3 (V2C_102_54),
	.V2C_4 (V2C_170_54),
	.V2C_5 (V2C_204_54),
	.V2C_6 (V2C_283_54),
	.V2C_7 (V2C_336_54),
	.V2C_8 (V2C_440_54),
	.V2C_9 (V2C_537_54),
	.V2C_10 (V2C_618_54),
	.V2C_11 (V2C_774_54),
	.V2C_12 (V2C_850_54),
	.V2C_13 (V2C_883_54),
	.V2C_14 (V2C_945_54),
	.V2C_15 (V2C_980_54),
	.V2C_16 (V2C_1047_54),
	.V2C_17 (V2C_1063_54),
	.V2C_18 (V2C_1113_54),
	.V2C_19 (V2C_1205_54),
	.V2C_20 (V2C_1206_54),
	.C2V_1 (C2V_54_38),
	.C2V_2 (C2V_54_62),
	.C2V_3 (C2V_54_102),
	.C2V_4 (C2V_54_170),
	.C2V_5 (C2V_54_204),
	.C2V_6 (C2V_54_283),
	.C2V_7 (C2V_54_336),
	.C2V_8 (C2V_54_440),
	.C2V_9 (C2V_54_537),
	.C2V_10 (C2V_54_618),
	.C2V_11 (C2V_54_774),
	.C2V_12 (C2V_54_850),
	.C2V_13 (C2V_54_883),
	.C2V_14 (C2V_54_945),
	.C2V_15 (C2V_54_980),
	.C2V_16 (C2V_54_1047),
	.C2V_17 (C2V_54_1063),
	.C2V_18 (C2V_54_1113),
	.C2V_19 (C2V_54_1205),
	.C2V_20 (C2V_54_1206),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU55 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_14_55),
	.V2C_2 (V2C_50_55),
	.V2C_3 (V2C_118_55),
	.V2C_4 (V2C_179_55),
	.V2C_5 (V2C_193_55),
	.V2C_6 (V2C_284_55),
	.V2C_7 (V2C_384_55),
	.V2C_8 (V2C_390_55),
	.V2C_9 (V2C_487_55),
	.V2C_10 (V2C_723_55),
	.V2C_11 (V2C_771_55),
	.V2C_12 (V2C_819_55),
	.V2C_13 (V2C_908_55),
	.V2C_14 (V2C_949_55),
	.V2C_15 (V2C_983_55),
	.V2C_16 (V2C_1022_55),
	.V2C_17 (V2C_1096_55),
	.V2C_18 (V2C_1107_55),
	.V2C_19 (V2C_1206_55),
	.V2C_20 (V2C_1207_55),
	.C2V_1 (C2V_55_14),
	.C2V_2 (C2V_55_50),
	.C2V_3 (C2V_55_118),
	.C2V_4 (C2V_55_179),
	.C2V_5 (C2V_55_193),
	.C2V_6 (C2V_55_284),
	.C2V_7 (C2V_55_384),
	.C2V_8 (C2V_55_390),
	.C2V_9 (C2V_55_487),
	.C2V_10 (C2V_55_723),
	.C2V_11 (C2V_55_771),
	.C2V_12 (C2V_55_819),
	.C2V_13 (C2V_55_908),
	.C2V_14 (C2V_55_949),
	.C2V_15 (C2V_55_983),
	.C2V_16 (C2V_55_1022),
	.C2V_17 (C2V_55_1096),
	.C2V_18 (C2V_55_1107),
	.C2V_19 (C2V_55_1206),
	.C2V_20 (C2V_55_1207),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU56 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_23_56),
	.V2C_2 (V2C_72_56),
	.V2C_3 (V2C_128_56),
	.V2C_4 (V2C_176_56),
	.V2C_5 (V2C_205_56),
	.V2C_6 (V2C_274_56),
	.V2C_7 (V2C_325_56),
	.V2C_8 (V2C_432_56),
	.V2C_9 (V2C_521_56),
	.V2C_10 (V2C_633_56),
	.V2C_11 (V2C_694_56),
	.V2C_12 (V2C_862_56),
	.V2C_13 (V2C_904_56),
	.V2C_14 (V2C_919_56),
	.V2C_15 (V2C_998_56),
	.V2C_16 (V2C_1030_56),
	.V2C_17 (V2C_1097_56),
	.V2C_18 (V2C_1128_56),
	.V2C_19 (V2C_1207_56),
	.V2C_20 (V2C_1208_56),
	.C2V_1 (C2V_56_23),
	.C2V_2 (C2V_56_72),
	.C2V_3 (C2V_56_128),
	.C2V_4 (C2V_56_176),
	.C2V_5 (C2V_56_205),
	.C2V_6 (C2V_56_274),
	.C2V_7 (C2V_56_325),
	.C2V_8 (C2V_56_432),
	.C2V_9 (C2V_56_521),
	.C2V_10 (C2V_56_633),
	.C2V_11 (C2V_56_694),
	.C2V_12 (C2V_56_862),
	.C2V_13 (C2V_56_904),
	.C2V_14 (C2V_56_919),
	.C2V_15 (C2V_56_998),
	.C2V_16 (C2V_56_1030),
	.C2V_17 (C2V_56_1097),
	.C2V_18 (C2V_56_1128),
	.C2V_19 (C2V_56_1207),
	.C2V_20 (C2V_56_1208),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU57 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_18_57),
	.V2C_2 (V2C_93_57),
	.V2C_3 (V2C_110_57),
	.V2C_4 (V2C_192_57),
	.V2C_5 (V2C_210_57),
	.V2C_6 (V2C_277_57),
	.V2C_7 (V2C_374_57),
	.V2C_8 (V2C_429_57),
	.V2C_9 (V2C_540_57),
	.V2C_10 (V2C_597_57),
	.V2C_11 (V2C_625_57),
	.V2C_12 (V2C_729_57),
	.V2C_13 (V2C_908_57),
	.V2C_14 (V2C_952_57),
	.V2C_15 (V2C_977_57),
	.V2C_16 (V2C_1037_57),
	.V2C_17 (V2C_1067_57),
	.V2C_18 (V2C_1112_57),
	.V2C_19 (V2C_1208_57),
	.V2C_20 (V2C_1209_57),
	.C2V_1 (C2V_57_18),
	.C2V_2 (C2V_57_93),
	.C2V_3 (C2V_57_110),
	.C2V_4 (C2V_57_192),
	.C2V_5 (C2V_57_210),
	.C2V_6 (C2V_57_277),
	.C2V_7 (C2V_57_374),
	.C2V_8 (C2V_57_429),
	.C2V_9 (C2V_57_540),
	.C2V_10 (C2V_57_597),
	.C2V_11 (C2V_57_625),
	.C2V_12 (C2V_57_729),
	.C2V_13 (C2V_57_908),
	.C2V_14 (C2V_57_952),
	.C2V_15 (C2V_57_977),
	.C2V_16 (C2V_57_1037),
	.C2V_17 (C2V_57_1067),
	.C2V_18 (C2V_57_1112),
	.C2V_19 (C2V_57_1208),
	.C2V_20 (C2V_57_1209),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU58 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_37_58),
	.V2C_2 (V2C_96_58),
	.V2C_3 (V2C_135_58),
	.V2C_4 (V2C_191_58),
	.V2C_5 (V2C_208_58),
	.V2C_6 (V2C_262_58),
	.V2C_7 (V2C_438_58),
	.V2C_8 (V2C_526_58),
	.V2C_9 (V2C_562_58),
	.V2C_10 (V2C_624_58),
	.V2C_11 (V2C_649_58),
	.V2C_12 (V2C_695_58),
	.V2C_13 (V2C_912_58),
	.V2C_14 (V2C_936_58),
	.V2C_15 (V2C_972_58),
	.V2C_16 (V2C_1050_58),
	.V2C_17 (V2C_1077_58),
	.V2C_18 (V2C_1141_58),
	.V2C_19 (V2C_1209_58),
	.V2C_20 (V2C_1210_58),
	.C2V_1 (C2V_58_37),
	.C2V_2 (C2V_58_96),
	.C2V_3 (C2V_58_135),
	.C2V_4 (C2V_58_191),
	.C2V_5 (C2V_58_208),
	.C2V_6 (C2V_58_262),
	.C2V_7 (C2V_58_438),
	.C2V_8 (C2V_58_526),
	.C2V_9 (C2V_58_562),
	.C2V_10 (C2V_58_624),
	.C2V_11 (C2V_58_649),
	.C2V_12 (C2V_58_695),
	.C2V_13 (C2V_58_912),
	.C2V_14 (C2V_58_936),
	.C2V_15 (C2V_58_972),
	.C2V_16 (C2V_58_1050),
	.C2V_17 (C2V_58_1077),
	.C2V_18 (C2V_58_1141),
	.C2V_19 (C2V_58_1209),
	.C2V_20 (C2V_58_1210),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU59 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_8_59),
	.V2C_2 (V2C_66_59),
	.V2C_3 (V2C_101_59),
	.V2C_4 (V2C_172_59),
	.V2C_5 (V2C_236_59),
	.V2C_6 (V2C_254_59),
	.V2C_7 (V2C_303_59),
	.V2C_8 (V2C_370_59),
	.V2C_9 (V2C_449_59),
	.V2C_10 (V2C_683_59),
	.V2C_11 (V2C_747_59),
	.V2C_12 (V2C_801_59),
	.V2C_13 (V2C_879_59),
	.V2C_14 (V2C_927_59),
	.V2C_15 (V2C_970_59),
	.V2C_16 (V2C_1022_59),
	.V2C_17 (V2C_1071_59),
	.V2C_18 (V2C_1119_59),
	.V2C_19 (V2C_1210_59),
	.V2C_20 (V2C_1211_59),
	.C2V_1 (C2V_59_8),
	.C2V_2 (C2V_59_66),
	.C2V_3 (C2V_59_101),
	.C2V_4 (C2V_59_172),
	.C2V_5 (C2V_59_236),
	.C2V_6 (C2V_59_254),
	.C2V_7 (C2V_59_303),
	.C2V_8 (C2V_59_370),
	.C2V_9 (C2V_59_449),
	.C2V_10 (C2V_59_683),
	.C2V_11 (C2V_59_747),
	.C2V_12 (C2V_59_801),
	.C2V_13 (C2V_59_879),
	.C2V_14 (C2V_59_927),
	.C2V_15 (C2V_59_970),
	.C2V_16 (C2V_59_1022),
	.C2V_17 (C2V_59_1071),
	.C2V_18 (C2V_59_1119),
	.C2V_19 (C2V_59_1210),
	.C2V_20 (C2V_59_1211),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU60 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_39_60),
	.V2C_2 (V2C_63_60),
	.V2C_3 (V2C_103_60),
	.V2C_4 (V2C_171_60),
	.V2C_5 (V2C_205_60),
	.V2C_6 (V2C_284_60),
	.V2C_7 (V2C_289_60),
	.V2C_8 (V2C_441_60),
	.V2C_9 (V2C_538_60),
	.V2C_10 (V2C_619_60),
	.V2C_11 (V2C_775_60),
	.V2C_12 (V2C_851_60),
	.V2C_13 (V2C_884_60),
	.V2C_14 (V2C_946_60),
	.V2C_15 (V2C_981_60),
	.V2C_16 (V2C_1048_60),
	.V2C_17 (V2C_1064_60),
	.V2C_18 (V2C_1114_60),
	.V2C_19 (V2C_1211_60),
	.V2C_20 (V2C_1212_60),
	.C2V_1 (C2V_60_39),
	.C2V_2 (C2V_60_63),
	.C2V_3 (C2V_60_103),
	.C2V_4 (C2V_60_171),
	.C2V_5 (C2V_60_205),
	.C2V_6 (C2V_60_284),
	.C2V_7 (C2V_60_289),
	.C2V_8 (C2V_60_441),
	.C2V_9 (C2V_60_538),
	.C2V_10 (C2V_60_619),
	.C2V_11 (C2V_60_775),
	.C2V_12 (C2V_60_851),
	.C2V_13 (C2V_60_884),
	.C2V_14 (C2V_60_946),
	.C2V_15 (C2V_60_981),
	.C2V_16 (C2V_60_1048),
	.C2V_17 (C2V_60_1064),
	.C2V_18 (C2V_60_1114),
	.C2V_19 (C2V_60_1211),
	.C2V_20 (C2V_60_1212),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU61 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_15_61),
	.V2C_2 (V2C_51_61),
	.V2C_3 (V2C_119_61),
	.V2C_4 (V2C_180_61),
	.V2C_5 (V2C_194_61),
	.V2C_6 (V2C_285_61),
	.V2C_7 (V2C_337_61),
	.V2C_8 (V2C_391_61),
	.V2C_9 (V2C_488_61),
	.V2C_10 (V2C_724_61),
	.V2C_11 (V2C_772_61),
	.V2C_12 (V2C_820_61),
	.V2C_13 (V2C_909_61),
	.V2C_14 (V2C_950_61),
	.V2C_15 (V2C_984_61),
	.V2C_16 (V2C_1023_61),
	.V2C_17 (V2C_1097_61),
	.V2C_18 (V2C_1108_61),
	.V2C_19 (V2C_1212_61),
	.V2C_20 (V2C_1213_61),
	.C2V_1 (C2V_61_15),
	.C2V_2 (C2V_61_51),
	.C2V_3 (C2V_61_119),
	.C2V_4 (C2V_61_180),
	.C2V_5 (C2V_61_194),
	.C2V_6 (C2V_61_285),
	.C2V_7 (C2V_61_337),
	.C2V_8 (C2V_61_391),
	.C2V_9 (C2V_61_488),
	.C2V_10 (C2V_61_724),
	.C2V_11 (C2V_61_772),
	.C2V_12 (C2V_61_820),
	.C2V_13 (C2V_61_909),
	.C2V_14 (C2V_61_950),
	.C2V_15 (C2V_61_984),
	.C2V_16 (C2V_61_1023),
	.C2V_17 (C2V_61_1097),
	.C2V_18 (C2V_61_1108),
	.C2V_19 (C2V_61_1212),
	.C2V_20 (C2V_61_1213),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU62 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_24_62),
	.V2C_2 (V2C_73_62),
	.V2C_3 (V2C_129_62),
	.V2C_4 (V2C_177_62),
	.V2C_5 (V2C_206_62),
	.V2C_6 (V2C_275_62),
	.V2C_7 (V2C_326_62),
	.V2C_8 (V2C_385_62),
	.V2C_9 (V2C_522_62),
	.V2C_10 (V2C_634_62),
	.V2C_11 (V2C_695_62),
	.V2C_12 (V2C_863_62),
	.V2C_13 (V2C_905_62),
	.V2C_14 (V2C_920_62),
	.V2C_15 (V2C_999_62),
	.V2C_16 (V2C_1031_62),
	.V2C_17 (V2C_1098_62),
	.V2C_18 (V2C_1129_62),
	.V2C_19 (V2C_1213_62),
	.V2C_20 (V2C_1214_62),
	.C2V_1 (C2V_62_24),
	.C2V_2 (C2V_62_73),
	.C2V_3 (C2V_62_129),
	.C2V_4 (C2V_62_177),
	.C2V_5 (C2V_62_206),
	.C2V_6 (C2V_62_275),
	.C2V_7 (C2V_62_326),
	.C2V_8 (C2V_62_385),
	.C2V_9 (C2V_62_522),
	.C2V_10 (C2V_62_634),
	.C2V_11 (C2V_62_695),
	.C2V_12 (C2V_62_863),
	.C2V_13 (C2V_62_905),
	.C2V_14 (C2V_62_920),
	.C2V_15 (C2V_62_999),
	.C2V_16 (C2V_62_1031),
	.C2V_17 (C2V_62_1098),
	.C2V_18 (C2V_62_1129),
	.C2V_19 (C2V_62_1213),
	.C2V_20 (C2V_62_1214),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU63 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_19_63),
	.V2C_2 (V2C_94_63),
	.V2C_3 (V2C_111_63),
	.V2C_4 (V2C_145_63),
	.V2C_5 (V2C_211_63),
	.V2C_6 (V2C_278_63),
	.V2C_7 (V2C_375_63),
	.V2C_8 (V2C_430_63),
	.V2C_9 (V2C_541_63),
	.V2C_10 (V2C_598_63),
	.V2C_11 (V2C_626_63),
	.V2C_12 (V2C_730_63),
	.V2C_13 (V2C_909_63),
	.V2C_14 (V2C_953_63),
	.V2C_15 (V2C_978_63),
	.V2C_16 (V2C_1038_63),
	.V2C_17 (V2C_1068_63),
	.V2C_18 (V2C_1113_63),
	.V2C_19 (V2C_1214_63),
	.V2C_20 (V2C_1215_63),
	.C2V_1 (C2V_63_19),
	.C2V_2 (C2V_63_94),
	.C2V_3 (C2V_63_111),
	.C2V_4 (C2V_63_145),
	.C2V_5 (C2V_63_211),
	.C2V_6 (C2V_63_278),
	.C2V_7 (C2V_63_375),
	.C2V_8 (C2V_63_430),
	.C2V_9 (C2V_63_541),
	.C2V_10 (C2V_63_598),
	.C2V_11 (C2V_63_626),
	.C2V_12 (C2V_63_730),
	.C2V_13 (C2V_63_909),
	.C2V_14 (C2V_63_953),
	.C2V_15 (C2V_63_978),
	.C2V_16 (C2V_63_1038),
	.C2V_17 (C2V_63_1068),
	.C2V_18 (C2V_63_1113),
	.C2V_19 (C2V_63_1214),
	.C2V_20 (C2V_63_1215),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU64 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_38_64),
	.V2C_2 (V2C_49_64),
	.V2C_3 (V2C_136_64),
	.V2C_4 (V2C_192_64),
	.V2C_5 (V2C_209_64),
	.V2C_6 (V2C_263_64),
	.V2C_7 (V2C_439_64),
	.V2C_8 (V2C_527_64),
	.V2C_9 (V2C_563_64),
	.V2C_10 (V2C_577_64),
	.V2C_11 (V2C_650_64),
	.V2C_12 (V2C_696_64),
	.V2C_13 (V2C_865_64),
	.V2C_14 (V2C_937_64),
	.V2C_15 (V2C_973_64),
	.V2C_16 (V2C_1051_64),
	.V2C_17 (V2C_1078_64),
	.V2C_18 (V2C_1142_64),
	.V2C_19 (V2C_1215_64),
	.V2C_20 (V2C_1216_64),
	.C2V_1 (C2V_64_38),
	.C2V_2 (C2V_64_49),
	.C2V_3 (C2V_64_136),
	.C2V_4 (C2V_64_192),
	.C2V_5 (C2V_64_209),
	.C2V_6 (C2V_64_263),
	.C2V_7 (C2V_64_439),
	.C2V_8 (C2V_64_527),
	.C2V_9 (C2V_64_563),
	.C2V_10 (C2V_64_577),
	.C2V_11 (C2V_64_650),
	.C2V_12 (C2V_64_696),
	.C2V_13 (C2V_64_865),
	.C2V_14 (C2V_64_937),
	.C2V_15 (C2V_64_973),
	.C2V_16 (C2V_64_1051),
	.C2V_17 (C2V_64_1078),
	.C2V_18 (C2V_64_1142),
	.C2V_19 (C2V_64_1215),
	.C2V_20 (C2V_64_1216),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU65 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_9_65),
	.V2C_2 (V2C_67_65),
	.V2C_3 (V2C_102_65),
	.V2C_4 (V2C_173_65),
	.V2C_5 (V2C_237_65),
	.V2C_6 (V2C_255_65),
	.V2C_7 (V2C_304_65),
	.V2C_8 (V2C_371_65),
	.V2C_9 (V2C_450_65),
	.V2C_10 (V2C_684_65),
	.V2C_11 (V2C_748_65),
	.V2C_12 (V2C_802_65),
	.V2C_13 (V2C_880_65),
	.V2C_14 (V2C_928_65),
	.V2C_15 (V2C_971_65),
	.V2C_16 (V2C_1023_65),
	.V2C_17 (V2C_1072_65),
	.V2C_18 (V2C_1120_65),
	.V2C_19 (V2C_1216_65),
	.V2C_20 (V2C_1217_65),
	.C2V_1 (C2V_65_9),
	.C2V_2 (C2V_65_67),
	.C2V_3 (C2V_65_102),
	.C2V_4 (C2V_65_173),
	.C2V_5 (C2V_65_237),
	.C2V_6 (C2V_65_255),
	.C2V_7 (C2V_65_304),
	.C2V_8 (C2V_65_371),
	.C2V_9 (C2V_65_450),
	.C2V_10 (C2V_65_684),
	.C2V_11 (C2V_65_748),
	.C2V_12 (C2V_65_802),
	.C2V_13 (C2V_65_880),
	.C2V_14 (C2V_65_928),
	.C2V_15 (C2V_65_971),
	.C2V_16 (C2V_65_1023),
	.C2V_17 (C2V_65_1072),
	.C2V_18 (C2V_65_1120),
	.C2V_19 (C2V_65_1216),
	.C2V_20 (C2V_65_1217),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU66 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_40_66),
	.V2C_2 (V2C_64_66),
	.V2C_3 (V2C_104_66),
	.V2C_4 (V2C_172_66),
	.V2C_5 (V2C_206_66),
	.V2C_6 (V2C_285_66),
	.V2C_7 (V2C_290_66),
	.V2C_8 (V2C_442_66),
	.V2C_9 (V2C_539_66),
	.V2C_10 (V2C_620_66),
	.V2C_11 (V2C_776_66),
	.V2C_12 (V2C_852_66),
	.V2C_13 (V2C_885_66),
	.V2C_14 (V2C_947_66),
	.V2C_15 (V2C_982_66),
	.V2C_16 (V2C_1049_66),
	.V2C_17 (V2C_1065_66),
	.V2C_18 (V2C_1115_66),
	.V2C_19 (V2C_1217_66),
	.V2C_20 (V2C_1218_66),
	.C2V_1 (C2V_66_40),
	.C2V_2 (C2V_66_64),
	.C2V_3 (C2V_66_104),
	.C2V_4 (C2V_66_172),
	.C2V_5 (C2V_66_206),
	.C2V_6 (C2V_66_285),
	.C2V_7 (C2V_66_290),
	.C2V_8 (C2V_66_442),
	.C2V_9 (C2V_66_539),
	.C2V_10 (C2V_66_620),
	.C2V_11 (C2V_66_776),
	.C2V_12 (C2V_66_852),
	.C2V_13 (C2V_66_885),
	.C2V_14 (C2V_66_947),
	.C2V_15 (C2V_66_982),
	.C2V_16 (C2V_66_1049),
	.C2V_17 (C2V_66_1065),
	.C2V_18 (C2V_66_1115),
	.C2V_19 (C2V_66_1217),
	.C2V_20 (C2V_66_1218),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU67 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_16_67),
	.V2C_2 (V2C_52_67),
	.V2C_3 (V2C_120_67),
	.V2C_4 (V2C_181_67),
	.V2C_5 (V2C_195_67),
	.V2C_6 (V2C_286_67),
	.V2C_7 (V2C_338_67),
	.V2C_8 (V2C_392_67),
	.V2C_9 (V2C_489_67),
	.V2C_10 (V2C_725_67),
	.V2C_11 (V2C_773_67),
	.V2C_12 (V2C_821_67),
	.V2C_13 (V2C_910_67),
	.V2C_14 (V2C_951_67),
	.V2C_15 (V2C_985_67),
	.V2C_16 (V2C_1024_67),
	.V2C_17 (V2C_1098_67),
	.V2C_18 (V2C_1109_67),
	.V2C_19 (V2C_1218_67),
	.V2C_20 (V2C_1219_67),
	.C2V_1 (C2V_67_16),
	.C2V_2 (C2V_67_52),
	.C2V_3 (C2V_67_120),
	.C2V_4 (C2V_67_181),
	.C2V_5 (C2V_67_195),
	.C2V_6 (C2V_67_286),
	.C2V_7 (C2V_67_338),
	.C2V_8 (C2V_67_392),
	.C2V_9 (C2V_67_489),
	.C2V_10 (C2V_67_725),
	.C2V_11 (C2V_67_773),
	.C2V_12 (C2V_67_821),
	.C2V_13 (C2V_67_910),
	.C2V_14 (C2V_67_951),
	.C2V_15 (C2V_67_985),
	.C2V_16 (C2V_67_1024),
	.C2V_17 (C2V_67_1098),
	.C2V_18 (C2V_67_1109),
	.C2V_19 (C2V_67_1218),
	.C2V_20 (C2V_67_1219),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU68 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_25_68),
	.V2C_2 (V2C_74_68),
	.V2C_3 (V2C_130_68),
	.V2C_4 (V2C_178_68),
	.V2C_5 (V2C_207_68),
	.V2C_6 (V2C_276_68),
	.V2C_7 (V2C_327_68),
	.V2C_8 (V2C_386_68),
	.V2C_9 (V2C_523_68),
	.V2C_10 (V2C_635_68),
	.V2C_11 (V2C_696_68),
	.V2C_12 (V2C_864_68),
	.V2C_13 (V2C_906_68),
	.V2C_14 (V2C_921_68),
	.V2C_15 (V2C_1000_68),
	.V2C_16 (V2C_1032_68),
	.V2C_17 (V2C_1099_68),
	.V2C_18 (V2C_1130_68),
	.V2C_19 (V2C_1219_68),
	.V2C_20 (V2C_1220_68),
	.C2V_1 (C2V_68_25),
	.C2V_2 (C2V_68_74),
	.C2V_3 (C2V_68_130),
	.C2V_4 (C2V_68_178),
	.C2V_5 (C2V_68_207),
	.C2V_6 (C2V_68_276),
	.C2V_7 (C2V_68_327),
	.C2V_8 (C2V_68_386),
	.C2V_9 (C2V_68_523),
	.C2V_10 (C2V_68_635),
	.C2V_11 (C2V_68_696),
	.C2V_12 (C2V_68_864),
	.C2V_13 (C2V_68_906),
	.C2V_14 (C2V_68_921),
	.C2V_15 (C2V_68_1000),
	.C2V_16 (C2V_68_1032),
	.C2V_17 (C2V_68_1099),
	.C2V_18 (C2V_68_1130),
	.C2V_19 (C2V_68_1219),
	.C2V_20 (C2V_68_1220),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU69 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_20_69),
	.V2C_2 (V2C_95_69),
	.V2C_3 (V2C_112_69),
	.V2C_4 (V2C_146_69),
	.V2C_5 (V2C_212_69),
	.V2C_6 (V2C_279_69),
	.V2C_7 (V2C_376_69),
	.V2C_8 (V2C_431_69),
	.V2C_9 (V2C_542_69),
	.V2C_10 (V2C_599_69),
	.V2C_11 (V2C_627_69),
	.V2C_12 (V2C_731_69),
	.V2C_13 (V2C_910_69),
	.V2C_14 (V2C_954_69),
	.V2C_15 (V2C_979_69),
	.V2C_16 (V2C_1039_69),
	.V2C_17 (V2C_1069_69),
	.V2C_18 (V2C_1114_69),
	.V2C_19 (V2C_1220_69),
	.V2C_20 (V2C_1221_69),
	.C2V_1 (C2V_69_20),
	.C2V_2 (C2V_69_95),
	.C2V_3 (C2V_69_112),
	.C2V_4 (C2V_69_146),
	.C2V_5 (C2V_69_212),
	.C2V_6 (C2V_69_279),
	.C2V_7 (C2V_69_376),
	.C2V_8 (C2V_69_431),
	.C2V_9 (C2V_69_542),
	.C2V_10 (C2V_69_599),
	.C2V_11 (C2V_69_627),
	.C2V_12 (C2V_69_731),
	.C2V_13 (C2V_69_910),
	.C2V_14 (C2V_69_954),
	.C2V_15 (C2V_69_979),
	.C2V_16 (C2V_69_1039),
	.C2V_17 (C2V_69_1069),
	.C2V_18 (C2V_69_1114),
	.C2V_19 (C2V_69_1220),
	.C2V_20 (C2V_69_1221),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU70 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_39_70),
	.V2C_2 (V2C_50_70),
	.V2C_3 (V2C_137_70),
	.V2C_4 (V2C_145_70),
	.V2C_5 (V2C_210_70),
	.V2C_6 (V2C_264_70),
	.V2C_7 (V2C_440_70),
	.V2C_8 (V2C_528_70),
	.V2C_9 (V2C_564_70),
	.V2C_10 (V2C_578_70),
	.V2C_11 (V2C_651_70),
	.V2C_12 (V2C_697_70),
	.V2C_13 (V2C_866_70),
	.V2C_14 (V2C_938_70),
	.V2C_15 (V2C_974_70),
	.V2C_16 (V2C_1052_70),
	.V2C_17 (V2C_1079_70),
	.V2C_18 (V2C_1143_70),
	.V2C_19 (V2C_1221_70),
	.V2C_20 (V2C_1222_70),
	.C2V_1 (C2V_70_39),
	.C2V_2 (C2V_70_50),
	.C2V_3 (C2V_70_137),
	.C2V_4 (C2V_70_145),
	.C2V_5 (C2V_70_210),
	.C2V_6 (C2V_70_264),
	.C2V_7 (C2V_70_440),
	.C2V_8 (C2V_70_528),
	.C2V_9 (C2V_70_564),
	.C2V_10 (C2V_70_578),
	.C2V_11 (C2V_70_651),
	.C2V_12 (C2V_70_697),
	.C2V_13 (C2V_70_866),
	.C2V_14 (C2V_70_938),
	.C2V_15 (C2V_70_974),
	.C2V_16 (C2V_70_1052),
	.C2V_17 (C2V_70_1079),
	.C2V_18 (C2V_70_1143),
	.C2V_19 (C2V_70_1221),
	.C2V_20 (C2V_70_1222),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU71 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_10_71),
	.V2C_2 (V2C_68_71),
	.V2C_3 (V2C_103_71),
	.V2C_4 (V2C_174_71),
	.V2C_5 (V2C_238_71),
	.V2C_6 (V2C_256_71),
	.V2C_7 (V2C_305_71),
	.V2C_8 (V2C_372_71),
	.V2C_9 (V2C_451_71),
	.V2C_10 (V2C_685_71),
	.V2C_11 (V2C_749_71),
	.V2C_12 (V2C_803_71),
	.V2C_13 (V2C_881_71),
	.V2C_14 (V2C_929_71),
	.V2C_15 (V2C_972_71),
	.V2C_16 (V2C_1024_71),
	.V2C_17 (V2C_1073_71),
	.V2C_18 (V2C_1121_71),
	.V2C_19 (V2C_1222_71),
	.V2C_20 (V2C_1223_71),
	.C2V_1 (C2V_71_10),
	.C2V_2 (C2V_71_68),
	.C2V_3 (C2V_71_103),
	.C2V_4 (C2V_71_174),
	.C2V_5 (C2V_71_238),
	.C2V_6 (C2V_71_256),
	.C2V_7 (C2V_71_305),
	.C2V_8 (C2V_71_372),
	.C2V_9 (C2V_71_451),
	.C2V_10 (C2V_71_685),
	.C2V_11 (C2V_71_749),
	.C2V_12 (C2V_71_803),
	.C2V_13 (C2V_71_881),
	.C2V_14 (C2V_71_929),
	.C2V_15 (C2V_71_972),
	.C2V_16 (C2V_71_1024),
	.C2V_17 (C2V_71_1073),
	.C2V_18 (C2V_71_1121),
	.C2V_19 (C2V_71_1222),
	.C2V_20 (C2V_71_1223),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU72 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_41_72),
	.V2C_2 (V2C_65_72),
	.V2C_3 (V2C_105_72),
	.V2C_4 (V2C_173_72),
	.V2C_5 (V2C_207_72),
	.V2C_6 (V2C_286_72),
	.V2C_7 (V2C_291_72),
	.V2C_8 (V2C_443_72),
	.V2C_9 (V2C_540_72),
	.V2C_10 (V2C_621_72),
	.V2C_11 (V2C_777_72),
	.V2C_12 (V2C_853_72),
	.V2C_13 (V2C_886_72),
	.V2C_14 (V2C_948_72),
	.V2C_15 (V2C_983_72),
	.V2C_16 (V2C_1050_72),
	.V2C_17 (V2C_1066_72),
	.V2C_18 (V2C_1116_72),
	.V2C_19 (V2C_1223_72),
	.V2C_20 (V2C_1224_72),
	.C2V_1 (C2V_72_41),
	.C2V_2 (C2V_72_65),
	.C2V_3 (C2V_72_105),
	.C2V_4 (C2V_72_173),
	.C2V_5 (C2V_72_207),
	.C2V_6 (C2V_72_286),
	.C2V_7 (C2V_72_291),
	.C2V_8 (C2V_72_443),
	.C2V_9 (C2V_72_540),
	.C2V_10 (C2V_72_621),
	.C2V_11 (C2V_72_777),
	.C2V_12 (C2V_72_853),
	.C2V_13 (C2V_72_886),
	.C2V_14 (C2V_72_948),
	.C2V_15 (C2V_72_983),
	.C2V_16 (C2V_72_1050),
	.C2V_17 (C2V_72_1066),
	.C2V_18 (C2V_72_1116),
	.C2V_19 (C2V_72_1223),
	.C2V_20 (C2V_72_1224),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU73 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_17_73),
	.V2C_2 (V2C_53_73),
	.V2C_3 (V2C_121_73),
	.V2C_4 (V2C_182_73),
	.V2C_5 (V2C_196_73),
	.V2C_6 (V2C_287_73),
	.V2C_7 (V2C_339_73),
	.V2C_8 (V2C_393_73),
	.V2C_9 (V2C_490_73),
	.V2C_10 (V2C_726_73),
	.V2C_11 (V2C_774_73),
	.V2C_12 (V2C_822_73),
	.V2C_13 (V2C_911_73),
	.V2C_14 (V2C_952_73),
	.V2C_15 (V2C_986_73),
	.V2C_16 (V2C_1025_73),
	.V2C_17 (V2C_1099_73),
	.V2C_18 (V2C_1110_73),
	.V2C_19 (V2C_1224_73),
	.V2C_20 (V2C_1225_73),
	.C2V_1 (C2V_73_17),
	.C2V_2 (C2V_73_53),
	.C2V_3 (C2V_73_121),
	.C2V_4 (C2V_73_182),
	.C2V_5 (C2V_73_196),
	.C2V_6 (C2V_73_287),
	.C2V_7 (C2V_73_339),
	.C2V_8 (C2V_73_393),
	.C2V_9 (C2V_73_490),
	.C2V_10 (C2V_73_726),
	.C2V_11 (C2V_73_774),
	.C2V_12 (C2V_73_822),
	.C2V_13 (C2V_73_911),
	.C2V_14 (C2V_73_952),
	.C2V_15 (C2V_73_986),
	.C2V_16 (C2V_73_1025),
	.C2V_17 (C2V_73_1099),
	.C2V_18 (C2V_73_1110),
	.C2V_19 (C2V_73_1224),
	.C2V_20 (C2V_73_1225),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU74 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_26_74),
	.V2C_2 (V2C_75_74),
	.V2C_3 (V2C_131_74),
	.V2C_4 (V2C_179_74),
	.V2C_5 (V2C_208_74),
	.V2C_6 (V2C_277_74),
	.V2C_7 (V2C_328_74),
	.V2C_8 (V2C_387_74),
	.V2C_9 (V2C_524_74),
	.V2C_10 (V2C_636_74),
	.V2C_11 (V2C_697_74),
	.V2C_12 (V2C_817_74),
	.V2C_13 (V2C_907_74),
	.V2C_14 (V2C_922_74),
	.V2C_15 (V2C_1001_74),
	.V2C_16 (V2C_1033_74),
	.V2C_17 (V2C_1100_74),
	.V2C_18 (V2C_1131_74),
	.V2C_19 (V2C_1225_74),
	.V2C_20 (V2C_1226_74),
	.C2V_1 (C2V_74_26),
	.C2V_2 (C2V_74_75),
	.C2V_3 (C2V_74_131),
	.C2V_4 (C2V_74_179),
	.C2V_5 (C2V_74_208),
	.C2V_6 (C2V_74_277),
	.C2V_7 (C2V_74_328),
	.C2V_8 (C2V_74_387),
	.C2V_9 (C2V_74_524),
	.C2V_10 (C2V_74_636),
	.C2V_11 (C2V_74_697),
	.C2V_12 (C2V_74_817),
	.C2V_13 (C2V_74_907),
	.C2V_14 (C2V_74_922),
	.C2V_15 (C2V_74_1001),
	.C2V_16 (C2V_74_1033),
	.C2V_17 (C2V_74_1100),
	.C2V_18 (C2V_74_1131),
	.C2V_19 (C2V_74_1225),
	.C2V_20 (C2V_74_1226),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU75 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_21_75),
	.V2C_2 (V2C_96_75),
	.V2C_3 (V2C_113_75),
	.V2C_4 (V2C_147_75),
	.V2C_5 (V2C_213_75),
	.V2C_6 (V2C_280_75),
	.V2C_7 (V2C_377_75),
	.V2C_8 (V2C_432_75),
	.V2C_9 (V2C_543_75),
	.V2C_10 (V2C_600_75),
	.V2C_11 (V2C_628_75),
	.V2C_12 (V2C_732_75),
	.V2C_13 (V2C_911_75),
	.V2C_14 (V2C_955_75),
	.V2C_15 (V2C_980_75),
	.V2C_16 (V2C_1040_75),
	.V2C_17 (V2C_1070_75),
	.V2C_18 (V2C_1115_75),
	.V2C_19 (V2C_1226_75),
	.V2C_20 (V2C_1227_75),
	.C2V_1 (C2V_75_21),
	.C2V_2 (C2V_75_96),
	.C2V_3 (C2V_75_113),
	.C2V_4 (C2V_75_147),
	.C2V_5 (C2V_75_213),
	.C2V_6 (C2V_75_280),
	.C2V_7 (C2V_75_377),
	.C2V_8 (C2V_75_432),
	.C2V_9 (C2V_75_543),
	.C2V_10 (C2V_75_600),
	.C2V_11 (C2V_75_628),
	.C2V_12 (C2V_75_732),
	.C2V_13 (C2V_75_911),
	.C2V_14 (C2V_75_955),
	.C2V_15 (C2V_75_980),
	.C2V_16 (C2V_75_1040),
	.C2V_17 (C2V_75_1070),
	.C2V_18 (C2V_75_1115),
	.C2V_19 (C2V_75_1226),
	.C2V_20 (C2V_75_1227),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU76 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_40_76),
	.V2C_2 (V2C_51_76),
	.V2C_3 (V2C_138_76),
	.V2C_4 (V2C_146_76),
	.V2C_5 (V2C_211_76),
	.V2C_6 (V2C_265_76),
	.V2C_7 (V2C_441_76),
	.V2C_8 (V2C_481_76),
	.V2C_9 (V2C_565_76),
	.V2C_10 (V2C_579_76),
	.V2C_11 (V2C_652_76),
	.V2C_12 (V2C_698_76),
	.V2C_13 (V2C_867_76),
	.V2C_14 (V2C_939_76),
	.V2C_15 (V2C_975_76),
	.V2C_16 (V2C_1053_76),
	.V2C_17 (V2C_1080_76),
	.V2C_18 (V2C_1144_76),
	.V2C_19 (V2C_1227_76),
	.V2C_20 (V2C_1228_76),
	.C2V_1 (C2V_76_40),
	.C2V_2 (C2V_76_51),
	.C2V_3 (C2V_76_138),
	.C2V_4 (C2V_76_146),
	.C2V_5 (C2V_76_211),
	.C2V_6 (C2V_76_265),
	.C2V_7 (C2V_76_441),
	.C2V_8 (C2V_76_481),
	.C2V_9 (C2V_76_565),
	.C2V_10 (C2V_76_579),
	.C2V_11 (C2V_76_652),
	.C2V_12 (C2V_76_698),
	.C2V_13 (C2V_76_867),
	.C2V_14 (C2V_76_939),
	.C2V_15 (C2V_76_975),
	.C2V_16 (C2V_76_1053),
	.C2V_17 (C2V_76_1080),
	.C2V_18 (C2V_76_1144),
	.C2V_19 (C2V_76_1227),
	.C2V_20 (C2V_76_1228),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU77 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_11_77),
	.V2C_2 (V2C_69_77),
	.V2C_3 (V2C_104_77),
	.V2C_4 (V2C_175_77),
	.V2C_5 (V2C_239_77),
	.V2C_6 (V2C_257_77),
	.V2C_7 (V2C_306_77),
	.V2C_8 (V2C_373_77),
	.V2C_9 (V2C_452_77),
	.V2C_10 (V2C_686_77),
	.V2C_11 (V2C_750_77),
	.V2C_12 (V2C_804_77),
	.V2C_13 (V2C_882_77),
	.V2C_14 (V2C_930_77),
	.V2C_15 (V2C_973_77),
	.V2C_16 (V2C_1025_77),
	.V2C_17 (V2C_1074_77),
	.V2C_18 (V2C_1122_77),
	.V2C_19 (V2C_1228_77),
	.V2C_20 (V2C_1229_77),
	.C2V_1 (C2V_77_11),
	.C2V_2 (C2V_77_69),
	.C2V_3 (C2V_77_104),
	.C2V_4 (C2V_77_175),
	.C2V_5 (C2V_77_239),
	.C2V_6 (C2V_77_257),
	.C2V_7 (C2V_77_306),
	.C2V_8 (C2V_77_373),
	.C2V_9 (C2V_77_452),
	.C2V_10 (C2V_77_686),
	.C2V_11 (C2V_77_750),
	.C2V_12 (C2V_77_804),
	.C2V_13 (C2V_77_882),
	.C2V_14 (C2V_77_930),
	.C2V_15 (C2V_77_973),
	.C2V_16 (C2V_77_1025),
	.C2V_17 (C2V_77_1074),
	.C2V_18 (C2V_77_1122),
	.C2V_19 (C2V_77_1228),
	.C2V_20 (C2V_77_1229),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU78 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_42_78),
	.V2C_2 (V2C_66_78),
	.V2C_3 (V2C_106_78),
	.V2C_4 (V2C_174_78),
	.V2C_5 (V2C_208_78),
	.V2C_6 (V2C_287_78),
	.V2C_7 (V2C_292_78),
	.V2C_8 (V2C_444_78),
	.V2C_9 (V2C_541_78),
	.V2C_10 (V2C_622_78),
	.V2C_11 (V2C_778_78),
	.V2C_12 (V2C_854_78),
	.V2C_13 (V2C_887_78),
	.V2C_14 (V2C_949_78),
	.V2C_15 (V2C_984_78),
	.V2C_16 (V2C_1051_78),
	.V2C_17 (V2C_1067_78),
	.V2C_18 (V2C_1117_78),
	.V2C_19 (V2C_1229_78),
	.V2C_20 (V2C_1230_78),
	.C2V_1 (C2V_78_42),
	.C2V_2 (C2V_78_66),
	.C2V_3 (C2V_78_106),
	.C2V_4 (C2V_78_174),
	.C2V_5 (C2V_78_208),
	.C2V_6 (C2V_78_287),
	.C2V_7 (C2V_78_292),
	.C2V_8 (C2V_78_444),
	.C2V_9 (C2V_78_541),
	.C2V_10 (C2V_78_622),
	.C2V_11 (C2V_78_778),
	.C2V_12 (C2V_78_854),
	.C2V_13 (C2V_78_887),
	.C2V_14 (C2V_78_949),
	.C2V_15 (C2V_78_984),
	.C2V_16 (C2V_78_1051),
	.C2V_17 (C2V_78_1067),
	.C2V_18 (C2V_78_1117),
	.C2V_19 (C2V_78_1229),
	.C2V_20 (C2V_78_1230),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU79 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_18_79),
	.V2C_2 (V2C_54_79),
	.V2C_3 (V2C_122_79),
	.V2C_4 (V2C_183_79),
	.V2C_5 (V2C_197_79),
	.V2C_6 (V2C_288_79),
	.V2C_7 (V2C_340_79),
	.V2C_8 (V2C_394_79),
	.V2C_9 (V2C_491_79),
	.V2C_10 (V2C_727_79),
	.V2C_11 (V2C_775_79),
	.V2C_12 (V2C_823_79),
	.V2C_13 (V2C_912_79),
	.V2C_14 (V2C_953_79),
	.V2C_15 (V2C_987_79),
	.V2C_16 (V2C_1026_79),
	.V2C_17 (V2C_1100_79),
	.V2C_18 (V2C_1111_79),
	.V2C_19 (V2C_1230_79),
	.V2C_20 (V2C_1231_79),
	.C2V_1 (C2V_79_18),
	.C2V_2 (C2V_79_54),
	.C2V_3 (C2V_79_122),
	.C2V_4 (C2V_79_183),
	.C2V_5 (C2V_79_197),
	.C2V_6 (C2V_79_288),
	.C2V_7 (C2V_79_340),
	.C2V_8 (C2V_79_394),
	.C2V_9 (C2V_79_491),
	.C2V_10 (C2V_79_727),
	.C2V_11 (C2V_79_775),
	.C2V_12 (C2V_79_823),
	.C2V_13 (C2V_79_912),
	.C2V_14 (C2V_79_953),
	.C2V_15 (C2V_79_987),
	.C2V_16 (C2V_79_1026),
	.C2V_17 (C2V_79_1100),
	.C2V_18 (C2V_79_1111),
	.C2V_19 (C2V_79_1230),
	.C2V_20 (C2V_79_1231),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU80 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_27_80),
	.V2C_2 (V2C_76_80),
	.V2C_3 (V2C_132_80),
	.V2C_4 (V2C_180_80),
	.V2C_5 (V2C_209_80),
	.V2C_6 (V2C_278_80),
	.V2C_7 (V2C_329_80),
	.V2C_8 (V2C_388_80),
	.V2C_9 (V2C_525_80),
	.V2C_10 (V2C_637_80),
	.V2C_11 (V2C_698_80),
	.V2C_12 (V2C_818_80),
	.V2C_13 (V2C_908_80),
	.V2C_14 (V2C_923_80),
	.V2C_15 (V2C_1002_80),
	.V2C_16 (V2C_1034_80),
	.V2C_17 (V2C_1101_80),
	.V2C_18 (V2C_1132_80),
	.V2C_19 (V2C_1231_80),
	.V2C_20 (V2C_1232_80),
	.C2V_1 (C2V_80_27),
	.C2V_2 (C2V_80_76),
	.C2V_3 (C2V_80_132),
	.C2V_4 (C2V_80_180),
	.C2V_5 (C2V_80_209),
	.C2V_6 (C2V_80_278),
	.C2V_7 (C2V_80_329),
	.C2V_8 (C2V_80_388),
	.C2V_9 (C2V_80_525),
	.C2V_10 (C2V_80_637),
	.C2V_11 (C2V_80_698),
	.C2V_12 (C2V_80_818),
	.C2V_13 (C2V_80_908),
	.C2V_14 (C2V_80_923),
	.C2V_15 (C2V_80_1002),
	.C2V_16 (C2V_80_1034),
	.C2V_17 (C2V_80_1101),
	.C2V_18 (C2V_80_1132),
	.C2V_19 (C2V_80_1231),
	.C2V_20 (C2V_80_1232),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU81 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_22_81),
	.V2C_2 (V2C_49_81),
	.V2C_3 (V2C_114_81),
	.V2C_4 (V2C_148_81),
	.V2C_5 (V2C_214_81),
	.V2C_6 (V2C_281_81),
	.V2C_7 (V2C_378_81),
	.V2C_8 (V2C_385_81),
	.V2C_9 (V2C_544_81),
	.V2C_10 (V2C_601_81),
	.V2C_11 (V2C_629_81),
	.V2C_12 (V2C_733_81),
	.V2C_13 (V2C_912_81),
	.V2C_14 (V2C_956_81),
	.V2C_15 (V2C_981_81),
	.V2C_16 (V2C_1041_81),
	.V2C_17 (V2C_1071_81),
	.V2C_18 (V2C_1116_81),
	.V2C_19 (V2C_1232_81),
	.V2C_20 (V2C_1233_81),
	.C2V_1 (C2V_81_22),
	.C2V_2 (C2V_81_49),
	.C2V_3 (C2V_81_114),
	.C2V_4 (C2V_81_148),
	.C2V_5 (C2V_81_214),
	.C2V_6 (C2V_81_281),
	.C2V_7 (C2V_81_378),
	.C2V_8 (C2V_81_385),
	.C2V_9 (C2V_81_544),
	.C2V_10 (C2V_81_601),
	.C2V_11 (C2V_81_629),
	.C2V_12 (C2V_81_733),
	.C2V_13 (C2V_81_912),
	.C2V_14 (C2V_81_956),
	.C2V_15 (C2V_81_981),
	.C2V_16 (C2V_81_1041),
	.C2V_17 (C2V_81_1071),
	.C2V_18 (C2V_81_1116),
	.C2V_19 (C2V_81_1232),
	.C2V_20 (C2V_81_1233),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU82 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_41_82),
	.V2C_2 (V2C_52_82),
	.V2C_3 (V2C_139_82),
	.V2C_4 (V2C_147_82),
	.V2C_5 (V2C_212_82),
	.V2C_6 (V2C_266_82),
	.V2C_7 (V2C_442_82),
	.V2C_8 (V2C_482_82),
	.V2C_9 (V2C_566_82),
	.V2C_10 (V2C_580_82),
	.V2C_11 (V2C_653_82),
	.V2C_12 (V2C_699_82),
	.V2C_13 (V2C_868_82),
	.V2C_14 (V2C_940_82),
	.V2C_15 (V2C_976_82),
	.V2C_16 (V2C_1054_82),
	.V2C_17 (V2C_1081_82),
	.V2C_18 (V2C_1145_82),
	.V2C_19 (V2C_1233_82),
	.V2C_20 (V2C_1234_82),
	.C2V_1 (C2V_82_41),
	.C2V_2 (C2V_82_52),
	.C2V_3 (C2V_82_139),
	.C2V_4 (C2V_82_147),
	.C2V_5 (C2V_82_212),
	.C2V_6 (C2V_82_266),
	.C2V_7 (C2V_82_442),
	.C2V_8 (C2V_82_482),
	.C2V_9 (C2V_82_566),
	.C2V_10 (C2V_82_580),
	.C2V_11 (C2V_82_653),
	.C2V_12 (C2V_82_699),
	.C2V_13 (C2V_82_868),
	.C2V_14 (C2V_82_940),
	.C2V_15 (C2V_82_976),
	.C2V_16 (C2V_82_1054),
	.C2V_17 (C2V_82_1081),
	.C2V_18 (C2V_82_1145),
	.C2V_19 (C2V_82_1233),
	.C2V_20 (C2V_82_1234),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU83 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_12_83),
	.V2C_2 (V2C_70_83),
	.V2C_3 (V2C_105_83),
	.V2C_4 (V2C_176_83),
	.V2C_5 (V2C_240_83),
	.V2C_6 (V2C_258_83),
	.V2C_7 (V2C_307_83),
	.V2C_8 (V2C_374_83),
	.V2C_9 (V2C_453_83),
	.V2C_10 (V2C_687_83),
	.V2C_11 (V2C_751_83),
	.V2C_12 (V2C_805_83),
	.V2C_13 (V2C_883_83),
	.V2C_14 (V2C_931_83),
	.V2C_15 (V2C_974_83),
	.V2C_16 (V2C_1026_83),
	.V2C_17 (V2C_1075_83),
	.V2C_18 (V2C_1123_83),
	.V2C_19 (V2C_1234_83),
	.V2C_20 (V2C_1235_83),
	.C2V_1 (C2V_83_12),
	.C2V_2 (C2V_83_70),
	.C2V_3 (C2V_83_105),
	.C2V_4 (C2V_83_176),
	.C2V_5 (C2V_83_240),
	.C2V_6 (C2V_83_258),
	.C2V_7 (C2V_83_307),
	.C2V_8 (C2V_83_374),
	.C2V_9 (C2V_83_453),
	.C2V_10 (C2V_83_687),
	.C2V_11 (C2V_83_751),
	.C2V_12 (C2V_83_805),
	.C2V_13 (C2V_83_883),
	.C2V_14 (C2V_83_931),
	.C2V_15 (C2V_83_974),
	.C2V_16 (C2V_83_1026),
	.C2V_17 (C2V_83_1075),
	.C2V_18 (C2V_83_1123),
	.C2V_19 (C2V_83_1234),
	.C2V_20 (C2V_83_1235),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU84 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_43_84),
	.V2C_2 (V2C_67_84),
	.V2C_3 (V2C_107_84),
	.V2C_4 (V2C_175_84),
	.V2C_5 (V2C_209_84),
	.V2C_6 (V2C_288_84),
	.V2C_7 (V2C_293_84),
	.V2C_8 (V2C_445_84),
	.V2C_9 (V2C_542_84),
	.V2C_10 (V2C_623_84),
	.V2C_11 (V2C_779_84),
	.V2C_12 (V2C_855_84),
	.V2C_13 (V2C_888_84),
	.V2C_14 (V2C_950_84),
	.V2C_15 (V2C_985_84),
	.V2C_16 (V2C_1052_84),
	.V2C_17 (V2C_1068_84),
	.V2C_18 (V2C_1118_84),
	.V2C_19 (V2C_1235_84),
	.V2C_20 (V2C_1236_84),
	.C2V_1 (C2V_84_43),
	.C2V_2 (C2V_84_67),
	.C2V_3 (C2V_84_107),
	.C2V_4 (C2V_84_175),
	.C2V_5 (C2V_84_209),
	.C2V_6 (C2V_84_288),
	.C2V_7 (C2V_84_293),
	.C2V_8 (C2V_84_445),
	.C2V_9 (C2V_84_542),
	.C2V_10 (C2V_84_623),
	.C2V_11 (C2V_84_779),
	.C2V_12 (C2V_84_855),
	.C2V_13 (C2V_84_888),
	.C2V_14 (C2V_84_950),
	.C2V_15 (C2V_84_985),
	.C2V_16 (C2V_84_1052),
	.C2V_17 (C2V_84_1068),
	.C2V_18 (C2V_84_1118),
	.C2V_19 (C2V_84_1235),
	.C2V_20 (C2V_84_1236),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU85 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_19_85),
	.V2C_2 (V2C_55_85),
	.V2C_3 (V2C_123_85),
	.V2C_4 (V2C_184_85),
	.V2C_5 (V2C_198_85),
	.V2C_6 (V2C_241_85),
	.V2C_7 (V2C_341_85),
	.V2C_8 (V2C_395_85),
	.V2C_9 (V2C_492_85),
	.V2C_10 (V2C_728_85),
	.V2C_11 (V2C_776_85),
	.V2C_12 (V2C_824_85),
	.V2C_13 (V2C_865_85),
	.V2C_14 (V2C_954_85),
	.V2C_15 (V2C_988_85),
	.V2C_16 (V2C_1027_85),
	.V2C_17 (V2C_1101_85),
	.V2C_18 (V2C_1112_85),
	.V2C_19 (V2C_1236_85),
	.V2C_20 (V2C_1237_85),
	.C2V_1 (C2V_85_19),
	.C2V_2 (C2V_85_55),
	.C2V_3 (C2V_85_123),
	.C2V_4 (C2V_85_184),
	.C2V_5 (C2V_85_198),
	.C2V_6 (C2V_85_241),
	.C2V_7 (C2V_85_341),
	.C2V_8 (C2V_85_395),
	.C2V_9 (C2V_85_492),
	.C2V_10 (C2V_85_728),
	.C2V_11 (C2V_85_776),
	.C2V_12 (C2V_85_824),
	.C2V_13 (C2V_85_865),
	.C2V_14 (C2V_85_954),
	.C2V_15 (C2V_85_988),
	.C2V_16 (C2V_85_1027),
	.C2V_17 (C2V_85_1101),
	.C2V_18 (C2V_85_1112),
	.C2V_19 (C2V_85_1236),
	.C2V_20 (C2V_85_1237),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU86 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_28_86),
	.V2C_2 (V2C_77_86),
	.V2C_3 (V2C_133_86),
	.V2C_4 (V2C_181_86),
	.V2C_5 (V2C_210_86),
	.V2C_6 (V2C_279_86),
	.V2C_7 (V2C_330_86),
	.V2C_8 (V2C_389_86),
	.V2C_9 (V2C_526_86),
	.V2C_10 (V2C_638_86),
	.V2C_11 (V2C_699_86),
	.V2C_12 (V2C_819_86),
	.V2C_13 (V2C_909_86),
	.V2C_14 (V2C_924_86),
	.V2C_15 (V2C_1003_86),
	.V2C_16 (V2C_1035_86),
	.V2C_17 (V2C_1102_86),
	.V2C_18 (V2C_1133_86),
	.V2C_19 (V2C_1237_86),
	.V2C_20 (V2C_1238_86),
	.C2V_1 (C2V_86_28),
	.C2V_2 (C2V_86_77),
	.C2V_3 (C2V_86_133),
	.C2V_4 (C2V_86_181),
	.C2V_5 (C2V_86_210),
	.C2V_6 (C2V_86_279),
	.C2V_7 (C2V_86_330),
	.C2V_8 (C2V_86_389),
	.C2V_9 (C2V_86_526),
	.C2V_10 (C2V_86_638),
	.C2V_11 (C2V_86_699),
	.C2V_12 (C2V_86_819),
	.C2V_13 (C2V_86_909),
	.C2V_14 (C2V_86_924),
	.C2V_15 (C2V_86_1003),
	.C2V_16 (C2V_86_1035),
	.C2V_17 (C2V_86_1102),
	.C2V_18 (C2V_86_1133),
	.C2V_19 (C2V_86_1237),
	.C2V_20 (C2V_86_1238),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU87 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_23_87),
	.V2C_2 (V2C_50_87),
	.V2C_3 (V2C_115_87),
	.V2C_4 (V2C_149_87),
	.V2C_5 (V2C_215_87),
	.V2C_6 (V2C_282_87),
	.V2C_7 (V2C_379_87),
	.V2C_8 (V2C_386_87),
	.V2C_9 (V2C_545_87),
	.V2C_10 (V2C_602_87),
	.V2C_11 (V2C_630_87),
	.V2C_12 (V2C_734_87),
	.V2C_13 (V2C_865_87),
	.V2C_14 (V2C_957_87),
	.V2C_15 (V2C_982_87),
	.V2C_16 (V2C_1042_87),
	.V2C_17 (V2C_1072_87),
	.V2C_18 (V2C_1117_87),
	.V2C_19 (V2C_1238_87),
	.V2C_20 (V2C_1239_87),
	.C2V_1 (C2V_87_23),
	.C2V_2 (C2V_87_50),
	.C2V_3 (C2V_87_115),
	.C2V_4 (C2V_87_149),
	.C2V_5 (C2V_87_215),
	.C2V_6 (C2V_87_282),
	.C2V_7 (C2V_87_379),
	.C2V_8 (C2V_87_386),
	.C2V_9 (C2V_87_545),
	.C2V_10 (C2V_87_602),
	.C2V_11 (C2V_87_630),
	.C2V_12 (C2V_87_734),
	.C2V_13 (C2V_87_865),
	.C2V_14 (C2V_87_957),
	.C2V_15 (C2V_87_982),
	.C2V_16 (C2V_87_1042),
	.C2V_17 (C2V_87_1072),
	.C2V_18 (C2V_87_1117),
	.C2V_19 (C2V_87_1238),
	.C2V_20 (C2V_87_1239),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU88 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_42_88),
	.V2C_2 (V2C_53_88),
	.V2C_3 (V2C_140_88),
	.V2C_4 (V2C_148_88),
	.V2C_5 (V2C_213_88),
	.V2C_6 (V2C_267_88),
	.V2C_7 (V2C_443_88),
	.V2C_8 (V2C_483_88),
	.V2C_9 (V2C_567_88),
	.V2C_10 (V2C_581_88),
	.V2C_11 (V2C_654_88),
	.V2C_12 (V2C_700_88),
	.V2C_13 (V2C_869_88),
	.V2C_14 (V2C_941_88),
	.V2C_15 (V2C_977_88),
	.V2C_16 (V2C_1055_88),
	.V2C_17 (V2C_1082_88),
	.V2C_18 (V2C_1146_88),
	.V2C_19 (V2C_1239_88),
	.V2C_20 (V2C_1240_88),
	.C2V_1 (C2V_88_42),
	.C2V_2 (C2V_88_53),
	.C2V_3 (C2V_88_140),
	.C2V_4 (C2V_88_148),
	.C2V_5 (C2V_88_213),
	.C2V_6 (C2V_88_267),
	.C2V_7 (C2V_88_443),
	.C2V_8 (C2V_88_483),
	.C2V_9 (C2V_88_567),
	.C2V_10 (C2V_88_581),
	.C2V_11 (C2V_88_654),
	.C2V_12 (C2V_88_700),
	.C2V_13 (C2V_88_869),
	.C2V_14 (C2V_88_941),
	.C2V_15 (C2V_88_977),
	.C2V_16 (C2V_88_1055),
	.C2V_17 (C2V_88_1082),
	.C2V_18 (C2V_88_1146),
	.C2V_19 (C2V_88_1239),
	.C2V_20 (C2V_88_1240),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU89 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_13_89),
	.V2C_2 (V2C_71_89),
	.V2C_3 (V2C_106_89),
	.V2C_4 (V2C_177_89),
	.V2C_5 (V2C_193_89),
	.V2C_6 (V2C_259_89),
	.V2C_7 (V2C_308_89),
	.V2C_8 (V2C_375_89),
	.V2C_9 (V2C_454_89),
	.V2C_10 (V2C_688_89),
	.V2C_11 (V2C_752_89),
	.V2C_12 (V2C_806_89),
	.V2C_13 (V2C_884_89),
	.V2C_14 (V2C_932_89),
	.V2C_15 (V2C_975_89),
	.V2C_16 (V2C_1027_89),
	.V2C_17 (V2C_1076_89),
	.V2C_18 (V2C_1124_89),
	.V2C_19 (V2C_1240_89),
	.V2C_20 (V2C_1241_89),
	.C2V_1 (C2V_89_13),
	.C2V_2 (C2V_89_71),
	.C2V_3 (C2V_89_106),
	.C2V_4 (C2V_89_177),
	.C2V_5 (C2V_89_193),
	.C2V_6 (C2V_89_259),
	.C2V_7 (C2V_89_308),
	.C2V_8 (C2V_89_375),
	.C2V_9 (C2V_89_454),
	.C2V_10 (C2V_89_688),
	.C2V_11 (C2V_89_752),
	.C2V_12 (C2V_89_806),
	.C2V_13 (C2V_89_884),
	.C2V_14 (C2V_89_932),
	.C2V_15 (C2V_89_975),
	.C2V_16 (C2V_89_1027),
	.C2V_17 (C2V_89_1076),
	.C2V_18 (C2V_89_1124),
	.C2V_19 (C2V_89_1240),
	.C2V_20 (C2V_89_1241),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU90 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_44_90),
	.V2C_2 (V2C_68_90),
	.V2C_3 (V2C_108_90),
	.V2C_4 (V2C_176_90),
	.V2C_5 (V2C_210_90),
	.V2C_6 (V2C_241_90),
	.V2C_7 (V2C_294_90),
	.V2C_8 (V2C_446_90),
	.V2C_9 (V2C_543_90),
	.V2C_10 (V2C_624_90),
	.V2C_11 (V2C_780_90),
	.V2C_12 (V2C_856_90),
	.V2C_13 (V2C_889_90),
	.V2C_14 (V2C_951_90),
	.V2C_15 (V2C_986_90),
	.V2C_16 (V2C_1053_90),
	.V2C_17 (V2C_1069_90),
	.V2C_18 (V2C_1119_90),
	.V2C_19 (V2C_1241_90),
	.V2C_20 (V2C_1242_90),
	.C2V_1 (C2V_90_44),
	.C2V_2 (C2V_90_68),
	.C2V_3 (C2V_90_108),
	.C2V_4 (C2V_90_176),
	.C2V_5 (C2V_90_210),
	.C2V_6 (C2V_90_241),
	.C2V_7 (C2V_90_294),
	.C2V_8 (C2V_90_446),
	.C2V_9 (C2V_90_543),
	.C2V_10 (C2V_90_624),
	.C2V_11 (C2V_90_780),
	.C2V_12 (C2V_90_856),
	.C2V_13 (C2V_90_889),
	.C2V_14 (C2V_90_951),
	.C2V_15 (C2V_90_986),
	.C2V_16 (C2V_90_1053),
	.C2V_17 (C2V_90_1069),
	.C2V_18 (C2V_90_1119),
	.C2V_19 (C2V_90_1241),
	.C2V_20 (C2V_90_1242),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU91 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_20_91),
	.V2C_2 (V2C_56_91),
	.V2C_3 (V2C_124_91),
	.V2C_4 (V2C_185_91),
	.V2C_5 (V2C_199_91),
	.V2C_6 (V2C_242_91),
	.V2C_7 (V2C_342_91),
	.V2C_8 (V2C_396_91),
	.V2C_9 (V2C_493_91),
	.V2C_10 (V2C_729_91),
	.V2C_11 (V2C_777_91),
	.V2C_12 (V2C_825_91),
	.V2C_13 (V2C_866_91),
	.V2C_14 (V2C_955_91),
	.V2C_15 (V2C_989_91),
	.V2C_16 (V2C_1028_91),
	.V2C_17 (V2C_1102_91),
	.V2C_18 (V2C_1113_91),
	.V2C_19 (V2C_1242_91),
	.V2C_20 (V2C_1243_91),
	.C2V_1 (C2V_91_20),
	.C2V_2 (C2V_91_56),
	.C2V_3 (C2V_91_124),
	.C2V_4 (C2V_91_185),
	.C2V_5 (C2V_91_199),
	.C2V_6 (C2V_91_242),
	.C2V_7 (C2V_91_342),
	.C2V_8 (C2V_91_396),
	.C2V_9 (C2V_91_493),
	.C2V_10 (C2V_91_729),
	.C2V_11 (C2V_91_777),
	.C2V_12 (C2V_91_825),
	.C2V_13 (C2V_91_866),
	.C2V_14 (C2V_91_955),
	.C2V_15 (C2V_91_989),
	.C2V_16 (C2V_91_1028),
	.C2V_17 (C2V_91_1102),
	.C2V_18 (C2V_91_1113),
	.C2V_19 (C2V_91_1242),
	.C2V_20 (C2V_91_1243),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU92 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_29_92),
	.V2C_2 (V2C_78_92),
	.V2C_3 (V2C_134_92),
	.V2C_4 (V2C_182_92),
	.V2C_5 (V2C_211_92),
	.V2C_6 (V2C_280_92),
	.V2C_7 (V2C_331_92),
	.V2C_8 (V2C_390_92),
	.V2C_9 (V2C_527_92),
	.V2C_10 (V2C_639_92),
	.V2C_11 (V2C_700_92),
	.V2C_12 (V2C_820_92),
	.V2C_13 (V2C_910_92),
	.V2C_14 (V2C_925_92),
	.V2C_15 (V2C_1004_92),
	.V2C_16 (V2C_1036_92),
	.V2C_17 (V2C_1103_92),
	.V2C_18 (V2C_1134_92),
	.V2C_19 (V2C_1243_92),
	.V2C_20 (V2C_1244_92),
	.C2V_1 (C2V_92_29),
	.C2V_2 (C2V_92_78),
	.C2V_3 (C2V_92_134),
	.C2V_4 (C2V_92_182),
	.C2V_5 (C2V_92_211),
	.C2V_6 (C2V_92_280),
	.C2V_7 (C2V_92_331),
	.C2V_8 (C2V_92_390),
	.C2V_9 (C2V_92_527),
	.C2V_10 (C2V_92_639),
	.C2V_11 (C2V_92_700),
	.C2V_12 (C2V_92_820),
	.C2V_13 (C2V_92_910),
	.C2V_14 (C2V_92_925),
	.C2V_15 (C2V_92_1004),
	.C2V_16 (C2V_92_1036),
	.C2V_17 (C2V_92_1103),
	.C2V_18 (C2V_92_1134),
	.C2V_19 (C2V_92_1243),
	.C2V_20 (C2V_92_1244),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU93 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_24_93),
	.V2C_2 (V2C_51_93),
	.V2C_3 (V2C_116_93),
	.V2C_4 (V2C_150_93),
	.V2C_5 (V2C_216_93),
	.V2C_6 (V2C_283_93),
	.V2C_7 (V2C_380_93),
	.V2C_8 (V2C_387_93),
	.V2C_9 (V2C_546_93),
	.V2C_10 (V2C_603_93),
	.V2C_11 (V2C_631_93),
	.V2C_12 (V2C_735_93),
	.V2C_13 (V2C_866_93),
	.V2C_14 (V2C_958_93),
	.V2C_15 (V2C_983_93),
	.V2C_16 (V2C_1043_93),
	.V2C_17 (V2C_1073_93),
	.V2C_18 (V2C_1118_93),
	.V2C_19 (V2C_1244_93),
	.V2C_20 (V2C_1245_93),
	.C2V_1 (C2V_93_24),
	.C2V_2 (C2V_93_51),
	.C2V_3 (C2V_93_116),
	.C2V_4 (C2V_93_150),
	.C2V_5 (C2V_93_216),
	.C2V_6 (C2V_93_283),
	.C2V_7 (C2V_93_380),
	.C2V_8 (C2V_93_387),
	.C2V_9 (C2V_93_546),
	.C2V_10 (C2V_93_603),
	.C2V_11 (C2V_93_631),
	.C2V_12 (C2V_93_735),
	.C2V_13 (C2V_93_866),
	.C2V_14 (C2V_93_958),
	.C2V_15 (C2V_93_983),
	.C2V_16 (C2V_93_1043),
	.C2V_17 (C2V_93_1073),
	.C2V_18 (C2V_93_1118),
	.C2V_19 (C2V_93_1244),
	.C2V_20 (C2V_93_1245),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU94 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_43_94),
	.V2C_2 (V2C_54_94),
	.V2C_3 (V2C_141_94),
	.V2C_4 (V2C_149_94),
	.V2C_5 (V2C_214_94),
	.V2C_6 (V2C_268_94),
	.V2C_7 (V2C_444_94),
	.V2C_8 (V2C_484_94),
	.V2C_9 (V2C_568_94),
	.V2C_10 (V2C_582_94),
	.V2C_11 (V2C_655_94),
	.V2C_12 (V2C_701_94),
	.V2C_13 (V2C_870_94),
	.V2C_14 (V2C_942_94),
	.V2C_15 (V2C_978_94),
	.V2C_16 (V2C_1056_94),
	.V2C_17 (V2C_1083_94),
	.V2C_18 (V2C_1147_94),
	.V2C_19 (V2C_1245_94),
	.V2C_20 (V2C_1246_94),
	.C2V_1 (C2V_94_43),
	.C2V_2 (C2V_94_54),
	.C2V_3 (C2V_94_141),
	.C2V_4 (C2V_94_149),
	.C2V_5 (C2V_94_214),
	.C2V_6 (C2V_94_268),
	.C2V_7 (C2V_94_444),
	.C2V_8 (C2V_94_484),
	.C2V_9 (C2V_94_568),
	.C2V_10 (C2V_94_582),
	.C2V_11 (C2V_94_655),
	.C2V_12 (C2V_94_701),
	.C2V_13 (C2V_94_870),
	.C2V_14 (C2V_94_942),
	.C2V_15 (C2V_94_978),
	.C2V_16 (C2V_94_1056),
	.C2V_17 (C2V_94_1083),
	.C2V_18 (C2V_94_1147),
	.C2V_19 (C2V_94_1245),
	.C2V_20 (C2V_94_1246),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU95 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_14_95),
	.V2C_2 (V2C_72_95),
	.V2C_3 (V2C_107_95),
	.V2C_4 (V2C_178_95),
	.V2C_5 (V2C_194_95),
	.V2C_6 (V2C_260_95),
	.V2C_7 (V2C_309_95),
	.V2C_8 (V2C_376_95),
	.V2C_9 (V2C_455_95),
	.V2C_10 (V2C_689_95),
	.V2C_11 (V2C_753_95),
	.V2C_12 (V2C_807_95),
	.V2C_13 (V2C_885_95),
	.V2C_14 (V2C_933_95),
	.V2C_15 (V2C_976_95),
	.V2C_16 (V2C_1028_95),
	.V2C_17 (V2C_1077_95),
	.V2C_18 (V2C_1125_95),
	.V2C_19 (V2C_1246_95),
	.V2C_20 (V2C_1247_95),
	.C2V_1 (C2V_95_14),
	.C2V_2 (C2V_95_72),
	.C2V_3 (C2V_95_107),
	.C2V_4 (C2V_95_178),
	.C2V_5 (C2V_95_194),
	.C2V_6 (C2V_95_260),
	.C2V_7 (C2V_95_309),
	.C2V_8 (C2V_95_376),
	.C2V_9 (C2V_95_455),
	.C2V_10 (C2V_95_689),
	.C2V_11 (C2V_95_753),
	.C2V_12 (C2V_95_807),
	.C2V_13 (C2V_95_885),
	.C2V_14 (C2V_95_933),
	.C2V_15 (C2V_95_976),
	.C2V_16 (C2V_95_1028),
	.C2V_17 (C2V_95_1077),
	.C2V_18 (C2V_95_1125),
	.C2V_19 (C2V_95_1246),
	.C2V_20 (C2V_95_1247),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU96 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_45_96),
	.V2C_2 (V2C_69_96),
	.V2C_3 (V2C_109_96),
	.V2C_4 (V2C_177_96),
	.V2C_5 (V2C_211_96),
	.V2C_6 (V2C_242_96),
	.V2C_7 (V2C_295_96),
	.V2C_8 (V2C_447_96),
	.V2C_9 (V2C_544_96),
	.V2C_10 (V2C_577_96),
	.V2C_11 (V2C_781_96),
	.V2C_12 (V2C_857_96),
	.V2C_13 (V2C_890_96),
	.V2C_14 (V2C_952_96),
	.V2C_15 (V2C_987_96),
	.V2C_16 (V2C_1054_96),
	.V2C_17 (V2C_1070_96),
	.V2C_18 (V2C_1120_96),
	.V2C_19 (V2C_1247_96),
	.V2C_20 (V2C_1248_96),
	.C2V_1 (C2V_96_45),
	.C2V_2 (C2V_96_69),
	.C2V_3 (C2V_96_109),
	.C2V_4 (C2V_96_177),
	.C2V_5 (C2V_96_211),
	.C2V_6 (C2V_96_242),
	.C2V_7 (C2V_96_295),
	.C2V_8 (C2V_96_447),
	.C2V_9 (C2V_96_544),
	.C2V_10 (C2V_96_577),
	.C2V_11 (C2V_96_781),
	.C2V_12 (C2V_96_857),
	.C2V_13 (C2V_96_890),
	.C2V_14 (C2V_96_952),
	.C2V_15 (C2V_96_987),
	.C2V_16 (C2V_96_1054),
	.C2V_17 (C2V_96_1070),
	.C2V_18 (C2V_96_1120),
	.C2V_19 (C2V_96_1247),
	.C2V_20 (C2V_96_1248),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU97 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_21_97),
	.V2C_2 (V2C_57_97),
	.V2C_3 (V2C_125_97),
	.V2C_4 (V2C_186_97),
	.V2C_5 (V2C_200_97),
	.V2C_6 (V2C_243_97),
	.V2C_7 (V2C_343_97),
	.V2C_8 (V2C_397_97),
	.V2C_9 (V2C_494_97),
	.V2C_10 (V2C_730_97),
	.V2C_11 (V2C_778_97),
	.V2C_12 (V2C_826_97),
	.V2C_13 (V2C_867_97),
	.V2C_14 (V2C_956_97),
	.V2C_15 (V2C_990_97),
	.V2C_16 (V2C_1029_97),
	.V2C_17 (V2C_1103_97),
	.V2C_18 (V2C_1114_97),
	.V2C_19 (V2C_1248_97),
	.V2C_20 (V2C_1249_97),
	.C2V_1 (C2V_97_21),
	.C2V_2 (C2V_97_57),
	.C2V_3 (C2V_97_125),
	.C2V_4 (C2V_97_186),
	.C2V_5 (C2V_97_200),
	.C2V_6 (C2V_97_243),
	.C2V_7 (C2V_97_343),
	.C2V_8 (C2V_97_397),
	.C2V_9 (C2V_97_494),
	.C2V_10 (C2V_97_730),
	.C2V_11 (C2V_97_778),
	.C2V_12 (C2V_97_826),
	.C2V_13 (C2V_97_867),
	.C2V_14 (C2V_97_956),
	.C2V_15 (C2V_97_990),
	.C2V_16 (C2V_97_1029),
	.C2V_17 (C2V_97_1103),
	.C2V_18 (C2V_97_1114),
	.C2V_19 (C2V_97_1248),
	.C2V_20 (C2V_97_1249),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU98 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_30_98),
	.V2C_2 (V2C_79_98),
	.V2C_3 (V2C_135_98),
	.V2C_4 (V2C_183_98),
	.V2C_5 (V2C_212_98),
	.V2C_6 (V2C_281_98),
	.V2C_7 (V2C_332_98),
	.V2C_8 (V2C_391_98),
	.V2C_9 (V2C_528_98),
	.V2C_10 (V2C_640_98),
	.V2C_11 (V2C_701_98),
	.V2C_12 (V2C_821_98),
	.V2C_13 (V2C_911_98),
	.V2C_14 (V2C_926_98),
	.V2C_15 (V2C_1005_98),
	.V2C_16 (V2C_1037_98),
	.V2C_17 (V2C_1104_98),
	.V2C_18 (V2C_1135_98),
	.V2C_19 (V2C_1249_98),
	.V2C_20 (V2C_1250_98),
	.C2V_1 (C2V_98_30),
	.C2V_2 (C2V_98_79),
	.C2V_3 (C2V_98_135),
	.C2V_4 (C2V_98_183),
	.C2V_5 (C2V_98_212),
	.C2V_6 (C2V_98_281),
	.C2V_7 (C2V_98_332),
	.C2V_8 (C2V_98_391),
	.C2V_9 (C2V_98_528),
	.C2V_10 (C2V_98_640),
	.C2V_11 (C2V_98_701),
	.C2V_12 (C2V_98_821),
	.C2V_13 (C2V_98_911),
	.C2V_14 (C2V_98_926),
	.C2V_15 (C2V_98_1005),
	.C2V_16 (C2V_98_1037),
	.C2V_17 (C2V_98_1104),
	.C2V_18 (C2V_98_1135),
	.C2V_19 (C2V_98_1249),
	.C2V_20 (C2V_98_1250),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU99 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_25_99),
	.V2C_2 (V2C_52_99),
	.V2C_3 (V2C_117_99),
	.V2C_4 (V2C_151_99),
	.V2C_5 (V2C_217_99),
	.V2C_6 (V2C_284_99),
	.V2C_7 (V2C_381_99),
	.V2C_8 (V2C_388_99),
	.V2C_9 (V2C_547_99),
	.V2C_10 (V2C_604_99),
	.V2C_11 (V2C_632_99),
	.V2C_12 (V2C_736_99),
	.V2C_13 (V2C_867_99),
	.V2C_14 (V2C_959_99),
	.V2C_15 (V2C_984_99),
	.V2C_16 (V2C_1044_99),
	.V2C_17 (V2C_1074_99),
	.V2C_18 (V2C_1119_99),
	.V2C_19 (V2C_1250_99),
	.V2C_20 (V2C_1251_99),
	.C2V_1 (C2V_99_25),
	.C2V_2 (C2V_99_52),
	.C2V_3 (C2V_99_117),
	.C2V_4 (C2V_99_151),
	.C2V_5 (C2V_99_217),
	.C2V_6 (C2V_99_284),
	.C2V_7 (C2V_99_381),
	.C2V_8 (C2V_99_388),
	.C2V_9 (C2V_99_547),
	.C2V_10 (C2V_99_604),
	.C2V_11 (C2V_99_632),
	.C2V_12 (C2V_99_736),
	.C2V_13 (C2V_99_867),
	.C2V_14 (C2V_99_959),
	.C2V_15 (C2V_99_984),
	.C2V_16 (C2V_99_1044),
	.C2V_17 (C2V_99_1074),
	.C2V_18 (C2V_99_1119),
	.C2V_19 (C2V_99_1250),
	.C2V_20 (C2V_99_1251),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU100 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_44_100),
	.V2C_2 (V2C_55_100),
	.V2C_3 (V2C_142_100),
	.V2C_4 (V2C_150_100),
	.V2C_5 (V2C_215_100),
	.V2C_6 (V2C_269_100),
	.V2C_7 (V2C_445_100),
	.V2C_8 (V2C_485_100),
	.V2C_9 (V2C_569_100),
	.V2C_10 (V2C_583_100),
	.V2C_11 (V2C_656_100),
	.V2C_12 (V2C_702_100),
	.V2C_13 (V2C_871_100),
	.V2C_14 (V2C_943_100),
	.V2C_15 (V2C_979_100),
	.V2C_16 (V2C_1009_100),
	.V2C_17 (V2C_1084_100),
	.V2C_18 (V2C_1148_100),
	.V2C_19 (V2C_1251_100),
	.V2C_20 (V2C_1252_100),
	.C2V_1 (C2V_100_44),
	.C2V_2 (C2V_100_55),
	.C2V_3 (C2V_100_142),
	.C2V_4 (C2V_100_150),
	.C2V_5 (C2V_100_215),
	.C2V_6 (C2V_100_269),
	.C2V_7 (C2V_100_445),
	.C2V_8 (C2V_100_485),
	.C2V_9 (C2V_100_569),
	.C2V_10 (C2V_100_583),
	.C2V_11 (C2V_100_656),
	.C2V_12 (C2V_100_702),
	.C2V_13 (C2V_100_871),
	.C2V_14 (C2V_100_943),
	.C2V_15 (C2V_100_979),
	.C2V_16 (C2V_100_1009),
	.C2V_17 (C2V_100_1084),
	.C2V_18 (C2V_100_1148),
	.C2V_19 (C2V_100_1251),
	.C2V_20 (C2V_100_1252),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU101 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_15_101),
	.V2C_2 (V2C_73_101),
	.V2C_3 (V2C_108_101),
	.V2C_4 (V2C_179_101),
	.V2C_5 (V2C_195_101),
	.V2C_6 (V2C_261_101),
	.V2C_7 (V2C_310_101),
	.V2C_8 (V2C_377_101),
	.V2C_9 (V2C_456_101),
	.V2C_10 (V2C_690_101),
	.V2C_11 (V2C_754_101),
	.V2C_12 (V2C_808_101),
	.V2C_13 (V2C_886_101),
	.V2C_14 (V2C_934_101),
	.V2C_15 (V2C_977_101),
	.V2C_16 (V2C_1029_101),
	.V2C_17 (V2C_1078_101),
	.V2C_18 (V2C_1126_101),
	.V2C_19 (V2C_1252_101),
	.V2C_20 (V2C_1253_101),
	.C2V_1 (C2V_101_15),
	.C2V_2 (C2V_101_73),
	.C2V_3 (C2V_101_108),
	.C2V_4 (C2V_101_179),
	.C2V_5 (C2V_101_195),
	.C2V_6 (C2V_101_261),
	.C2V_7 (C2V_101_310),
	.C2V_8 (C2V_101_377),
	.C2V_9 (C2V_101_456),
	.C2V_10 (C2V_101_690),
	.C2V_11 (C2V_101_754),
	.C2V_12 (C2V_101_808),
	.C2V_13 (C2V_101_886),
	.C2V_14 (C2V_101_934),
	.C2V_15 (C2V_101_977),
	.C2V_16 (C2V_101_1029),
	.C2V_17 (C2V_101_1078),
	.C2V_18 (C2V_101_1126),
	.C2V_19 (C2V_101_1252),
	.C2V_20 (C2V_101_1253),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU102 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_46_102),
	.V2C_2 (V2C_70_102),
	.V2C_3 (V2C_110_102),
	.V2C_4 (V2C_178_102),
	.V2C_5 (V2C_212_102),
	.V2C_6 (V2C_243_102),
	.V2C_7 (V2C_296_102),
	.V2C_8 (V2C_448_102),
	.V2C_9 (V2C_545_102),
	.V2C_10 (V2C_578_102),
	.V2C_11 (V2C_782_102),
	.V2C_12 (V2C_858_102),
	.V2C_13 (V2C_891_102),
	.V2C_14 (V2C_953_102),
	.V2C_15 (V2C_988_102),
	.V2C_16 (V2C_1055_102),
	.V2C_17 (V2C_1071_102),
	.V2C_18 (V2C_1121_102),
	.V2C_19 (V2C_1253_102),
	.V2C_20 (V2C_1254_102),
	.C2V_1 (C2V_102_46),
	.C2V_2 (C2V_102_70),
	.C2V_3 (C2V_102_110),
	.C2V_4 (C2V_102_178),
	.C2V_5 (C2V_102_212),
	.C2V_6 (C2V_102_243),
	.C2V_7 (C2V_102_296),
	.C2V_8 (C2V_102_448),
	.C2V_9 (C2V_102_545),
	.C2V_10 (C2V_102_578),
	.C2V_11 (C2V_102_782),
	.C2V_12 (C2V_102_858),
	.C2V_13 (C2V_102_891),
	.C2V_14 (C2V_102_953),
	.C2V_15 (C2V_102_988),
	.C2V_16 (C2V_102_1055),
	.C2V_17 (C2V_102_1071),
	.C2V_18 (C2V_102_1121),
	.C2V_19 (C2V_102_1253),
	.C2V_20 (C2V_102_1254),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU103 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_22_103),
	.V2C_2 (V2C_58_103),
	.V2C_3 (V2C_126_103),
	.V2C_4 (V2C_187_103),
	.V2C_5 (V2C_201_103),
	.V2C_6 (V2C_244_103),
	.V2C_7 (V2C_344_103),
	.V2C_8 (V2C_398_103),
	.V2C_9 (V2C_495_103),
	.V2C_10 (V2C_731_103),
	.V2C_11 (V2C_779_103),
	.V2C_12 (V2C_827_103),
	.V2C_13 (V2C_868_103),
	.V2C_14 (V2C_957_103),
	.V2C_15 (V2C_991_103),
	.V2C_16 (V2C_1030_103),
	.V2C_17 (V2C_1104_103),
	.V2C_18 (V2C_1115_103),
	.V2C_19 (V2C_1254_103),
	.V2C_20 (V2C_1255_103),
	.C2V_1 (C2V_103_22),
	.C2V_2 (C2V_103_58),
	.C2V_3 (C2V_103_126),
	.C2V_4 (C2V_103_187),
	.C2V_5 (C2V_103_201),
	.C2V_6 (C2V_103_244),
	.C2V_7 (C2V_103_344),
	.C2V_8 (C2V_103_398),
	.C2V_9 (C2V_103_495),
	.C2V_10 (C2V_103_731),
	.C2V_11 (C2V_103_779),
	.C2V_12 (C2V_103_827),
	.C2V_13 (C2V_103_868),
	.C2V_14 (C2V_103_957),
	.C2V_15 (C2V_103_991),
	.C2V_16 (C2V_103_1030),
	.C2V_17 (C2V_103_1104),
	.C2V_18 (C2V_103_1115),
	.C2V_19 (C2V_103_1254),
	.C2V_20 (C2V_103_1255),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU104 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_31_104),
	.V2C_2 (V2C_80_104),
	.V2C_3 (V2C_136_104),
	.V2C_4 (V2C_184_104),
	.V2C_5 (V2C_213_104),
	.V2C_6 (V2C_282_104),
	.V2C_7 (V2C_333_104),
	.V2C_8 (V2C_392_104),
	.V2C_9 (V2C_481_104),
	.V2C_10 (V2C_641_104),
	.V2C_11 (V2C_702_104),
	.V2C_12 (V2C_822_104),
	.V2C_13 (V2C_912_104),
	.V2C_14 (V2C_927_104),
	.V2C_15 (V2C_1006_104),
	.V2C_16 (V2C_1038_104),
	.V2C_17 (V2C_1057_104),
	.V2C_18 (V2C_1136_104),
	.V2C_19 (V2C_1255_104),
	.V2C_20 (V2C_1256_104),
	.C2V_1 (C2V_104_31),
	.C2V_2 (C2V_104_80),
	.C2V_3 (C2V_104_136),
	.C2V_4 (C2V_104_184),
	.C2V_5 (C2V_104_213),
	.C2V_6 (C2V_104_282),
	.C2V_7 (C2V_104_333),
	.C2V_8 (C2V_104_392),
	.C2V_9 (C2V_104_481),
	.C2V_10 (C2V_104_641),
	.C2V_11 (C2V_104_702),
	.C2V_12 (C2V_104_822),
	.C2V_13 (C2V_104_912),
	.C2V_14 (C2V_104_927),
	.C2V_15 (C2V_104_1006),
	.C2V_16 (C2V_104_1038),
	.C2V_17 (C2V_104_1057),
	.C2V_18 (C2V_104_1136),
	.C2V_19 (C2V_104_1255),
	.C2V_20 (C2V_104_1256),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU105 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_26_105),
	.V2C_2 (V2C_53_105),
	.V2C_3 (V2C_118_105),
	.V2C_4 (V2C_152_105),
	.V2C_5 (V2C_218_105),
	.V2C_6 (V2C_285_105),
	.V2C_7 (V2C_382_105),
	.V2C_8 (V2C_389_105),
	.V2C_9 (V2C_548_105),
	.V2C_10 (V2C_605_105),
	.V2C_11 (V2C_633_105),
	.V2C_12 (V2C_737_105),
	.V2C_13 (V2C_868_105),
	.V2C_14 (V2C_960_105),
	.V2C_15 (V2C_985_105),
	.V2C_16 (V2C_1045_105),
	.V2C_17 (V2C_1075_105),
	.V2C_18 (V2C_1120_105),
	.V2C_19 (V2C_1256_105),
	.V2C_20 (V2C_1257_105),
	.C2V_1 (C2V_105_26),
	.C2V_2 (C2V_105_53),
	.C2V_3 (C2V_105_118),
	.C2V_4 (C2V_105_152),
	.C2V_5 (C2V_105_218),
	.C2V_6 (C2V_105_285),
	.C2V_7 (C2V_105_382),
	.C2V_8 (C2V_105_389),
	.C2V_9 (C2V_105_548),
	.C2V_10 (C2V_105_605),
	.C2V_11 (C2V_105_633),
	.C2V_12 (C2V_105_737),
	.C2V_13 (C2V_105_868),
	.C2V_14 (C2V_105_960),
	.C2V_15 (C2V_105_985),
	.C2V_16 (C2V_105_1045),
	.C2V_17 (C2V_105_1075),
	.C2V_18 (C2V_105_1120),
	.C2V_19 (C2V_105_1256),
	.C2V_20 (C2V_105_1257),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU106 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_45_106),
	.V2C_2 (V2C_56_106),
	.V2C_3 (V2C_143_106),
	.V2C_4 (V2C_151_106),
	.V2C_5 (V2C_216_106),
	.V2C_6 (V2C_270_106),
	.V2C_7 (V2C_446_106),
	.V2C_8 (V2C_486_106),
	.V2C_9 (V2C_570_106),
	.V2C_10 (V2C_584_106),
	.V2C_11 (V2C_657_106),
	.V2C_12 (V2C_703_106),
	.V2C_13 (V2C_872_106),
	.V2C_14 (V2C_944_106),
	.V2C_15 (V2C_980_106),
	.V2C_16 (V2C_1010_106),
	.V2C_17 (V2C_1085_106),
	.V2C_18 (V2C_1149_106),
	.V2C_19 (V2C_1257_106),
	.V2C_20 (V2C_1258_106),
	.C2V_1 (C2V_106_45),
	.C2V_2 (C2V_106_56),
	.C2V_3 (C2V_106_143),
	.C2V_4 (C2V_106_151),
	.C2V_5 (C2V_106_216),
	.C2V_6 (C2V_106_270),
	.C2V_7 (C2V_106_446),
	.C2V_8 (C2V_106_486),
	.C2V_9 (C2V_106_570),
	.C2V_10 (C2V_106_584),
	.C2V_11 (C2V_106_657),
	.C2V_12 (C2V_106_703),
	.C2V_13 (C2V_106_872),
	.C2V_14 (C2V_106_944),
	.C2V_15 (C2V_106_980),
	.C2V_16 (C2V_106_1010),
	.C2V_17 (C2V_106_1085),
	.C2V_18 (C2V_106_1149),
	.C2V_19 (C2V_106_1257),
	.C2V_20 (C2V_106_1258),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU107 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_16_107),
	.V2C_2 (V2C_74_107),
	.V2C_3 (V2C_109_107),
	.V2C_4 (V2C_180_107),
	.V2C_5 (V2C_196_107),
	.V2C_6 (V2C_262_107),
	.V2C_7 (V2C_311_107),
	.V2C_8 (V2C_378_107),
	.V2C_9 (V2C_457_107),
	.V2C_10 (V2C_691_107),
	.V2C_11 (V2C_755_107),
	.V2C_12 (V2C_809_107),
	.V2C_13 (V2C_887_107),
	.V2C_14 (V2C_935_107),
	.V2C_15 (V2C_978_107),
	.V2C_16 (V2C_1030_107),
	.V2C_17 (V2C_1079_107),
	.V2C_18 (V2C_1127_107),
	.V2C_19 (V2C_1258_107),
	.V2C_20 (V2C_1259_107),
	.C2V_1 (C2V_107_16),
	.C2V_2 (C2V_107_74),
	.C2V_3 (C2V_107_109),
	.C2V_4 (C2V_107_180),
	.C2V_5 (C2V_107_196),
	.C2V_6 (C2V_107_262),
	.C2V_7 (C2V_107_311),
	.C2V_8 (C2V_107_378),
	.C2V_9 (C2V_107_457),
	.C2V_10 (C2V_107_691),
	.C2V_11 (C2V_107_755),
	.C2V_12 (C2V_107_809),
	.C2V_13 (C2V_107_887),
	.C2V_14 (C2V_107_935),
	.C2V_15 (C2V_107_978),
	.C2V_16 (C2V_107_1030),
	.C2V_17 (C2V_107_1079),
	.C2V_18 (C2V_107_1127),
	.C2V_19 (C2V_107_1258),
	.C2V_20 (C2V_107_1259),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU108 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_47_108),
	.V2C_2 (V2C_71_108),
	.V2C_3 (V2C_111_108),
	.V2C_4 (V2C_179_108),
	.V2C_5 (V2C_213_108),
	.V2C_6 (V2C_244_108),
	.V2C_7 (V2C_297_108),
	.V2C_8 (V2C_449_108),
	.V2C_9 (V2C_546_108),
	.V2C_10 (V2C_579_108),
	.V2C_11 (V2C_783_108),
	.V2C_12 (V2C_859_108),
	.V2C_13 (V2C_892_108),
	.V2C_14 (V2C_954_108),
	.V2C_15 (V2C_989_108),
	.V2C_16 (V2C_1056_108),
	.V2C_17 (V2C_1072_108),
	.V2C_18 (V2C_1122_108),
	.V2C_19 (V2C_1259_108),
	.V2C_20 (V2C_1260_108),
	.C2V_1 (C2V_108_47),
	.C2V_2 (C2V_108_71),
	.C2V_3 (C2V_108_111),
	.C2V_4 (C2V_108_179),
	.C2V_5 (C2V_108_213),
	.C2V_6 (C2V_108_244),
	.C2V_7 (C2V_108_297),
	.C2V_8 (C2V_108_449),
	.C2V_9 (C2V_108_546),
	.C2V_10 (C2V_108_579),
	.C2V_11 (C2V_108_783),
	.C2V_12 (C2V_108_859),
	.C2V_13 (C2V_108_892),
	.C2V_14 (C2V_108_954),
	.C2V_15 (C2V_108_989),
	.C2V_16 (C2V_108_1056),
	.C2V_17 (C2V_108_1072),
	.C2V_18 (C2V_108_1122),
	.C2V_19 (C2V_108_1259),
	.C2V_20 (C2V_108_1260),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU109 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_23_109),
	.V2C_2 (V2C_59_109),
	.V2C_3 (V2C_127_109),
	.V2C_4 (V2C_188_109),
	.V2C_5 (V2C_202_109),
	.V2C_6 (V2C_245_109),
	.V2C_7 (V2C_345_109),
	.V2C_8 (V2C_399_109),
	.V2C_9 (V2C_496_109),
	.V2C_10 (V2C_732_109),
	.V2C_11 (V2C_780_109),
	.V2C_12 (V2C_828_109),
	.V2C_13 (V2C_869_109),
	.V2C_14 (V2C_958_109),
	.V2C_15 (V2C_992_109),
	.V2C_16 (V2C_1031_109),
	.V2C_17 (V2C_1057_109),
	.V2C_18 (V2C_1116_109),
	.V2C_19 (V2C_1260_109),
	.V2C_20 (V2C_1261_109),
	.C2V_1 (C2V_109_23),
	.C2V_2 (C2V_109_59),
	.C2V_3 (C2V_109_127),
	.C2V_4 (C2V_109_188),
	.C2V_5 (C2V_109_202),
	.C2V_6 (C2V_109_245),
	.C2V_7 (C2V_109_345),
	.C2V_8 (C2V_109_399),
	.C2V_9 (C2V_109_496),
	.C2V_10 (C2V_109_732),
	.C2V_11 (C2V_109_780),
	.C2V_12 (C2V_109_828),
	.C2V_13 (C2V_109_869),
	.C2V_14 (C2V_109_958),
	.C2V_15 (C2V_109_992),
	.C2V_16 (C2V_109_1031),
	.C2V_17 (C2V_109_1057),
	.C2V_18 (C2V_109_1116),
	.C2V_19 (C2V_109_1260),
	.C2V_20 (C2V_109_1261),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU110 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_32_110),
	.V2C_2 (V2C_81_110),
	.V2C_3 (V2C_137_110),
	.V2C_4 (V2C_185_110),
	.V2C_5 (V2C_214_110),
	.V2C_6 (V2C_283_110),
	.V2C_7 (V2C_334_110),
	.V2C_8 (V2C_393_110),
	.V2C_9 (V2C_482_110),
	.V2C_10 (V2C_642_110),
	.V2C_11 (V2C_703_110),
	.V2C_12 (V2C_823_110),
	.V2C_13 (V2C_865_110),
	.V2C_14 (V2C_928_110),
	.V2C_15 (V2C_1007_110),
	.V2C_16 (V2C_1039_110),
	.V2C_17 (V2C_1058_110),
	.V2C_18 (V2C_1137_110),
	.V2C_19 (V2C_1261_110),
	.V2C_20 (V2C_1262_110),
	.C2V_1 (C2V_110_32),
	.C2V_2 (C2V_110_81),
	.C2V_3 (C2V_110_137),
	.C2V_4 (C2V_110_185),
	.C2V_5 (C2V_110_214),
	.C2V_6 (C2V_110_283),
	.C2V_7 (C2V_110_334),
	.C2V_8 (C2V_110_393),
	.C2V_9 (C2V_110_482),
	.C2V_10 (C2V_110_642),
	.C2V_11 (C2V_110_703),
	.C2V_12 (C2V_110_823),
	.C2V_13 (C2V_110_865),
	.C2V_14 (C2V_110_928),
	.C2V_15 (C2V_110_1007),
	.C2V_16 (C2V_110_1039),
	.C2V_17 (C2V_110_1058),
	.C2V_18 (C2V_110_1137),
	.C2V_19 (C2V_110_1261),
	.C2V_20 (C2V_110_1262),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU111 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_27_111),
	.V2C_2 (V2C_54_111),
	.V2C_3 (V2C_119_111),
	.V2C_4 (V2C_153_111),
	.V2C_5 (V2C_219_111),
	.V2C_6 (V2C_286_111),
	.V2C_7 (V2C_383_111),
	.V2C_8 (V2C_390_111),
	.V2C_9 (V2C_549_111),
	.V2C_10 (V2C_606_111),
	.V2C_11 (V2C_634_111),
	.V2C_12 (V2C_738_111),
	.V2C_13 (V2C_869_111),
	.V2C_14 (V2C_913_111),
	.V2C_15 (V2C_986_111),
	.V2C_16 (V2C_1046_111),
	.V2C_17 (V2C_1076_111),
	.V2C_18 (V2C_1121_111),
	.V2C_19 (V2C_1262_111),
	.V2C_20 (V2C_1263_111),
	.C2V_1 (C2V_111_27),
	.C2V_2 (C2V_111_54),
	.C2V_3 (C2V_111_119),
	.C2V_4 (C2V_111_153),
	.C2V_5 (C2V_111_219),
	.C2V_6 (C2V_111_286),
	.C2V_7 (C2V_111_383),
	.C2V_8 (C2V_111_390),
	.C2V_9 (C2V_111_549),
	.C2V_10 (C2V_111_606),
	.C2V_11 (C2V_111_634),
	.C2V_12 (C2V_111_738),
	.C2V_13 (C2V_111_869),
	.C2V_14 (C2V_111_913),
	.C2V_15 (C2V_111_986),
	.C2V_16 (C2V_111_1046),
	.C2V_17 (C2V_111_1076),
	.C2V_18 (C2V_111_1121),
	.C2V_19 (C2V_111_1262),
	.C2V_20 (C2V_111_1263),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU112 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_46_112),
	.V2C_2 (V2C_57_112),
	.V2C_3 (V2C_144_112),
	.V2C_4 (V2C_152_112),
	.V2C_5 (V2C_217_112),
	.V2C_6 (V2C_271_112),
	.V2C_7 (V2C_447_112),
	.V2C_8 (V2C_487_112),
	.V2C_9 (V2C_571_112),
	.V2C_10 (V2C_585_112),
	.V2C_11 (V2C_658_112),
	.V2C_12 (V2C_704_112),
	.V2C_13 (V2C_873_112),
	.V2C_14 (V2C_945_112),
	.V2C_15 (V2C_981_112),
	.V2C_16 (V2C_1011_112),
	.V2C_17 (V2C_1086_112),
	.V2C_18 (V2C_1150_112),
	.V2C_19 (V2C_1263_112),
	.V2C_20 (V2C_1264_112),
	.C2V_1 (C2V_112_46),
	.C2V_2 (C2V_112_57),
	.C2V_3 (C2V_112_144),
	.C2V_4 (C2V_112_152),
	.C2V_5 (C2V_112_217),
	.C2V_6 (C2V_112_271),
	.C2V_7 (C2V_112_447),
	.C2V_8 (C2V_112_487),
	.C2V_9 (C2V_112_571),
	.C2V_10 (C2V_112_585),
	.C2V_11 (C2V_112_658),
	.C2V_12 (C2V_112_704),
	.C2V_13 (C2V_112_873),
	.C2V_14 (C2V_112_945),
	.C2V_15 (C2V_112_981),
	.C2V_16 (C2V_112_1011),
	.C2V_17 (C2V_112_1086),
	.C2V_18 (C2V_112_1150),
	.C2V_19 (C2V_112_1263),
	.C2V_20 (C2V_112_1264),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU113 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_17_113),
	.V2C_2 (V2C_75_113),
	.V2C_3 (V2C_110_113),
	.V2C_4 (V2C_181_113),
	.V2C_5 (V2C_197_113),
	.V2C_6 (V2C_263_113),
	.V2C_7 (V2C_312_113),
	.V2C_8 (V2C_379_113),
	.V2C_9 (V2C_458_113),
	.V2C_10 (V2C_692_113),
	.V2C_11 (V2C_756_113),
	.V2C_12 (V2C_810_113),
	.V2C_13 (V2C_888_113),
	.V2C_14 (V2C_936_113),
	.V2C_15 (V2C_979_113),
	.V2C_16 (V2C_1031_113),
	.V2C_17 (V2C_1080_113),
	.V2C_18 (V2C_1128_113),
	.V2C_19 (V2C_1264_113),
	.V2C_20 (V2C_1265_113),
	.C2V_1 (C2V_113_17),
	.C2V_2 (C2V_113_75),
	.C2V_3 (C2V_113_110),
	.C2V_4 (C2V_113_181),
	.C2V_5 (C2V_113_197),
	.C2V_6 (C2V_113_263),
	.C2V_7 (C2V_113_312),
	.C2V_8 (C2V_113_379),
	.C2V_9 (C2V_113_458),
	.C2V_10 (C2V_113_692),
	.C2V_11 (C2V_113_756),
	.C2V_12 (C2V_113_810),
	.C2V_13 (C2V_113_888),
	.C2V_14 (C2V_113_936),
	.C2V_15 (C2V_113_979),
	.C2V_16 (C2V_113_1031),
	.C2V_17 (C2V_113_1080),
	.C2V_18 (C2V_113_1128),
	.C2V_19 (C2V_113_1264),
	.C2V_20 (C2V_113_1265),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU114 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_48_114),
	.V2C_2 (V2C_72_114),
	.V2C_3 (V2C_112_114),
	.V2C_4 (V2C_180_114),
	.V2C_5 (V2C_214_114),
	.V2C_6 (V2C_245_114),
	.V2C_7 (V2C_298_114),
	.V2C_8 (V2C_450_114),
	.V2C_9 (V2C_547_114),
	.V2C_10 (V2C_580_114),
	.V2C_11 (V2C_784_114),
	.V2C_12 (V2C_860_114),
	.V2C_13 (V2C_893_114),
	.V2C_14 (V2C_955_114),
	.V2C_15 (V2C_990_114),
	.V2C_16 (V2C_1009_114),
	.V2C_17 (V2C_1073_114),
	.V2C_18 (V2C_1123_114),
	.V2C_19 (V2C_1265_114),
	.V2C_20 (V2C_1266_114),
	.C2V_1 (C2V_114_48),
	.C2V_2 (C2V_114_72),
	.C2V_3 (C2V_114_112),
	.C2V_4 (C2V_114_180),
	.C2V_5 (C2V_114_214),
	.C2V_6 (C2V_114_245),
	.C2V_7 (C2V_114_298),
	.C2V_8 (C2V_114_450),
	.C2V_9 (C2V_114_547),
	.C2V_10 (C2V_114_580),
	.C2V_11 (C2V_114_784),
	.C2V_12 (C2V_114_860),
	.C2V_13 (C2V_114_893),
	.C2V_14 (C2V_114_955),
	.C2V_15 (C2V_114_990),
	.C2V_16 (C2V_114_1009),
	.C2V_17 (C2V_114_1073),
	.C2V_18 (C2V_114_1123),
	.C2V_19 (C2V_114_1265),
	.C2V_20 (C2V_114_1266),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU115 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_24_115),
	.V2C_2 (V2C_60_115),
	.V2C_3 (V2C_128_115),
	.V2C_4 (V2C_189_115),
	.V2C_5 (V2C_203_115),
	.V2C_6 (V2C_246_115),
	.V2C_7 (V2C_346_115),
	.V2C_8 (V2C_400_115),
	.V2C_9 (V2C_497_115),
	.V2C_10 (V2C_733_115),
	.V2C_11 (V2C_781_115),
	.V2C_12 (V2C_829_115),
	.V2C_13 (V2C_870_115),
	.V2C_14 (V2C_959_115),
	.V2C_15 (V2C_993_115),
	.V2C_16 (V2C_1032_115),
	.V2C_17 (V2C_1058_115),
	.V2C_18 (V2C_1117_115),
	.V2C_19 (V2C_1266_115),
	.V2C_20 (V2C_1267_115),
	.C2V_1 (C2V_115_24),
	.C2V_2 (C2V_115_60),
	.C2V_3 (C2V_115_128),
	.C2V_4 (C2V_115_189),
	.C2V_5 (C2V_115_203),
	.C2V_6 (C2V_115_246),
	.C2V_7 (C2V_115_346),
	.C2V_8 (C2V_115_400),
	.C2V_9 (C2V_115_497),
	.C2V_10 (C2V_115_733),
	.C2V_11 (C2V_115_781),
	.C2V_12 (C2V_115_829),
	.C2V_13 (C2V_115_870),
	.C2V_14 (C2V_115_959),
	.C2V_15 (C2V_115_993),
	.C2V_16 (C2V_115_1032),
	.C2V_17 (C2V_115_1058),
	.C2V_18 (C2V_115_1117),
	.C2V_19 (C2V_115_1266),
	.C2V_20 (C2V_115_1267),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU116 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_33_116),
	.V2C_2 (V2C_82_116),
	.V2C_3 (V2C_138_116),
	.V2C_4 (V2C_186_116),
	.V2C_5 (V2C_215_116),
	.V2C_6 (V2C_284_116),
	.V2C_7 (V2C_335_116),
	.V2C_8 (V2C_394_116),
	.V2C_9 (V2C_483_116),
	.V2C_10 (V2C_643_116),
	.V2C_11 (V2C_704_116),
	.V2C_12 (V2C_824_116),
	.V2C_13 (V2C_866_116),
	.V2C_14 (V2C_929_116),
	.V2C_15 (V2C_1008_116),
	.V2C_16 (V2C_1040_116),
	.V2C_17 (V2C_1059_116),
	.V2C_18 (V2C_1138_116),
	.V2C_19 (V2C_1267_116),
	.V2C_20 (V2C_1268_116),
	.C2V_1 (C2V_116_33),
	.C2V_2 (C2V_116_82),
	.C2V_3 (C2V_116_138),
	.C2V_4 (C2V_116_186),
	.C2V_5 (C2V_116_215),
	.C2V_6 (C2V_116_284),
	.C2V_7 (C2V_116_335),
	.C2V_8 (C2V_116_394),
	.C2V_9 (C2V_116_483),
	.C2V_10 (C2V_116_643),
	.C2V_11 (C2V_116_704),
	.C2V_12 (C2V_116_824),
	.C2V_13 (C2V_116_866),
	.C2V_14 (C2V_116_929),
	.C2V_15 (C2V_116_1008),
	.C2V_16 (C2V_116_1040),
	.C2V_17 (C2V_116_1059),
	.C2V_18 (C2V_116_1138),
	.C2V_19 (C2V_116_1267),
	.C2V_20 (C2V_116_1268),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU117 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_28_117),
	.V2C_2 (V2C_55_117),
	.V2C_3 (V2C_120_117),
	.V2C_4 (V2C_154_117),
	.V2C_5 (V2C_220_117),
	.V2C_6 (V2C_287_117),
	.V2C_7 (V2C_384_117),
	.V2C_8 (V2C_391_117),
	.V2C_9 (V2C_550_117),
	.V2C_10 (V2C_607_117),
	.V2C_11 (V2C_635_117),
	.V2C_12 (V2C_739_117),
	.V2C_13 (V2C_870_117),
	.V2C_14 (V2C_914_117),
	.V2C_15 (V2C_987_117),
	.V2C_16 (V2C_1047_117),
	.V2C_17 (V2C_1077_117),
	.V2C_18 (V2C_1122_117),
	.V2C_19 (V2C_1268_117),
	.V2C_20 (V2C_1269_117),
	.C2V_1 (C2V_117_28),
	.C2V_2 (C2V_117_55),
	.C2V_3 (C2V_117_120),
	.C2V_4 (C2V_117_154),
	.C2V_5 (C2V_117_220),
	.C2V_6 (C2V_117_287),
	.C2V_7 (C2V_117_384),
	.C2V_8 (C2V_117_391),
	.C2V_9 (C2V_117_550),
	.C2V_10 (C2V_117_607),
	.C2V_11 (C2V_117_635),
	.C2V_12 (C2V_117_739),
	.C2V_13 (C2V_117_870),
	.C2V_14 (C2V_117_914),
	.C2V_15 (C2V_117_987),
	.C2V_16 (C2V_117_1047),
	.C2V_17 (C2V_117_1077),
	.C2V_18 (C2V_117_1122),
	.C2V_19 (C2V_117_1268),
	.C2V_20 (C2V_117_1269),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU118 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_47_118),
	.V2C_2 (V2C_58_118),
	.V2C_3 (V2C_97_118),
	.V2C_4 (V2C_153_118),
	.V2C_5 (V2C_218_118),
	.V2C_6 (V2C_272_118),
	.V2C_7 (V2C_448_118),
	.V2C_8 (V2C_488_118),
	.V2C_9 (V2C_572_118),
	.V2C_10 (V2C_586_118),
	.V2C_11 (V2C_659_118),
	.V2C_12 (V2C_705_118),
	.V2C_13 (V2C_874_118),
	.V2C_14 (V2C_946_118),
	.V2C_15 (V2C_982_118),
	.V2C_16 (V2C_1012_118),
	.V2C_17 (V2C_1087_118),
	.V2C_18 (V2C_1151_118),
	.V2C_19 (V2C_1269_118),
	.V2C_20 (V2C_1270_118),
	.C2V_1 (C2V_118_47),
	.C2V_2 (C2V_118_58),
	.C2V_3 (C2V_118_97),
	.C2V_4 (C2V_118_153),
	.C2V_5 (C2V_118_218),
	.C2V_6 (C2V_118_272),
	.C2V_7 (C2V_118_448),
	.C2V_8 (C2V_118_488),
	.C2V_9 (C2V_118_572),
	.C2V_10 (C2V_118_586),
	.C2V_11 (C2V_118_659),
	.C2V_12 (C2V_118_705),
	.C2V_13 (C2V_118_874),
	.C2V_14 (C2V_118_946),
	.C2V_15 (C2V_118_982),
	.C2V_16 (C2V_118_1012),
	.C2V_17 (C2V_118_1087),
	.C2V_18 (C2V_118_1151),
	.C2V_19 (C2V_118_1269),
	.C2V_20 (C2V_118_1270),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU119 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_18_119),
	.V2C_2 (V2C_76_119),
	.V2C_3 (V2C_111_119),
	.V2C_4 (V2C_182_119),
	.V2C_5 (V2C_198_119),
	.V2C_6 (V2C_264_119),
	.V2C_7 (V2C_313_119),
	.V2C_8 (V2C_380_119),
	.V2C_9 (V2C_459_119),
	.V2C_10 (V2C_693_119),
	.V2C_11 (V2C_757_119),
	.V2C_12 (V2C_811_119),
	.V2C_13 (V2C_889_119),
	.V2C_14 (V2C_937_119),
	.V2C_15 (V2C_980_119),
	.V2C_16 (V2C_1032_119),
	.V2C_17 (V2C_1081_119),
	.V2C_18 (V2C_1129_119),
	.V2C_19 (V2C_1270_119),
	.V2C_20 (V2C_1271_119),
	.C2V_1 (C2V_119_18),
	.C2V_2 (C2V_119_76),
	.C2V_3 (C2V_119_111),
	.C2V_4 (C2V_119_182),
	.C2V_5 (C2V_119_198),
	.C2V_6 (C2V_119_264),
	.C2V_7 (C2V_119_313),
	.C2V_8 (C2V_119_380),
	.C2V_9 (C2V_119_459),
	.C2V_10 (C2V_119_693),
	.C2V_11 (C2V_119_757),
	.C2V_12 (C2V_119_811),
	.C2V_13 (C2V_119_889),
	.C2V_14 (C2V_119_937),
	.C2V_15 (C2V_119_980),
	.C2V_16 (C2V_119_1032),
	.C2V_17 (C2V_119_1081),
	.C2V_18 (C2V_119_1129),
	.C2V_19 (C2V_119_1270),
	.C2V_20 (C2V_119_1271),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU120 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_1_120),
	.V2C_2 (V2C_73_120),
	.V2C_3 (V2C_113_120),
	.V2C_4 (V2C_181_120),
	.V2C_5 (V2C_215_120),
	.V2C_6 (V2C_246_120),
	.V2C_7 (V2C_299_120),
	.V2C_8 (V2C_451_120),
	.V2C_9 (V2C_548_120),
	.V2C_10 (V2C_581_120),
	.V2C_11 (V2C_785_120),
	.V2C_12 (V2C_861_120),
	.V2C_13 (V2C_894_120),
	.V2C_14 (V2C_956_120),
	.V2C_15 (V2C_991_120),
	.V2C_16 (V2C_1010_120),
	.V2C_17 (V2C_1074_120),
	.V2C_18 (V2C_1124_120),
	.V2C_19 (V2C_1271_120),
	.V2C_20 (V2C_1272_120),
	.C2V_1 (C2V_120_1),
	.C2V_2 (C2V_120_73),
	.C2V_3 (C2V_120_113),
	.C2V_4 (C2V_120_181),
	.C2V_5 (C2V_120_215),
	.C2V_6 (C2V_120_246),
	.C2V_7 (C2V_120_299),
	.C2V_8 (C2V_120_451),
	.C2V_9 (C2V_120_548),
	.C2V_10 (C2V_120_581),
	.C2V_11 (C2V_120_785),
	.C2V_12 (C2V_120_861),
	.C2V_13 (C2V_120_894),
	.C2V_14 (C2V_120_956),
	.C2V_15 (C2V_120_991),
	.C2V_16 (C2V_120_1010),
	.C2V_17 (C2V_120_1074),
	.C2V_18 (C2V_120_1124),
	.C2V_19 (C2V_120_1271),
	.C2V_20 (C2V_120_1272),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU121 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_25_121),
	.V2C_2 (V2C_61_121),
	.V2C_3 (V2C_129_121),
	.V2C_4 (V2C_190_121),
	.V2C_5 (V2C_204_121),
	.V2C_6 (V2C_247_121),
	.V2C_7 (V2C_347_121),
	.V2C_8 (V2C_401_121),
	.V2C_9 (V2C_498_121),
	.V2C_10 (V2C_734_121),
	.V2C_11 (V2C_782_121),
	.V2C_12 (V2C_830_121),
	.V2C_13 (V2C_871_121),
	.V2C_14 (V2C_960_121),
	.V2C_15 (V2C_994_121),
	.V2C_16 (V2C_1033_121),
	.V2C_17 (V2C_1059_121),
	.V2C_18 (V2C_1118_121),
	.V2C_19 (V2C_1272_121),
	.V2C_20 (V2C_1273_121),
	.C2V_1 (C2V_121_25),
	.C2V_2 (C2V_121_61),
	.C2V_3 (C2V_121_129),
	.C2V_4 (C2V_121_190),
	.C2V_5 (C2V_121_204),
	.C2V_6 (C2V_121_247),
	.C2V_7 (C2V_121_347),
	.C2V_8 (C2V_121_401),
	.C2V_9 (C2V_121_498),
	.C2V_10 (C2V_121_734),
	.C2V_11 (C2V_121_782),
	.C2V_12 (C2V_121_830),
	.C2V_13 (C2V_121_871),
	.C2V_14 (C2V_121_960),
	.C2V_15 (C2V_121_994),
	.C2V_16 (C2V_121_1033),
	.C2V_17 (C2V_121_1059),
	.C2V_18 (C2V_121_1118),
	.C2V_19 (C2V_121_1272),
	.C2V_20 (C2V_121_1273),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU122 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_34_122),
	.V2C_2 (V2C_83_122),
	.V2C_3 (V2C_139_122),
	.V2C_4 (V2C_187_122),
	.V2C_5 (V2C_216_122),
	.V2C_6 (V2C_285_122),
	.V2C_7 (V2C_336_122),
	.V2C_8 (V2C_395_122),
	.V2C_9 (V2C_484_122),
	.V2C_10 (V2C_644_122),
	.V2C_11 (V2C_705_122),
	.V2C_12 (V2C_825_122),
	.V2C_13 (V2C_867_122),
	.V2C_14 (V2C_930_122),
	.V2C_15 (V2C_961_122),
	.V2C_16 (V2C_1041_122),
	.V2C_17 (V2C_1060_122),
	.V2C_18 (V2C_1139_122),
	.V2C_19 (V2C_1273_122),
	.V2C_20 (V2C_1274_122),
	.C2V_1 (C2V_122_34),
	.C2V_2 (C2V_122_83),
	.C2V_3 (C2V_122_139),
	.C2V_4 (C2V_122_187),
	.C2V_5 (C2V_122_216),
	.C2V_6 (C2V_122_285),
	.C2V_7 (C2V_122_336),
	.C2V_8 (C2V_122_395),
	.C2V_9 (C2V_122_484),
	.C2V_10 (C2V_122_644),
	.C2V_11 (C2V_122_705),
	.C2V_12 (C2V_122_825),
	.C2V_13 (C2V_122_867),
	.C2V_14 (C2V_122_930),
	.C2V_15 (C2V_122_961),
	.C2V_16 (C2V_122_1041),
	.C2V_17 (C2V_122_1060),
	.C2V_18 (C2V_122_1139),
	.C2V_19 (C2V_122_1273),
	.C2V_20 (C2V_122_1274),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU123 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_29_123),
	.V2C_2 (V2C_56_123),
	.V2C_3 (V2C_121_123),
	.V2C_4 (V2C_155_123),
	.V2C_5 (V2C_221_123),
	.V2C_6 (V2C_288_123),
	.V2C_7 (V2C_337_123),
	.V2C_8 (V2C_392_123),
	.V2C_9 (V2C_551_123),
	.V2C_10 (V2C_608_123),
	.V2C_11 (V2C_636_123),
	.V2C_12 (V2C_740_123),
	.V2C_13 (V2C_871_123),
	.V2C_14 (V2C_915_123),
	.V2C_15 (V2C_988_123),
	.V2C_16 (V2C_1048_123),
	.V2C_17 (V2C_1078_123),
	.V2C_18 (V2C_1123_123),
	.V2C_19 (V2C_1274_123),
	.V2C_20 (V2C_1275_123),
	.C2V_1 (C2V_123_29),
	.C2V_2 (C2V_123_56),
	.C2V_3 (C2V_123_121),
	.C2V_4 (C2V_123_155),
	.C2V_5 (C2V_123_221),
	.C2V_6 (C2V_123_288),
	.C2V_7 (C2V_123_337),
	.C2V_8 (C2V_123_392),
	.C2V_9 (C2V_123_551),
	.C2V_10 (C2V_123_608),
	.C2V_11 (C2V_123_636),
	.C2V_12 (C2V_123_740),
	.C2V_13 (C2V_123_871),
	.C2V_14 (C2V_123_915),
	.C2V_15 (C2V_123_988),
	.C2V_16 (C2V_123_1048),
	.C2V_17 (C2V_123_1078),
	.C2V_18 (C2V_123_1123),
	.C2V_19 (C2V_123_1274),
	.C2V_20 (C2V_123_1275),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU124 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_48_124),
	.V2C_2 (V2C_59_124),
	.V2C_3 (V2C_98_124),
	.V2C_4 (V2C_154_124),
	.V2C_5 (V2C_219_124),
	.V2C_6 (V2C_273_124),
	.V2C_7 (V2C_449_124),
	.V2C_8 (V2C_489_124),
	.V2C_9 (V2C_573_124),
	.V2C_10 (V2C_587_124),
	.V2C_11 (V2C_660_124),
	.V2C_12 (V2C_706_124),
	.V2C_13 (V2C_875_124),
	.V2C_14 (V2C_947_124),
	.V2C_15 (V2C_983_124),
	.V2C_16 (V2C_1013_124),
	.V2C_17 (V2C_1088_124),
	.V2C_18 (V2C_1152_124),
	.V2C_19 (V2C_1275_124),
	.V2C_20 (V2C_1276_124),
	.C2V_1 (C2V_124_48),
	.C2V_2 (C2V_124_59),
	.C2V_3 (C2V_124_98),
	.C2V_4 (C2V_124_154),
	.C2V_5 (C2V_124_219),
	.C2V_6 (C2V_124_273),
	.C2V_7 (C2V_124_449),
	.C2V_8 (C2V_124_489),
	.C2V_9 (C2V_124_573),
	.C2V_10 (C2V_124_587),
	.C2V_11 (C2V_124_660),
	.C2V_12 (C2V_124_706),
	.C2V_13 (C2V_124_875),
	.C2V_14 (C2V_124_947),
	.C2V_15 (C2V_124_983),
	.C2V_16 (C2V_124_1013),
	.C2V_17 (C2V_124_1088),
	.C2V_18 (C2V_124_1152),
	.C2V_19 (C2V_124_1275),
	.C2V_20 (C2V_124_1276),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU125 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_19_125),
	.V2C_2 (V2C_77_125),
	.V2C_3 (V2C_112_125),
	.V2C_4 (V2C_183_125),
	.V2C_5 (V2C_199_125),
	.V2C_6 (V2C_265_125),
	.V2C_7 (V2C_314_125),
	.V2C_8 (V2C_381_125),
	.V2C_9 (V2C_460_125),
	.V2C_10 (V2C_694_125),
	.V2C_11 (V2C_758_125),
	.V2C_12 (V2C_812_125),
	.V2C_13 (V2C_890_125),
	.V2C_14 (V2C_938_125),
	.V2C_15 (V2C_981_125),
	.V2C_16 (V2C_1033_125),
	.V2C_17 (V2C_1082_125),
	.V2C_18 (V2C_1130_125),
	.V2C_19 (V2C_1276_125),
	.V2C_20 (V2C_1277_125),
	.C2V_1 (C2V_125_19),
	.C2V_2 (C2V_125_77),
	.C2V_3 (C2V_125_112),
	.C2V_4 (C2V_125_183),
	.C2V_5 (C2V_125_199),
	.C2V_6 (C2V_125_265),
	.C2V_7 (C2V_125_314),
	.C2V_8 (C2V_125_381),
	.C2V_9 (C2V_125_460),
	.C2V_10 (C2V_125_694),
	.C2V_11 (C2V_125_758),
	.C2V_12 (C2V_125_812),
	.C2V_13 (C2V_125_890),
	.C2V_14 (C2V_125_938),
	.C2V_15 (C2V_125_981),
	.C2V_16 (C2V_125_1033),
	.C2V_17 (C2V_125_1082),
	.C2V_18 (C2V_125_1130),
	.C2V_19 (C2V_125_1276),
	.C2V_20 (C2V_125_1277),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU126 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_2_126),
	.V2C_2 (V2C_74_126),
	.V2C_3 (V2C_114_126),
	.V2C_4 (V2C_182_126),
	.V2C_5 (V2C_216_126),
	.V2C_6 (V2C_247_126),
	.V2C_7 (V2C_300_126),
	.V2C_8 (V2C_452_126),
	.V2C_9 (V2C_549_126),
	.V2C_10 (V2C_582_126),
	.V2C_11 (V2C_786_126),
	.V2C_12 (V2C_862_126),
	.V2C_13 (V2C_895_126),
	.V2C_14 (V2C_957_126),
	.V2C_15 (V2C_992_126),
	.V2C_16 (V2C_1011_126),
	.V2C_17 (V2C_1075_126),
	.V2C_18 (V2C_1125_126),
	.V2C_19 (V2C_1277_126),
	.V2C_20 (V2C_1278_126),
	.C2V_1 (C2V_126_2),
	.C2V_2 (C2V_126_74),
	.C2V_3 (C2V_126_114),
	.C2V_4 (C2V_126_182),
	.C2V_5 (C2V_126_216),
	.C2V_6 (C2V_126_247),
	.C2V_7 (C2V_126_300),
	.C2V_8 (C2V_126_452),
	.C2V_9 (C2V_126_549),
	.C2V_10 (C2V_126_582),
	.C2V_11 (C2V_126_786),
	.C2V_12 (C2V_126_862),
	.C2V_13 (C2V_126_895),
	.C2V_14 (C2V_126_957),
	.C2V_15 (C2V_126_992),
	.C2V_16 (C2V_126_1011),
	.C2V_17 (C2V_126_1075),
	.C2V_18 (C2V_126_1125),
	.C2V_19 (C2V_126_1277),
	.C2V_20 (C2V_126_1278),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU127 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_26_127),
	.V2C_2 (V2C_62_127),
	.V2C_3 (V2C_130_127),
	.V2C_4 (V2C_191_127),
	.V2C_5 (V2C_205_127),
	.V2C_6 (V2C_248_127),
	.V2C_7 (V2C_348_127),
	.V2C_8 (V2C_402_127),
	.V2C_9 (V2C_499_127),
	.V2C_10 (V2C_735_127),
	.V2C_11 (V2C_783_127),
	.V2C_12 (V2C_831_127),
	.V2C_13 (V2C_872_127),
	.V2C_14 (V2C_913_127),
	.V2C_15 (V2C_995_127),
	.V2C_16 (V2C_1034_127),
	.V2C_17 (V2C_1060_127),
	.V2C_18 (V2C_1119_127),
	.V2C_19 (V2C_1278_127),
	.V2C_20 (V2C_1279_127),
	.C2V_1 (C2V_127_26),
	.C2V_2 (C2V_127_62),
	.C2V_3 (C2V_127_130),
	.C2V_4 (C2V_127_191),
	.C2V_5 (C2V_127_205),
	.C2V_6 (C2V_127_248),
	.C2V_7 (C2V_127_348),
	.C2V_8 (C2V_127_402),
	.C2V_9 (C2V_127_499),
	.C2V_10 (C2V_127_735),
	.C2V_11 (C2V_127_783),
	.C2V_12 (C2V_127_831),
	.C2V_13 (C2V_127_872),
	.C2V_14 (C2V_127_913),
	.C2V_15 (C2V_127_995),
	.C2V_16 (C2V_127_1034),
	.C2V_17 (C2V_127_1060),
	.C2V_18 (C2V_127_1119),
	.C2V_19 (C2V_127_1278),
	.C2V_20 (C2V_127_1279),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU128 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_35_128),
	.V2C_2 (V2C_84_128),
	.V2C_3 (V2C_140_128),
	.V2C_4 (V2C_188_128),
	.V2C_5 (V2C_217_128),
	.V2C_6 (V2C_286_128),
	.V2C_7 (V2C_289_128),
	.V2C_8 (V2C_396_128),
	.V2C_9 (V2C_485_128),
	.V2C_10 (V2C_645_128),
	.V2C_11 (V2C_706_128),
	.V2C_12 (V2C_826_128),
	.V2C_13 (V2C_868_128),
	.V2C_14 (V2C_931_128),
	.V2C_15 (V2C_962_128),
	.V2C_16 (V2C_1042_128),
	.V2C_17 (V2C_1061_128),
	.V2C_18 (V2C_1140_128),
	.V2C_19 (V2C_1279_128),
	.V2C_20 (V2C_1280_128),
	.C2V_1 (C2V_128_35),
	.C2V_2 (C2V_128_84),
	.C2V_3 (C2V_128_140),
	.C2V_4 (C2V_128_188),
	.C2V_5 (C2V_128_217),
	.C2V_6 (C2V_128_286),
	.C2V_7 (C2V_128_289),
	.C2V_8 (C2V_128_396),
	.C2V_9 (C2V_128_485),
	.C2V_10 (C2V_128_645),
	.C2V_11 (C2V_128_706),
	.C2V_12 (C2V_128_826),
	.C2V_13 (C2V_128_868),
	.C2V_14 (C2V_128_931),
	.C2V_15 (C2V_128_962),
	.C2V_16 (C2V_128_1042),
	.C2V_17 (C2V_128_1061),
	.C2V_18 (C2V_128_1140),
	.C2V_19 (C2V_128_1279),
	.C2V_20 (C2V_128_1280),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU129 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_30_129),
	.V2C_2 (V2C_57_129),
	.V2C_3 (V2C_122_129),
	.V2C_4 (V2C_156_129),
	.V2C_5 (V2C_222_129),
	.V2C_6 (V2C_241_129),
	.V2C_7 (V2C_338_129),
	.V2C_8 (V2C_393_129),
	.V2C_9 (V2C_552_129),
	.V2C_10 (V2C_609_129),
	.V2C_11 (V2C_637_129),
	.V2C_12 (V2C_741_129),
	.V2C_13 (V2C_872_129),
	.V2C_14 (V2C_916_129),
	.V2C_15 (V2C_989_129),
	.V2C_16 (V2C_1049_129),
	.V2C_17 (V2C_1079_129),
	.V2C_18 (V2C_1124_129),
	.V2C_19 (V2C_1280_129),
	.V2C_20 (V2C_1281_129),
	.C2V_1 (C2V_129_30),
	.C2V_2 (C2V_129_57),
	.C2V_3 (C2V_129_122),
	.C2V_4 (C2V_129_156),
	.C2V_5 (C2V_129_222),
	.C2V_6 (C2V_129_241),
	.C2V_7 (C2V_129_338),
	.C2V_8 (C2V_129_393),
	.C2V_9 (C2V_129_552),
	.C2V_10 (C2V_129_609),
	.C2V_11 (C2V_129_637),
	.C2V_12 (C2V_129_741),
	.C2V_13 (C2V_129_872),
	.C2V_14 (C2V_129_916),
	.C2V_15 (C2V_129_989),
	.C2V_16 (C2V_129_1049),
	.C2V_17 (C2V_129_1079),
	.C2V_18 (C2V_129_1124),
	.C2V_19 (C2V_129_1280),
	.C2V_20 (C2V_129_1281),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU130 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_1_130),
	.V2C_2 (V2C_60_130),
	.V2C_3 (V2C_99_130),
	.V2C_4 (V2C_155_130),
	.V2C_5 (V2C_220_130),
	.V2C_6 (V2C_274_130),
	.V2C_7 (V2C_450_130),
	.V2C_8 (V2C_490_130),
	.V2C_9 (V2C_574_130),
	.V2C_10 (V2C_588_130),
	.V2C_11 (V2C_661_130),
	.V2C_12 (V2C_707_130),
	.V2C_13 (V2C_876_130),
	.V2C_14 (V2C_948_130),
	.V2C_15 (V2C_984_130),
	.V2C_16 (V2C_1014_130),
	.V2C_17 (V2C_1089_130),
	.V2C_18 (V2C_1105_130),
	.V2C_19 (V2C_1281_130),
	.V2C_20 (V2C_1282_130),
	.C2V_1 (C2V_130_1),
	.C2V_2 (C2V_130_60),
	.C2V_3 (C2V_130_99),
	.C2V_4 (C2V_130_155),
	.C2V_5 (C2V_130_220),
	.C2V_6 (C2V_130_274),
	.C2V_7 (C2V_130_450),
	.C2V_8 (C2V_130_490),
	.C2V_9 (C2V_130_574),
	.C2V_10 (C2V_130_588),
	.C2V_11 (C2V_130_661),
	.C2V_12 (C2V_130_707),
	.C2V_13 (C2V_130_876),
	.C2V_14 (C2V_130_948),
	.C2V_15 (C2V_130_984),
	.C2V_16 (C2V_130_1014),
	.C2V_17 (C2V_130_1089),
	.C2V_18 (C2V_130_1105),
	.C2V_19 (C2V_130_1281),
	.C2V_20 (C2V_130_1282),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU131 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_20_131),
	.V2C_2 (V2C_78_131),
	.V2C_3 (V2C_113_131),
	.V2C_4 (V2C_184_131),
	.V2C_5 (V2C_200_131),
	.V2C_6 (V2C_266_131),
	.V2C_7 (V2C_315_131),
	.V2C_8 (V2C_382_131),
	.V2C_9 (V2C_461_131),
	.V2C_10 (V2C_695_131),
	.V2C_11 (V2C_759_131),
	.V2C_12 (V2C_813_131),
	.V2C_13 (V2C_891_131),
	.V2C_14 (V2C_939_131),
	.V2C_15 (V2C_982_131),
	.V2C_16 (V2C_1034_131),
	.V2C_17 (V2C_1083_131),
	.V2C_18 (V2C_1131_131),
	.V2C_19 (V2C_1282_131),
	.V2C_20 (V2C_1283_131),
	.C2V_1 (C2V_131_20),
	.C2V_2 (C2V_131_78),
	.C2V_3 (C2V_131_113),
	.C2V_4 (C2V_131_184),
	.C2V_5 (C2V_131_200),
	.C2V_6 (C2V_131_266),
	.C2V_7 (C2V_131_315),
	.C2V_8 (C2V_131_382),
	.C2V_9 (C2V_131_461),
	.C2V_10 (C2V_131_695),
	.C2V_11 (C2V_131_759),
	.C2V_12 (C2V_131_813),
	.C2V_13 (C2V_131_891),
	.C2V_14 (C2V_131_939),
	.C2V_15 (C2V_131_982),
	.C2V_16 (C2V_131_1034),
	.C2V_17 (C2V_131_1083),
	.C2V_18 (C2V_131_1131),
	.C2V_19 (C2V_131_1282),
	.C2V_20 (C2V_131_1283),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU132 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_3_132),
	.V2C_2 (V2C_75_132),
	.V2C_3 (V2C_115_132),
	.V2C_4 (V2C_183_132),
	.V2C_5 (V2C_217_132),
	.V2C_6 (V2C_248_132),
	.V2C_7 (V2C_301_132),
	.V2C_8 (V2C_453_132),
	.V2C_9 (V2C_550_132),
	.V2C_10 (V2C_583_132),
	.V2C_11 (V2C_787_132),
	.V2C_12 (V2C_863_132),
	.V2C_13 (V2C_896_132),
	.V2C_14 (V2C_958_132),
	.V2C_15 (V2C_993_132),
	.V2C_16 (V2C_1012_132),
	.V2C_17 (V2C_1076_132),
	.V2C_18 (V2C_1126_132),
	.V2C_19 (V2C_1283_132),
	.V2C_20 (V2C_1284_132),
	.C2V_1 (C2V_132_3),
	.C2V_2 (C2V_132_75),
	.C2V_3 (C2V_132_115),
	.C2V_4 (C2V_132_183),
	.C2V_5 (C2V_132_217),
	.C2V_6 (C2V_132_248),
	.C2V_7 (C2V_132_301),
	.C2V_8 (C2V_132_453),
	.C2V_9 (C2V_132_550),
	.C2V_10 (C2V_132_583),
	.C2V_11 (C2V_132_787),
	.C2V_12 (C2V_132_863),
	.C2V_13 (C2V_132_896),
	.C2V_14 (C2V_132_958),
	.C2V_15 (C2V_132_993),
	.C2V_16 (C2V_132_1012),
	.C2V_17 (C2V_132_1076),
	.C2V_18 (C2V_132_1126),
	.C2V_19 (C2V_132_1283),
	.C2V_20 (C2V_132_1284),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU133 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_27_133),
	.V2C_2 (V2C_63_133),
	.V2C_3 (V2C_131_133),
	.V2C_4 (V2C_192_133),
	.V2C_5 (V2C_206_133),
	.V2C_6 (V2C_249_133),
	.V2C_7 (V2C_349_133),
	.V2C_8 (V2C_403_133),
	.V2C_9 (V2C_500_133),
	.V2C_10 (V2C_736_133),
	.V2C_11 (V2C_784_133),
	.V2C_12 (V2C_832_133),
	.V2C_13 (V2C_873_133),
	.V2C_14 (V2C_914_133),
	.V2C_15 (V2C_996_133),
	.V2C_16 (V2C_1035_133),
	.V2C_17 (V2C_1061_133),
	.V2C_18 (V2C_1120_133),
	.V2C_19 (V2C_1284_133),
	.V2C_20 (V2C_1285_133),
	.C2V_1 (C2V_133_27),
	.C2V_2 (C2V_133_63),
	.C2V_3 (C2V_133_131),
	.C2V_4 (C2V_133_192),
	.C2V_5 (C2V_133_206),
	.C2V_6 (C2V_133_249),
	.C2V_7 (C2V_133_349),
	.C2V_8 (C2V_133_403),
	.C2V_9 (C2V_133_500),
	.C2V_10 (C2V_133_736),
	.C2V_11 (C2V_133_784),
	.C2V_12 (C2V_133_832),
	.C2V_13 (C2V_133_873),
	.C2V_14 (C2V_133_914),
	.C2V_15 (C2V_133_996),
	.C2V_16 (C2V_133_1035),
	.C2V_17 (C2V_133_1061),
	.C2V_18 (C2V_133_1120),
	.C2V_19 (C2V_133_1284),
	.C2V_20 (C2V_133_1285),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU134 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_36_134),
	.V2C_2 (V2C_85_134),
	.V2C_3 (V2C_141_134),
	.V2C_4 (V2C_189_134),
	.V2C_5 (V2C_218_134),
	.V2C_6 (V2C_287_134),
	.V2C_7 (V2C_290_134),
	.V2C_8 (V2C_397_134),
	.V2C_9 (V2C_486_134),
	.V2C_10 (V2C_646_134),
	.V2C_11 (V2C_707_134),
	.V2C_12 (V2C_827_134),
	.V2C_13 (V2C_869_134),
	.V2C_14 (V2C_932_134),
	.V2C_15 (V2C_963_134),
	.V2C_16 (V2C_1043_134),
	.V2C_17 (V2C_1062_134),
	.V2C_18 (V2C_1141_134),
	.V2C_19 (V2C_1285_134),
	.V2C_20 (V2C_1286_134),
	.C2V_1 (C2V_134_36),
	.C2V_2 (C2V_134_85),
	.C2V_3 (C2V_134_141),
	.C2V_4 (C2V_134_189),
	.C2V_5 (C2V_134_218),
	.C2V_6 (C2V_134_287),
	.C2V_7 (C2V_134_290),
	.C2V_8 (C2V_134_397),
	.C2V_9 (C2V_134_486),
	.C2V_10 (C2V_134_646),
	.C2V_11 (C2V_134_707),
	.C2V_12 (C2V_134_827),
	.C2V_13 (C2V_134_869),
	.C2V_14 (C2V_134_932),
	.C2V_15 (C2V_134_963),
	.C2V_16 (C2V_134_1043),
	.C2V_17 (C2V_134_1062),
	.C2V_18 (C2V_134_1141),
	.C2V_19 (C2V_134_1285),
	.C2V_20 (C2V_134_1286),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU135 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_31_135),
	.V2C_2 (V2C_58_135),
	.V2C_3 (V2C_123_135),
	.V2C_4 (V2C_157_135),
	.V2C_5 (V2C_223_135),
	.V2C_6 (V2C_242_135),
	.V2C_7 (V2C_339_135),
	.V2C_8 (V2C_394_135),
	.V2C_9 (V2C_553_135),
	.V2C_10 (V2C_610_135),
	.V2C_11 (V2C_638_135),
	.V2C_12 (V2C_742_135),
	.V2C_13 (V2C_873_135),
	.V2C_14 (V2C_917_135),
	.V2C_15 (V2C_990_135),
	.V2C_16 (V2C_1050_135),
	.V2C_17 (V2C_1080_135),
	.V2C_18 (V2C_1125_135),
	.V2C_19 (V2C_1286_135),
	.V2C_20 (V2C_1287_135),
	.C2V_1 (C2V_135_31),
	.C2V_2 (C2V_135_58),
	.C2V_3 (C2V_135_123),
	.C2V_4 (C2V_135_157),
	.C2V_5 (C2V_135_223),
	.C2V_6 (C2V_135_242),
	.C2V_7 (C2V_135_339),
	.C2V_8 (C2V_135_394),
	.C2V_9 (C2V_135_553),
	.C2V_10 (C2V_135_610),
	.C2V_11 (C2V_135_638),
	.C2V_12 (C2V_135_742),
	.C2V_13 (C2V_135_873),
	.C2V_14 (C2V_135_917),
	.C2V_15 (C2V_135_990),
	.C2V_16 (C2V_135_1050),
	.C2V_17 (C2V_135_1080),
	.C2V_18 (C2V_135_1125),
	.C2V_19 (C2V_135_1286),
	.C2V_20 (C2V_135_1287),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU136 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_2_136),
	.V2C_2 (V2C_61_136),
	.V2C_3 (V2C_100_136),
	.V2C_4 (V2C_156_136),
	.V2C_5 (V2C_221_136),
	.V2C_6 (V2C_275_136),
	.V2C_7 (V2C_451_136),
	.V2C_8 (V2C_491_136),
	.V2C_9 (V2C_575_136),
	.V2C_10 (V2C_589_136),
	.V2C_11 (V2C_662_136),
	.V2C_12 (V2C_708_136),
	.V2C_13 (V2C_877_136),
	.V2C_14 (V2C_949_136),
	.V2C_15 (V2C_985_136),
	.V2C_16 (V2C_1015_136),
	.V2C_17 (V2C_1090_136),
	.V2C_18 (V2C_1106_136),
	.V2C_19 (V2C_1287_136),
	.V2C_20 (V2C_1288_136),
	.C2V_1 (C2V_136_2),
	.C2V_2 (C2V_136_61),
	.C2V_3 (C2V_136_100),
	.C2V_4 (C2V_136_156),
	.C2V_5 (C2V_136_221),
	.C2V_6 (C2V_136_275),
	.C2V_7 (C2V_136_451),
	.C2V_8 (C2V_136_491),
	.C2V_9 (C2V_136_575),
	.C2V_10 (C2V_136_589),
	.C2V_11 (C2V_136_662),
	.C2V_12 (C2V_136_708),
	.C2V_13 (C2V_136_877),
	.C2V_14 (C2V_136_949),
	.C2V_15 (C2V_136_985),
	.C2V_16 (C2V_136_1015),
	.C2V_17 (C2V_136_1090),
	.C2V_18 (C2V_136_1106),
	.C2V_19 (C2V_136_1287),
	.C2V_20 (C2V_136_1288),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU137 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_21_137),
	.V2C_2 (V2C_79_137),
	.V2C_3 (V2C_114_137),
	.V2C_4 (V2C_185_137),
	.V2C_5 (V2C_201_137),
	.V2C_6 (V2C_267_137),
	.V2C_7 (V2C_316_137),
	.V2C_8 (V2C_383_137),
	.V2C_9 (V2C_462_137),
	.V2C_10 (V2C_696_137),
	.V2C_11 (V2C_760_137),
	.V2C_12 (V2C_814_137),
	.V2C_13 (V2C_892_137),
	.V2C_14 (V2C_940_137),
	.V2C_15 (V2C_983_137),
	.V2C_16 (V2C_1035_137),
	.V2C_17 (V2C_1084_137),
	.V2C_18 (V2C_1132_137),
	.V2C_19 (V2C_1288_137),
	.V2C_20 (V2C_1289_137),
	.C2V_1 (C2V_137_21),
	.C2V_2 (C2V_137_79),
	.C2V_3 (C2V_137_114),
	.C2V_4 (C2V_137_185),
	.C2V_5 (C2V_137_201),
	.C2V_6 (C2V_137_267),
	.C2V_7 (C2V_137_316),
	.C2V_8 (C2V_137_383),
	.C2V_9 (C2V_137_462),
	.C2V_10 (C2V_137_696),
	.C2V_11 (C2V_137_760),
	.C2V_12 (C2V_137_814),
	.C2V_13 (C2V_137_892),
	.C2V_14 (C2V_137_940),
	.C2V_15 (C2V_137_983),
	.C2V_16 (C2V_137_1035),
	.C2V_17 (C2V_137_1084),
	.C2V_18 (C2V_137_1132),
	.C2V_19 (C2V_137_1288),
	.C2V_20 (C2V_137_1289),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU138 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_4_138),
	.V2C_2 (V2C_76_138),
	.V2C_3 (V2C_116_138),
	.V2C_4 (V2C_184_138),
	.V2C_5 (V2C_218_138),
	.V2C_6 (V2C_249_138),
	.V2C_7 (V2C_302_138),
	.V2C_8 (V2C_454_138),
	.V2C_9 (V2C_551_138),
	.V2C_10 (V2C_584_138),
	.V2C_11 (V2C_788_138),
	.V2C_12 (V2C_864_138),
	.V2C_13 (V2C_897_138),
	.V2C_14 (V2C_959_138),
	.V2C_15 (V2C_994_138),
	.V2C_16 (V2C_1013_138),
	.V2C_17 (V2C_1077_138),
	.V2C_18 (V2C_1127_138),
	.V2C_19 (V2C_1289_138),
	.V2C_20 (V2C_1290_138),
	.C2V_1 (C2V_138_4),
	.C2V_2 (C2V_138_76),
	.C2V_3 (C2V_138_116),
	.C2V_4 (C2V_138_184),
	.C2V_5 (C2V_138_218),
	.C2V_6 (C2V_138_249),
	.C2V_7 (C2V_138_302),
	.C2V_8 (C2V_138_454),
	.C2V_9 (C2V_138_551),
	.C2V_10 (C2V_138_584),
	.C2V_11 (C2V_138_788),
	.C2V_12 (C2V_138_864),
	.C2V_13 (C2V_138_897),
	.C2V_14 (C2V_138_959),
	.C2V_15 (C2V_138_994),
	.C2V_16 (C2V_138_1013),
	.C2V_17 (C2V_138_1077),
	.C2V_18 (C2V_138_1127),
	.C2V_19 (C2V_138_1289),
	.C2V_20 (C2V_138_1290),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU139 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_28_139),
	.V2C_2 (V2C_64_139),
	.V2C_3 (V2C_132_139),
	.V2C_4 (V2C_145_139),
	.V2C_5 (V2C_207_139),
	.V2C_6 (V2C_250_139),
	.V2C_7 (V2C_350_139),
	.V2C_8 (V2C_404_139),
	.V2C_9 (V2C_501_139),
	.V2C_10 (V2C_737_139),
	.V2C_11 (V2C_785_139),
	.V2C_12 (V2C_833_139),
	.V2C_13 (V2C_874_139),
	.V2C_14 (V2C_915_139),
	.V2C_15 (V2C_997_139),
	.V2C_16 (V2C_1036_139),
	.V2C_17 (V2C_1062_139),
	.V2C_18 (V2C_1121_139),
	.V2C_19 (V2C_1290_139),
	.V2C_20 (V2C_1291_139),
	.C2V_1 (C2V_139_28),
	.C2V_2 (C2V_139_64),
	.C2V_3 (C2V_139_132),
	.C2V_4 (C2V_139_145),
	.C2V_5 (C2V_139_207),
	.C2V_6 (C2V_139_250),
	.C2V_7 (C2V_139_350),
	.C2V_8 (C2V_139_404),
	.C2V_9 (C2V_139_501),
	.C2V_10 (C2V_139_737),
	.C2V_11 (C2V_139_785),
	.C2V_12 (C2V_139_833),
	.C2V_13 (C2V_139_874),
	.C2V_14 (C2V_139_915),
	.C2V_15 (C2V_139_997),
	.C2V_16 (C2V_139_1036),
	.C2V_17 (C2V_139_1062),
	.C2V_18 (C2V_139_1121),
	.C2V_19 (C2V_139_1290),
	.C2V_20 (C2V_139_1291),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU140 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_37_140),
	.V2C_2 (V2C_86_140),
	.V2C_3 (V2C_142_140),
	.V2C_4 (V2C_190_140),
	.V2C_5 (V2C_219_140),
	.V2C_6 (V2C_288_140),
	.V2C_7 (V2C_291_140),
	.V2C_8 (V2C_398_140),
	.V2C_9 (V2C_487_140),
	.V2C_10 (V2C_647_140),
	.V2C_11 (V2C_708_140),
	.V2C_12 (V2C_828_140),
	.V2C_13 (V2C_870_140),
	.V2C_14 (V2C_933_140),
	.V2C_15 (V2C_964_140),
	.V2C_16 (V2C_1044_140),
	.V2C_17 (V2C_1063_140),
	.V2C_18 (V2C_1142_140),
	.V2C_19 (V2C_1291_140),
	.V2C_20 (V2C_1292_140),
	.C2V_1 (C2V_140_37),
	.C2V_2 (C2V_140_86),
	.C2V_3 (C2V_140_142),
	.C2V_4 (C2V_140_190),
	.C2V_5 (C2V_140_219),
	.C2V_6 (C2V_140_288),
	.C2V_7 (C2V_140_291),
	.C2V_8 (C2V_140_398),
	.C2V_9 (C2V_140_487),
	.C2V_10 (C2V_140_647),
	.C2V_11 (C2V_140_708),
	.C2V_12 (C2V_140_828),
	.C2V_13 (C2V_140_870),
	.C2V_14 (C2V_140_933),
	.C2V_15 (C2V_140_964),
	.C2V_16 (C2V_140_1044),
	.C2V_17 (C2V_140_1063),
	.C2V_18 (C2V_140_1142),
	.C2V_19 (C2V_140_1291),
	.C2V_20 (C2V_140_1292),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU141 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_32_141),
	.V2C_2 (V2C_59_141),
	.V2C_3 (V2C_124_141),
	.V2C_4 (V2C_158_141),
	.V2C_5 (V2C_224_141),
	.V2C_6 (V2C_243_141),
	.V2C_7 (V2C_340_141),
	.V2C_8 (V2C_395_141),
	.V2C_9 (V2C_554_141),
	.V2C_10 (V2C_611_141),
	.V2C_11 (V2C_639_141),
	.V2C_12 (V2C_743_141),
	.V2C_13 (V2C_874_141),
	.V2C_14 (V2C_918_141),
	.V2C_15 (V2C_991_141),
	.V2C_16 (V2C_1051_141),
	.V2C_17 (V2C_1081_141),
	.V2C_18 (V2C_1126_141),
	.V2C_19 (V2C_1292_141),
	.V2C_20 (V2C_1293_141),
	.C2V_1 (C2V_141_32),
	.C2V_2 (C2V_141_59),
	.C2V_3 (C2V_141_124),
	.C2V_4 (C2V_141_158),
	.C2V_5 (C2V_141_224),
	.C2V_6 (C2V_141_243),
	.C2V_7 (C2V_141_340),
	.C2V_8 (C2V_141_395),
	.C2V_9 (C2V_141_554),
	.C2V_10 (C2V_141_611),
	.C2V_11 (C2V_141_639),
	.C2V_12 (C2V_141_743),
	.C2V_13 (C2V_141_874),
	.C2V_14 (C2V_141_918),
	.C2V_15 (C2V_141_991),
	.C2V_16 (C2V_141_1051),
	.C2V_17 (C2V_141_1081),
	.C2V_18 (C2V_141_1126),
	.C2V_19 (C2V_141_1292),
	.C2V_20 (C2V_141_1293),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU142 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_3_142),
	.V2C_2 (V2C_62_142),
	.V2C_3 (V2C_101_142),
	.V2C_4 (V2C_157_142),
	.V2C_5 (V2C_222_142),
	.V2C_6 (V2C_276_142),
	.V2C_7 (V2C_452_142),
	.V2C_8 (V2C_492_142),
	.V2C_9 (V2C_576_142),
	.V2C_10 (V2C_590_142),
	.V2C_11 (V2C_663_142),
	.V2C_12 (V2C_709_142),
	.V2C_13 (V2C_878_142),
	.V2C_14 (V2C_950_142),
	.V2C_15 (V2C_986_142),
	.V2C_16 (V2C_1016_142),
	.V2C_17 (V2C_1091_142),
	.V2C_18 (V2C_1107_142),
	.V2C_19 (V2C_1293_142),
	.V2C_20 (V2C_1294_142),
	.C2V_1 (C2V_142_3),
	.C2V_2 (C2V_142_62),
	.C2V_3 (C2V_142_101),
	.C2V_4 (C2V_142_157),
	.C2V_5 (C2V_142_222),
	.C2V_6 (C2V_142_276),
	.C2V_7 (C2V_142_452),
	.C2V_8 (C2V_142_492),
	.C2V_9 (C2V_142_576),
	.C2V_10 (C2V_142_590),
	.C2V_11 (C2V_142_663),
	.C2V_12 (C2V_142_709),
	.C2V_13 (C2V_142_878),
	.C2V_14 (C2V_142_950),
	.C2V_15 (C2V_142_986),
	.C2V_16 (C2V_142_1016),
	.C2V_17 (C2V_142_1091),
	.C2V_18 (C2V_142_1107),
	.C2V_19 (C2V_142_1293),
	.C2V_20 (C2V_142_1294),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU143 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_22_143),
	.V2C_2 (V2C_80_143),
	.V2C_3 (V2C_115_143),
	.V2C_4 (V2C_186_143),
	.V2C_5 (V2C_202_143),
	.V2C_6 (V2C_268_143),
	.V2C_7 (V2C_317_143),
	.V2C_8 (V2C_384_143),
	.V2C_9 (V2C_463_143),
	.V2C_10 (V2C_697_143),
	.V2C_11 (V2C_761_143),
	.V2C_12 (V2C_815_143),
	.V2C_13 (V2C_893_143),
	.V2C_14 (V2C_941_143),
	.V2C_15 (V2C_984_143),
	.V2C_16 (V2C_1036_143),
	.V2C_17 (V2C_1085_143),
	.V2C_18 (V2C_1133_143),
	.V2C_19 (V2C_1294_143),
	.V2C_20 (V2C_1295_143),
	.C2V_1 (C2V_143_22),
	.C2V_2 (C2V_143_80),
	.C2V_3 (C2V_143_115),
	.C2V_4 (C2V_143_186),
	.C2V_5 (C2V_143_202),
	.C2V_6 (C2V_143_268),
	.C2V_7 (C2V_143_317),
	.C2V_8 (C2V_143_384),
	.C2V_9 (C2V_143_463),
	.C2V_10 (C2V_143_697),
	.C2V_11 (C2V_143_761),
	.C2V_12 (C2V_143_815),
	.C2V_13 (C2V_143_893),
	.C2V_14 (C2V_143_941),
	.C2V_15 (C2V_143_984),
	.C2V_16 (C2V_143_1036),
	.C2V_17 (C2V_143_1085),
	.C2V_18 (C2V_143_1133),
	.C2V_19 (C2V_143_1294),
	.C2V_20 (C2V_143_1295),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU144 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_5_144),
	.V2C_2 (V2C_77_144),
	.V2C_3 (V2C_117_144),
	.V2C_4 (V2C_185_144),
	.V2C_5 (V2C_219_144),
	.V2C_6 (V2C_250_144),
	.V2C_7 (V2C_303_144),
	.V2C_8 (V2C_455_144),
	.V2C_9 (V2C_552_144),
	.V2C_10 (V2C_585_144),
	.V2C_11 (V2C_789_144),
	.V2C_12 (V2C_817_144),
	.V2C_13 (V2C_898_144),
	.V2C_14 (V2C_960_144),
	.V2C_15 (V2C_995_144),
	.V2C_16 (V2C_1014_144),
	.V2C_17 (V2C_1078_144),
	.V2C_18 (V2C_1128_144),
	.V2C_19 (V2C_1295_144),
	.V2C_20 (V2C_1296_144),
	.C2V_1 (C2V_144_5),
	.C2V_2 (C2V_144_77),
	.C2V_3 (C2V_144_117),
	.C2V_4 (C2V_144_185),
	.C2V_5 (C2V_144_219),
	.C2V_6 (C2V_144_250),
	.C2V_7 (C2V_144_303),
	.C2V_8 (C2V_144_455),
	.C2V_9 (C2V_144_552),
	.C2V_10 (C2V_144_585),
	.C2V_11 (C2V_144_789),
	.C2V_12 (C2V_144_817),
	.C2V_13 (C2V_144_898),
	.C2V_14 (C2V_144_960),
	.C2V_15 (C2V_144_995),
	.C2V_16 (C2V_144_1014),
	.C2V_17 (C2V_144_1078),
	.C2V_18 (C2V_144_1128),
	.C2V_19 (C2V_144_1295),
	.C2V_20 (C2V_144_1296),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU145 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_29_145),
	.V2C_2 (V2C_65_145),
	.V2C_3 (V2C_133_145),
	.V2C_4 (V2C_146_145),
	.V2C_5 (V2C_208_145),
	.V2C_6 (V2C_251_145),
	.V2C_7 (V2C_351_145),
	.V2C_8 (V2C_405_145),
	.V2C_9 (V2C_502_145),
	.V2C_10 (V2C_738_145),
	.V2C_11 (V2C_786_145),
	.V2C_12 (V2C_834_145),
	.V2C_13 (V2C_875_145),
	.V2C_14 (V2C_916_145),
	.V2C_15 (V2C_998_145),
	.V2C_16 (V2C_1037_145),
	.V2C_17 (V2C_1063_145),
	.V2C_18 (V2C_1122_145),
	.V2C_19 (V2C_1296_145),
	.V2C_20 (V2C_1297_145),
	.C2V_1 (C2V_145_29),
	.C2V_2 (C2V_145_65),
	.C2V_3 (C2V_145_133),
	.C2V_4 (C2V_145_146),
	.C2V_5 (C2V_145_208),
	.C2V_6 (C2V_145_251),
	.C2V_7 (C2V_145_351),
	.C2V_8 (C2V_145_405),
	.C2V_9 (C2V_145_502),
	.C2V_10 (C2V_145_738),
	.C2V_11 (C2V_145_786),
	.C2V_12 (C2V_145_834),
	.C2V_13 (C2V_145_875),
	.C2V_14 (C2V_145_916),
	.C2V_15 (C2V_145_998),
	.C2V_16 (C2V_145_1037),
	.C2V_17 (C2V_145_1063),
	.C2V_18 (C2V_145_1122),
	.C2V_19 (C2V_145_1296),
	.C2V_20 (C2V_145_1297),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU146 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_38_146),
	.V2C_2 (V2C_87_146),
	.V2C_3 (V2C_143_146),
	.V2C_4 (V2C_191_146),
	.V2C_5 (V2C_220_146),
	.V2C_6 (V2C_241_146),
	.V2C_7 (V2C_292_146),
	.V2C_8 (V2C_399_146),
	.V2C_9 (V2C_488_146),
	.V2C_10 (V2C_648_146),
	.V2C_11 (V2C_709_146),
	.V2C_12 (V2C_829_146),
	.V2C_13 (V2C_871_146),
	.V2C_14 (V2C_934_146),
	.V2C_15 (V2C_965_146),
	.V2C_16 (V2C_1045_146),
	.V2C_17 (V2C_1064_146),
	.V2C_18 (V2C_1143_146),
	.V2C_19 (V2C_1297_146),
	.V2C_20 (V2C_1298_146),
	.C2V_1 (C2V_146_38),
	.C2V_2 (C2V_146_87),
	.C2V_3 (C2V_146_143),
	.C2V_4 (C2V_146_191),
	.C2V_5 (C2V_146_220),
	.C2V_6 (C2V_146_241),
	.C2V_7 (C2V_146_292),
	.C2V_8 (C2V_146_399),
	.C2V_9 (C2V_146_488),
	.C2V_10 (C2V_146_648),
	.C2V_11 (C2V_146_709),
	.C2V_12 (C2V_146_829),
	.C2V_13 (C2V_146_871),
	.C2V_14 (C2V_146_934),
	.C2V_15 (C2V_146_965),
	.C2V_16 (C2V_146_1045),
	.C2V_17 (C2V_146_1064),
	.C2V_18 (C2V_146_1143),
	.C2V_19 (C2V_146_1297),
	.C2V_20 (C2V_146_1298),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU147 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_33_147),
	.V2C_2 (V2C_60_147),
	.V2C_3 (V2C_125_147),
	.V2C_4 (V2C_159_147),
	.V2C_5 (V2C_225_147),
	.V2C_6 (V2C_244_147),
	.V2C_7 (V2C_341_147),
	.V2C_8 (V2C_396_147),
	.V2C_9 (V2C_555_147),
	.V2C_10 (V2C_612_147),
	.V2C_11 (V2C_640_147),
	.V2C_12 (V2C_744_147),
	.V2C_13 (V2C_875_147),
	.V2C_14 (V2C_919_147),
	.V2C_15 (V2C_992_147),
	.V2C_16 (V2C_1052_147),
	.V2C_17 (V2C_1082_147),
	.V2C_18 (V2C_1127_147),
	.V2C_19 (V2C_1298_147),
	.V2C_20 (V2C_1299_147),
	.C2V_1 (C2V_147_33),
	.C2V_2 (C2V_147_60),
	.C2V_3 (C2V_147_125),
	.C2V_4 (C2V_147_159),
	.C2V_5 (C2V_147_225),
	.C2V_6 (C2V_147_244),
	.C2V_7 (C2V_147_341),
	.C2V_8 (C2V_147_396),
	.C2V_9 (C2V_147_555),
	.C2V_10 (C2V_147_612),
	.C2V_11 (C2V_147_640),
	.C2V_12 (C2V_147_744),
	.C2V_13 (C2V_147_875),
	.C2V_14 (C2V_147_919),
	.C2V_15 (C2V_147_992),
	.C2V_16 (C2V_147_1052),
	.C2V_17 (C2V_147_1082),
	.C2V_18 (C2V_147_1127),
	.C2V_19 (C2V_147_1298),
	.C2V_20 (C2V_147_1299),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU148 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_4_148),
	.V2C_2 (V2C_63_148),
	.V2C_3 (V2C_102_148),
	.V2C_4 (V2C_158_148),
	.V2C_5 (V2C_223_148),
	.V2C_6 (V2C_277_148),
	.V2C_7 (V2C_453_148),
	.V2C_8 (V2C_493_148),
	.V2C_9 (V2C_529_148),
	.V2C_10 (V2C_591_148),
	.V2C_11 (V2C_664_148),
	.V2C_12 (V2C_710_148),
	.V2C_13 (V2C_879_148),
	.V2C_14 (V2C_951_148),
	.V2C_15 (V2C_987_148),
	.V2C_16 (V2C_1017_148),
	.V2C_17 (V2C_1092_148),
	.V2C_18 (V2C_1108_148),
	.V2C_19 (V2C_1299_148),
	.V2C_20 (V2C_1300_148),
	.C2V_1 (C2V_148_4),
	.C2V_2 (C2V_148_63),
	.C2V_3 (C2V_148_102),
	.C2V_4 (C2V_148_158),
	.C2V_5 (C2V_148_223),
	.C2V_6 (C2V_148_277),
	.C2V_7 (C2V_148_453),
	.C2V_8 (C2V_148_493),
	.C2V_9 (C2V_148_529),
	.C2V_10 (C2V_148_591),
	.C2V_11 (C2V_148_664),
	.C2V_12 (C2V_148_710),
	.C2V_13 (C2V_148_879),
	.C2V_14 (C2V_148_951),
	.C2V_15 (C2V_148_987),
	.C2V_16 (C2V_148_1017),
	.C2V_17 (C2V_148_1092),
	.C2V_18 (C2V_148_1108),
	.C2V_19 (C2V_148_1299),
	.C2V_20 (C2V_148_1300),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU149 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_23_149),
	.V2C_2 (V2C_81_149),
	.V2C_3 (V2C_116_149),
	.V2C_4 (V2C_187_149),
	.V2C_5 (V2C_203_149),
	.V2C_6 (V2C_269_149),
	.V2C_7 (V2C_318_149),
	.V2C_8 (V2C_337_149),
	.V2C_9 (V2C_464_149),
	.V2C_10 (V2C_698_149),
	.V2C_11 (V2C_762_149),
	.V2C_12 (V2C_816_149),
	.V2C_13 (V2C_894_149),
	.V2C_14 (V2C_942_149),
	.V2C_15 (V2C_985_149),
	.V2C_16 (V2C_1037_149),
	.V2C_17 (V2C_1086_149),
	.V2C_18 (V2C_1134_149),
	.V2C_19 (V2C_1300_149),
	.V2C_20 (V2C_1301_149),
	.C2V_1 (C2V_149_23),
	.C2V_2 (C2V_149_81),
	.C2V_3 (C2V_149_116),
	.C2V_4 (C2V_149_187),
	.C2V_5 (C2V_149_203),
	.C2V_6 (C2V_149_269),
	.C2V_7 (C2V_149_318),
	.C2V_8 (C2V_149_337),
	.C2V_9 (C2V_149_464),
	.C2V_10 (C2V_149_698),
	.C2V_11 (C2V_149_762),
	.C2V_12 (C2V_149_816),
	.C2V_13 (C2V_149_894),
	.C2V_14 (C2V_149_942),
	.C2V_15 (C2V_149_985),
	.C2V_16 (C2V_149_1037),
	.C2V_17 (C2V_149_1086),
	.C2V_18 (C2V_149_1134),
	.C2V_19 (C2V_149_1300),
	.C2V_20 (C2V_149_1301),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU150 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_6_150),
	.V2C_2 (V2C_78_150),
	.V2C_3 (V2C_118_150),
	.V2C_4 (V2C_186_150),
	.V2C_5 (V2C_220_150),
	.V2C_6 (V2C_251_150),
	.V2C_7 (V2C_304_150),
	.V2C_8 (V2C_456_150),
	.V2C_9 (V2C_553_150),
	.V2C_10 (V2C_586_150),
	.V2C_11 (V2C_790_150),
	.V2C_12 (V2C_818_150),
	.V2C_13 (V2C_899_150),
	.V2C_14 (V2C_913_150),
	.V2C_15 (V2C_996_150),
	.V2C_16 (V2C_1015_150),
	.V2C_17 (V2C_1079_150),
	.V2C_18 (V2C_1129_150),
	.V2C_19 (V2C_1301_150),
	.V2C_20 (V2C_1302_150),
	.C2V_1 (C2V_150_6),
	.C2V_2 (C2V_150_78),
	.C2V_3 (C2V_150_118),
	.C2V_4 (C2V_150_186),
	.C2V_5 (C2V_150_220),
	.C2V_6 (C2V_150_251),
	.C2V_7 (C2V_150_304),
	.C2V_8 (C2V_150_456),
	.C2V_9 (C2V_150_553),
	.C2V_10 (C2V_150_586),
	.C2V_11 (C2V_150_790),
	.C2V_12 (C2V_150_818),
	.C2V_13 (C2V_150_899),
	.C2V_14 (C2V_150_913),
	.C2V_15 (C2V_150_996),
	.C2V_16 (C2V_150_1015),
	.C2V_17 (C2V_150_1079),
	.C2V_18 (C2V_150_1129),
	.C2V_19 (C2V_150_1301),
	.C2V_20 (C2V_150_1302),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU151 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_30_151),
	.V2C_2 (V2C_66_151),
	.V2C_3 (V2C_134_151),
	.V2C_4 (V2C_147_151),
	.V2C_5 (V2C_209_151),
	.V2C_6 (V2C_252_151),
	.V2C_7 (V2C_352_151),
	.V2C_8 (V2C_406_151),
	.V2C_9 (V2C_503_151),
	.V2C_10 (V2C_739_151),
	.V2C_11 (V2C_787_151),
	.V2C_12 (V2C_835_151),
	.V2C_13 (V2C_876_151),
	.V2C_14 (V2C_917_151),
	.V2C_15 (V2C_999_151),
	.V2C_16 (V2C_1038_151),
	.V2C_17 (V2C_1064_151),
	.V2C_18 (V2C_1123_151),
	.V2C_19 (V2C_1302_151),
	.V2C_20 (V2C_1303_151),
	.C2V_1 (C2V_151_30),
	.C2V_2 (C2V_151_66),
	.C2V_3 (C2V_151_134),
	.C2V_4 (C2V_151_147),
	.C2V_5 (C2V_151_209),
	.C2V_6 (C2V_151_252),
	.C2V_7 (C2V_151_352),
	.C2V_8 (C2V_151_406),
	.C2V_9 (C2V_151_503),
	.C2V_10 (C2V_151_739),
	.C2V_11 (C2V_151_787),
	.C2V_12 (C2V_151_835),
	.C2V_13 (C2V_151_876),
	.C2V_14 (C2V_151_917),
	.C2V_15 (C2V_151_999),
	.C2V_16 (C2V_151_1038),
	.C2V_17 (C2V_151_1064),
	.C2V_18 (C2V_151_1123),
	.C2V_19 (C2V_151_1302),
	.C2V_20 (C2V_151_1303),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU152 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_39_152),
	.V2C_2 (V2C_88_152),
	.V2C_3 (V2C_144_152),
	.V2C_4 (V2C_192_152),
	.V2C_5 (V2C_221_152),
	.V2C_6 (V2C_242_152),
	.V2C_7 (V2C_293_152),
	.V2C_8 (V2C_400_152),
	.V2C_9 (V2C_489_152),
	.V2C_10 (V2C_649_152),
	.V2C_11 (V2C_710_152),
	.V2C_12 (V2C_830_152),
	.V2C_13 (V2C_872_152),
	.V2C_14 (V2C_935_152),
	.V2C_15 (V2C_966_152),
	.V2C_16 (V2C_1046_152),
	.V2C_17 (V2C_1065_152),
	.V2C_18 (V2C_1144_152),
	.V2C_19 (V2C_1303_152),
	.V2C_20 (V2C_1304_152),
	.C2V_1 (C2V_152_39),
	.C2V_2 (C2V_152_88),
	.C2V_3 (C2V_152_144),
	.C2V_4 (C2V_152_192),
	.C2V_5 (C2V_152_221),
	.C2V_6 (C2V_152_242),
	.C2V_7 (C2V_152_293),
	.C2V_8 (C2V_152_400),
	.C2V_9 (C2V_152_489),
	.C2V_10 (C2V_152_649),
	.C2V_11 (C2V_152_710),
	.C2V_12 (C2V_152_830),
	.C2V_13 (C2V_152_872),
	.C2V_14 (C2V_152_935),
	.C2V_15 (C2V_152_966),
	.C2V_16 (C2V_152_1046),
	.C2V_17 (C2V_152_1065),
	.C2V_18 (C2V_152_1144),
	.C2V_19 (C2V_152_1303),
	.C2V_20 (C2V_152_1304),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU153 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_34_153),
	.V2C_2 (V2C_61_153),
	.V2C_3 (V2C_126_153),
	.V2C_4 (V2C_160_153),
	.V2C_5 (V2C_226_153),
	.V2C_6 (V2C_245_153),
	.V2C_7 (V2C_342_153),
	.V2C_8 (V2C_397_153),
	.V2C_9 (V2C_556_153),
	.V2C_10 (V2C_613_153),
	.V2C_11 (V2C_641_153),
	.V2C_12 (V2C_745_153),
	.V2C_13 (V2C_876_153),
	.V2C_14 (V2C_920_153),
	.V2C_15 (V2C_993_153),
	.V2C_16 (V2C_1053_153),
	.V2C_17 (V2C_1083_153),
	.V2C_18 (V2C_1128_153),
	.V2C_19 (V2C_1304_153),
	.V2C_20 (V2C_1305_153),
	.C2V_1 (C2V_153_34),
	.C2V_2 (C2V_153_61),
	.C2V_3 (C2V_153_126),
	.C2V_4 (C2V_153_160),
	.C2V_5 (C2V_153_226),
	.C2V_6 (C2V_153_245),
	.C2V_7 (C2V_153_342),
	.C2V_8 (C2V_153_397),
	.C2V_9 (C2V_153_556),
	.C2V_10 (C2V_153_613),
	.C2V_11 (C2V_153_641),
	.C2V_12 (C2V_153_745),
	.C2V_13 (C2V_153_876),
	.C2V_14 (C2V_153_920),
	.C2V_15 (C2V_153_993),
	.C2V_16 (C2V_153_1053),
	.C2V_17 (C2V_153_1083),
	.C2V_18 (C2V_153_1128),
	.C2V_19 (C2V_153_1304),
	.C2V_20 (C2V_153_1305),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU154 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_5_154),
	.V2C_2 (V2C_64_154),
	.V2C_3 (V2C_103_154),
	.V2C_4 (V2C_159_154),
	.V2C_5 (V2C_224_154),
	.V2C_6 (V2C_278_154),
	.V2C_7 (V2C_454_154),
	.V2C_8 (V2C_494_154),
	.V2C_9 (V2C_530_154),
	.V2C_10 (V2C_592_154),
	.V2C_11 (V2C_665_154),
	.V2C_12 (V2C_711_154),
	.V2C_13 (V2C_880_154),
	.V2C_14 (V2C_952_154),
	.V2C_15 (V2C_988_154),
	.V2C_16 (V2C_1018_154),
	.V2C_17 (V2C_1093_154),
	.V2C_18 (V2C_1109_154),
	.V2C_19 (V2C_1305_154),
	.V2C_20 (V2C_1306_154),
	.C2V_1 (C2V_154_5),
	.C2V_2 (C2V_154_64),
	.C2V_3 (C2V_154_103),
	.C2V_4 (C2V_154_159),
	.C2V_5 (C2V_154_224),
	.C2V_6 (C2V_154_278),
	.C2V_7 (C2V_154_454),
	.C2V_8 (C2V_154_494),
	.C2V_9 (C2V_154_530),
	.C2V_10 (C2V_154_592),
	.C2V_11 (C2V_154_665),
	.C2V_12 (C2V_154_711),
	.C2V_13 (C2V_154_880),
	.C2V_14 (C2V_154_952),
	.C2V_15 (C2V_154_988),
	.C2V_16 (C2V_154_1018),
	.C2V_17 (C2V_154_1093),
	.C2V_18 (C2V_154_1109),
	.C2V_19 (C2V_154_1305),
	.C2V_20 (C2V_154_1306),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU155 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_24_155),
	.V2C_2 (V2C_82_155),
	.V2C_3 (V2C_117_155),
	.V2C_4 (V2C_188_155),
	.V2C_5 (V2C_204_155),
	.V2C_6 (V2C_270_155),
	.V2C_7 (V2C_319_155),
	.V2C_8 (V2C_338_155),
	.V2C_9 (V2C_465_155),
	.V2C_10 (V2C_699_155),
	.V2C_11 (V2C_763_155),
	.V2C_12 (V2C_769_155),
	.V2C_13 (V2C_895_155),
	.V2C_14 (V2C_943_155),
	.V2C_15 (V2C_986_155),
	.V2C_16 (V2C_1038_155),
	.V2C_17 (V2C_1087_155),
	.V2C_18 (V2C_1135_155),
	.V2C_19 (V2C_1306_155),
	.V2C_20 (V2C_1307_155),
	.C2V_1 (C2V_155_24),
	.C2V_2 (C2V_155_82),
	.C2V_3 (C2V_155_117),
	.C2V_4 (C2V_155_188),
	.C2V_5 (C2V_155_204),
	.C2V_6 (C2V_155_270),
	.C2V_7 (C2V_155_319),
	.C2V_8 (C2V_155_338),
	.C2V_9 (C2V_155_465),
	.C2V_10 (C2V_155_699),
	.C2V_11 (C2V_155_763),
	.C2V_12 (C2V_155_769),
	.C2V_13 (C2V_155_895),
	.C2V_14 (C2V_155_943),
	.C2V_15 (C2V_155_986),
	.C2V_16 (C2V_155_1038),
	.C2V_17 (C2V_155_1087),
	.C2V_18 (C2V_155_1135),
	.C2V_19 (C2V_155_1306),
	.C2V_20 (C2V_155_1307),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU156 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_7_156),
	.V2C_2 (V2C_79_156),
	.V2C_3 (V2C_119_156),
	.V2C_4 (V2C_187_156),
	.V2C_5 (V2C_221_156),
	.V2C_6 (V2C_252_156),
	.V2C_7 (V2C_305_156),
	.V2C_8 (V2C_457_156),
	.V2C_9 (V2C_554_156),
	.V2C_10 (V2C_587_156),
	.V2C_11 (V2C_791_156),
	.V2C_12 (V2C_819_156),
	.V2C_13 (V2C_900_156),
	.V2C_14 (V2C_914_156),
	.V2C_15 (V2C_997_156),
	.V2C_16 (V2C_1016_156),
	.V2C_17 (V2C_1080_156),
	.V2C_18 (V2C_1130_156),
	.V2C_19 (V2C_1307_156),
	.V2C_20 (V2C_1308_156),
	.C2V_1 (C2V_156_7),
	.C2V_2 (C2V_156_79),
	.C2V_3 (C2V_156_119),
	.C2V_4 (C2V_156_187),
	.C2V_5 (C2V_156_221),
	.C2V_6 (C2V_156_252),
	.C2V_7 (C2V_156_305),
	.C2V_8 (C2V_156_457),
	.C2V_9 (C2V_156_554),
	.C2V_10 (C2V_156_587),
	.C2V_11 (C2V_156_791),
	.C2V_12 (C2V_156_819),
	.C2V_13 (C2V_156_900),
	.C2V_14 (C2V_156_914),
	.C2V_15 (C2V_156_997),
	.C2V_16 (C2V_156_1016),
	.C2V_17 (C2V_156_1080),
	.C2V_18 (C2V_156_1130),
	.C2V_19 (C2V_156_1307),
	.C2V_20 (C2V_156_1308),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU157 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_31_157),
	.V2C_2 (V2C_67_157),
	.V2C_3 (V2C_135_157),
	.V2C_4 (V2C_148_157),
	.V2C_5 (V2C_210_157),
	.V2C_6 (V2C_253_157),
	.V2C_7 (V2C_353_157),
	.V2C_8 (V2C_407_157),
	.V2C_9 (V2C_504_157),
	.V2C_10 (V2C_740_157),
	.V2C_11 (V2C_788_157),
	.V2C_12 (V2C_836_157),
	.V2C_13 (V2C_877_157),
	.V2C_14 (V2C_918_157),
	.V2C_15 (V2C_1000_157),
	.V2C_16 (V2C_1039_157),
	.V2C_17 (V2C_1065_157),
	.V2C_18 (V2C_1124_157),
	.V2C_19 (V2C_1308_157),
	.V2C_20 (V2C_1309_157),
	.C2V_1 (C2V_157_31),
	.C2V_2 (C2V_157_67),
	.C2V_3 (C2V_157_135),
	.C2V_4 (C2V_157_148),
	.C2V_5 (C2V_157_210),
	.C2V_6 (C2V_157_253),
	.C2V_7 (C2V_157_353),
	.C2V_8 (C2V_157_407),
	.C2V_9 (C2V_157_504),
	.C2V_10 (C2V_157_740),
	.C2V_11 (C2V_157_788),
	.C2V_12 (C2V_157_836),
	.C2V_13 (C2V_157_877),
	.C2V_14 (C2V_157_918),
	.C2V_15 (C2V_157_1000),
	.C2V_16 (C2V_157_1039),
	.C2V_17 (C2V_157_1065),
	.C2V_18 (C2V_157_1124),
	.C2V_19 (C2V_157_1308),
	.C2V_20 (C2V_157_1309),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU158 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_40_158),
	.V2C_2 (V2C_89_158),
	.V2C_3 (V2C_97_158),
	.V2C_4 (V2C_145_158),
	.V2C_5 (V2C_222_158),
	.V2C_6 (V2C_243_158),
	.V2C_7 (V2C_294_158),
	.V2C_8 (V2C_401_158),
	.V2C_9 (V2C_490_158),
	.V2C_10 (V2C_650_158),
	.V2C_11 (V2C_711_158),
	.V2C_12 (V2C_831_158),
	.V2C_13 (V2C_873_158),
	.V2C_14 (V2C_936_158),
	.V2C_15 (V2C_967_158),
	.V2C_16 (V2C_1047_158),
	.V2C_17 (V2C_1066_158),
	.V2C_18 (V2C_1145_158),
	.V2C_19 (V2C_1309_158),
	.V2C_20 (V2C_1310_158),
	.C2V_1 (C2V_158_40),
	.C2V_2 (C2V_158_89),
	.C2V_3 (C2V_158_97),
	.C2V_4 (C2V_158_145),
	.C2V_5 (C2V_158_222),
	.C2V_6 (C2V_158_243),
	.C2V_7 (C2V_158_294),
	.C2V_8 (C2V_158_401),
	.C2V_9 (C2V_158_490),
	.C2V_10 (C2V_158_650),
	.C2V_11 (C2V_158_711),
	.C2V_12 (C2V_158_831),
	.C2V_13 (C2V_158_873),
	.C2V_14 (C2V_158_936),
	.C2V_15 (C2V_158_967),
	.C2V_16 (C2V_158_1047),
	.C2V_17 (C2V_158_1066),
	.C2V_18 (C2V_158_1145),
	.C2V_19 (C2V_158_1309),
	.C2V_20 (C2V_158_1310),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU159 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_35_159),
	.V2C_2 (V2C_62_159),
	.V2C_3 (V2C_127_159),
	.V2C_4 (V2C_161_159),
	.V2C_5 (V2C_227_159),
	.V2C_6 (V2C_246_159),
	.V2C_7 (V2C_343_159),
	.V2C_8 (V2C_398_159),
	.V2C_9 (V2C_557_159),
	.V2C_10 (V2C_614_159),
	.V2C_11 (V2C_642_159),
	.V2C_12 (V2C_746_159),
	.V2C_13 (V2C_877_159),
	.V2C_14 (V2C_921_159),
	.V2C_15 (V2C_994_159),
	.V2C_16 (V2C_1054_159),
	.V2C_17 (V2C_1084_159),
	.V2C_18 (V2C_1129_159),
	.V2C_19 (V2C_1310_159),
	.V2C_20 (V2C_1311_159),
	.C2V_1 (C2V_159_35),
	.C2V_2 (C2V_159_62),
	.C2V_3 (C2V_159_127),
	.C2V_4 (C2V_159_161),
	.C2V_5 (C2V_159_227),
	.C2V_6 (C2V_159_246),
	.C2V_7 (C2V_159_343),
	.C2V_8 (C2V_159_398),
	.C2V_9 (C2V_159_557),
	.C2V_10 (C2V_159_614),
	.C2V_11 (C2V_159_642),
	.C2V_12 (C2V_159_746),
	.C2V_13 (C2V_159_877),
	.C2V_14 (C2V_159_921),
	.C2V_15 (C2V_159_994),
	.C2V_16 (C2V_159_1054),
	.C2V_17 (C2V_159_1084),
	.C2V_18 (C2V_159_1129),
	.C2V_19 (C2V_159_1310),
	.C2V_20 (C2V_159_1311),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU160 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_6_160),
	.V2C_2 (V2C_65_160),
	.V2C_3 (V2C_104_160),
	.V2C_4 (V2C_160_160),
	.V2C_5 (V2C_225_160),
	.V2C_6 (V2C_279_160),
	.V2C_7 (V2C_455_160),
	.V2C_8 (V2C_495_160),
	.V2C_9 (V2C_531_160),
	.V2C_10 (V2C_593_160),
	.V2C_11 (V2C_666_160),
	.V2C_12 (V2C_712_160),
	.V2C_13 (V2C_881_160),
	.V2C_14 (V2C_953_160),
	.V2C_15 (V2C_989_160),
	.V2C_16 (V2C_1019_160),
	.V2C_17 (V2C_1094_160),
	.V2C_18 (V2C_1110_160),
	.V2C_19 (V2C_1311_160),
	.V2C_20 (V2C_1312_160),
	.C2V_1 (C2V_160_6),
	.C2V_2 (C2V_160_65),
	.C2V_3 (C2V_160_104),
	.C2V_4 (C2V_160_160),
	.C2V_5 (C2V_160_225),
	.C2V_6 (C2V_160_279),
	.C2V_7 (C2V_160_455),
	.C2V_8 (C2V_160_495),
	.C2V_9 (C2V_160_531),
	.C2V_10 (C2V_160_593),
	.C2V_11 (C2V_160_666),
	.C2V_12 (C2V_160_712),
	.C2V_13 (C2V_160_881),
	.C2V_14 (C2V_160_953),
	.C2V_15 (C2V_160_989),
	.C2V_16 (C2V_160_1019),
	.C2V_17 (C2V_160_1094),
	.C2V_18 (C2V_160_1110),
	.C2V_19 (C2V_160_1311),
	.C2V_20 (C2V_160_1312),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU161 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_25_161),
	.V2C_2 (V2C_83_161),
	.V2C_3 (V2C_118_161),
	.V2C_4 (V2C_189_161),
	.V2C_5 (V2C_205_161),
	.V2C_6 (V2C_271_161),
	.V2C_7 (V2C_320_161),
	.V2C_8 (V2C_339_161),
	.V2C_9 (V2C_466_161),
	.V2C_10 (V2C_700_161),
	.V2C_11 (V2C_764_161),
	.V2C_12 (V2C_770_161),
	.V2C_13 (V2C_896_161),
	.V2C_14 (V2C_944_161),
	.V2C_15 (V2C_987_161),
	.V2C_16 (V2C_1039_161),
	.V2C_17 (V2C_1088_161),
	.V2C_18 (V2C_1136_161),
	.V2C_19 (V2C_1312_161),
	.V2C_20 (V2C_1313_161),
	.C2V_1 (C2V_161_25),
	.C2V_2 (C2V_161_83),
	.C2V_3 (C2V_161_118),
	.C2V_4 (C2V_161_189),
	.C2V_5 (C2V_161_205),
	.C2V_6 (C2V_161_271),
	.C2V_7 (C2V_161_320),
	.C2V_8 (C2V_161_339),
	.C2V_9 (C2V_161_466),
	.C2V_10 (C2V_161_700),
	.C2V_11 (C2V_161_764),
	.C2V_12 (C2V_161_770),
	.C2V_13 (C2V_161_896),
	.C2V_14 (C2V_161_944),
	.C2V_15 (C2V_161_987),
	.C2V_16 (C2V_161_1039),
	.C2V_17 (C2V_161_1088),
	.C2V_18 (C2V_161_1136),
	.C2V_19 (C2V_161_1312),
	.C2V_20 (C2V_161_1313),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU162 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_8_162),
	.V2C_2 (V2C_80_162),
	.V2C_3 (V2C_120_162),
	.V2C_4 (V2C_188_162),
	.V2C_5 (V2C_222_162),
	.V2C_6 (V2C_253_162),
	.V2C_7 (V2C_306_162),
	.V2C_8 (V2C_458_162),
	.V2C_9 (V2C_555_162),
	.V2C_10 (V2C_588_162),
	.V2C_11 (V2C_792_162),
	.V2C_12 (V2C_820_162),
	.V2C_13 (V2C_901_162),
	.V2C_14 (V2C_915_162),
	.V2C_15 (V2C_998_162),
	.V2C_16 (V2C_1017_162),
	.V2C_17 (V2C_1081_162),
	.V2C_18 (V2C_1131_162),
	.V2C_19 (V2C_1313_162),
	.V2C_20 (V2C_1314_162),
	.C2V_1 (C2V_162_8),
	.C2V_2 (C2V_162_80),
	.C2V_3 (C2V_162_120),
	.C2V_4 (C2V_162_188),
	.C2V_5 (C2V_162_222),
	.C2V_6 (C2V_162_253),
	.C2V_7 (C2V_162_306),
	.C2V_8 (C2V_162_458),
	.C2V_9 (C2V_162_555),
	.C2V_10 (C2V_162_588),
	.C2V_11 (C2V_162_792),
	.C2V_12 (C2V_162_820),
	.C2V_13 (C2V_162_901),
	.C2V_14 (C2V_162_915),
	.C2V_15 (C2V_162_998),
	.C2V_16 (C2V_162_1017),
	.C2V_17 (C2V_162_1081),
	.C2V_18 (C2V_162_1131),
	.C2V_19 (C2V_162_1313),
	.C2V_20 (C2V_162_1314),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU163 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_32_163),
	.V2C_2 (V2C_68_163),
	.V2C_3 (V2C_136_163),
	.V2C_4 (V2C_149_163),
	.V2C_5 (V2C_211_163),
	.V2C_6 (V2C_254_163),
	.V2C_7 (V2C_354_163),
	.V2C_8 (V2C_408_163),
	.V2C_9 (V2C_505_163),
	.V2C_10 (V2C_741_163),
	.V2C_11 (V2C_789_163),
	.V2C_12 (V2C_837_163),
	.V2C_13 (V2C_878_163),
	.V2C_14 (V2C_919_163),
	.V2C_15 (V2C_1001_163),
	.V2C_16 (V2C_1040_163),
	.V2C_17 (V2C_1066_163),
	.V2C_18 (V2C_1125_163),
	.V2C_19 (V2C_1314_163),
	.V2C_20 (V2C_1315_163),
	.C2V_1 (C2V_163_32),
	.C2V_2 (C2V_163_68),
	.C2V_3 (C2V_163_136),
	.C2V_4 (C2V_163_149),
	.C2V_5 (C2V_163_211),
	.C2V_6 (C2V_163_254),
	.C2V_7 (C2V_163_354),
	.C2V_8 (C2V_163_408),
	.C2V_9 (C2V_163_505),
	.C2V_10 (C2V_163_741),
	.C2V_11 (C2V_163_789),
	.C2V_12 (C2V_163_837),
	.C2V_13 (C2V_163_878),
	.C2V_14 (C2V_163_919),
	.C2V_15 (C2V_163_1001),
	.C2V_16 (C2V_163_1040),
	.C2V_17 (C2V_163_1066),
	.C2V_18 (C2V_163_1125),
	.C2V_19 (C2V_163_1314),
	.C2V_20 (C2V_163_1315),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU164 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_41_164),
	.V2C_2 (V2C_90_164),
	.V2C_3 (V2C_98_164),
	.V2C_4 (V2C_146_164),
	.V2C_5 (V2C_223_164),
	.V2C_6 (V2C_244_164),
	.V2C_7 (V2C_295_164),
	.V2C_8 (V2C_402_164),
	.V2C_9 (V2C_491_164),
	.V2C_10 (V2C_651_164),
	.V2C_11 (V2C_712_164),
	.V2C_12 (V2C_832_164),
	.V2C_13 (V2C_874_164),
	.V2C_14 (V2C_937_164),
	.V2C_15 (V2C_968_164),
	.V2C_16 (V2C_1048_164),
	.V2C_17 (V2C_1067_164),
	.V2C_18 (V2C_1146_164),
	.V2C_19 (V2C_1315_164),
	.V2C_20 (V2C_1316_164),
	.C2V_1 (C2V_164_41),
	.C2V_2 (C2V_164_90),
	.C2V_3 (C2V_164_98),
	.C2V_4 (C2V_164_146),
	.C2V_5 (C2V_164_223),
	.C2V_6 (C2V_164_244),
	.C2V_7 (C2V_164_295),
	.C2V_8 (C2V_164_402),
	.C2V_9 (C2V_164_491),
	.C2V_10 (C2V_164_651),
	.C2V_11 (C2V_164_712),
	.C2V_12 (C2V_164_832),
	.C2V_13 (C2V_164_874),
	.C2V_14 (C2V_164_937),
	.C2V_15 (C2V_164_968),
	.C2V_16 (C2V_164_1048),
	.C2V_17 (C2V_164_1067),
	.C2V_18 (C2V_164_1146),
	.C2V_19 (C2V_164_1315),
	.C2V_20 (C2V_164_1316),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU165 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_36_165),
	.V2C_2 (V2C_63_165),
	.V2C_3 (V2C_128_165),
	.V2C_4 (V2C_162_165),
	.V2C_5 (V2C_228_165),
	.V2C_6 (V2C_247_165),
	.V2C_7 (V2C_344_165),
	.V2C_8 (V2C_399_165),
	.V2C_9 (V2C_558_165),
	.V2C_10 (V2C_615_165),
	.V2C_11 (V2C_643_165),
	.V2C_12 (V2C_747_165),
	.V2C_13 (V2C_878_165),
	.V2C_14 (V2C_922_165),
	.V2C_15 (V2C_995_165),
	.V2C_16 (V2C_1055_165),
	.V2C_17 (V2C_1085_165),
	.V2C_18 (V2C_1130_165),
	.V2C_19 (V2C_1316_165),
	.V2C_20 (V2C_1317_165),
	.C2V_1 (C2V_165_36),
	.C2V_2 (C2V_165_63),
	.C2V_3 (C2V_165_128),
	.C2V_4 (C2V_165_162),
	.C2V_5 (C2V_165_228),
	.C2V_6 (C2V_165_247),
	.C2V_7 (C2V_165_344),
	.C2V_8 (C2V_165_399),
	.C2V_9 (C2V_165_558),
	.C2V_10 (C2V_165_615),
	.C2V_11 (C2V_165_643),
	.C2V_12 (C2V_165_747),
	.C2V_13 (C2V_165_878),
	.C2V_14 (C2V_165_922),
	.C2V_15 (C2V_165_995),
	.C2V_16 (C2V_165_1055),
	.C2V_17 (C2V_165_1085),
	.C2V_18 (C2V_165_1130),
	.C2V_19 (C2V_165_1316),
	.C2V_20 (C2V_165_1317),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU166 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_7_166),
	.V2C_2 (V2C_66_166),
	.V2C_3 (V2C_105_166),
	.V2C_4 (V2C_161_166),
	.V2C_5 (V2C_226_166),
	.V2C_6 (V2C_280_166),
	.V2C_7 (V2C_456_166),
	.V2C_8 (V2C_496_166),
	.V2C_9 (V2C_532_166),
	.V2C_10 (V2C_594_166),
	.V2C_11 (V2C_667_166),
	.V2C_12 (V2C_713_166),
	.V2C_13 (V2C_882_166),
	.V2C_14 (V2C_954_166),
	.V2C_15 (V2C_990_166),
	.V2C_16 (V2C_1020_166),
	.V2C_17 (V2C_1095_166),
	.V2C_18 (V2C_1111_166),
	.V2C_19 (V2C_1317_166),
	.V2C_20 (V2C_1318_166),
	.C2V_1 (C2V_166_7),
	.C2V_2 (C2V_166_66),
	.C2V_3 (C2V_166_105),
	.C2V_4 (C2V_166_161),
	.C2V_5 (C2V_166_226),
	.C2V_6 (C2V_166_280),
	.C2V_7 (C2V_166_456),
	.C2V_8 (C2V_166_496),
	.C2V_9 (C2V_166_532),
	.C2V_10 (C2V_166_594),
	.C2V_11 (C2V_166_667),
	.C2V_12 (C2V_166_713),
	.C2V_13 (C2V_166_882),
	.C2V_14 (C2V_166_954),
	.C2V_15 (C2V_166_990),
	.C2V_16 (C2V_166_1020),
	.C2V_17 (C2V_166_1095),
	.C2V_18 (C2V_166_1111),
	.C2V_19 (C2V_166_1317),
	.C2V_20 (C2V_166_1318),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU167 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_26_167),
	.V2C_2 (V2C_84_167),
	.V2C_3 (V2C_119_167),
	.V2C_4 (V2C_190_167),
	.V2C_5 (V2C_206_167),
	.V2C_6 (V2C_272_167),
	.V2C_7 (V2C_321_167),
	.V2C_8 (V2C_340_167),
	.V2C_9 (V2C_467_167),
	.V2C_10 (V2C_701_167),
	.V2C_11 (V2C_765_167),
	.V2C_12 (V2C_771_167),
	.V2C_13 (V2C_897_167),
	.V2C_14 (V2C_945_167),
	.V2C_15 (V2C_988_167),
	.V2C_16 (V2C_1040_167),
	.V2C_17 (V2C_1089_167),
	.V2C_18 (V2C_1137_167),
	.V2C_19 (V2C_1318_167),
	.V2C_20 (V2C_1319_167),
	.C2V_1 (C2V_167_26),
	.C2V_2 (C2V_167_84),
	.C2V_3 (C2V_167_119),
	.C2V_4 (C2V_167_190),
	.C2V_5 (C2V_167_206),
	.C2V_6 (C2V_167_272),
	.C2V_7 (C2V_167_321),
	.C2V_8 (C2V_167_340),
	.C2V_9 (C2V_167_467),
	.C2V_10 (C2V_167_701),
	.C2V_11 (C2V_167_765),
	.C2V_12 (C2V_167_771),
	.C2V_13 (C2V_167_897),
	.C2V_14 (C2V_167_945),
	.C2V_15 (C2V_167_988),
	.C2V_16 (C2V_167_1040),
	.C2V_17 (C2V_167_1089),
	.C2V_18 (C2V_167_1137),
	.C2V_19 (C2V_167_1318),
	.C2V_20 (C2V_167_1319),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU168 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_9_168),
	.V2C_2 (V2C_81_168),
	.V2C_3 (V2C_121_168),
	.V2C_4 (V2C_189_168),
	.V2C_5 (V2C_223_168),
	.V2C_6 (V2C_254_168),
	.V2C_7 (V2C_307_168),
	.V2C_8 (V2C_459_168),
	.V2C_9 (V2C_556_168),
	.V2C_10 (V2C_589_168),
	.V2C_11 (V2C_793_168),
	.V2C_12 (V2C_821_168),
	.V2C_13 (V2C_902_168),
	.V2C_14 (V2C_916_168),
	.V2C_15 (V2C_999_168),
	.V2C_16 (V2C_1018_168),
	.V2C_17 (V2C_1082_168),
	.V2C_18 (V2C_1132_168),
	.V2C_19 (V2C_1319_168),
	.V2C_20 (V2C_1320_168),
	.C2V_1 (C2V_168_9),
	.C2V_2 (C2V_168_81),
	.C2V_3 (C2V_168_121),
	.C2V_4 (C2V_168_189),
	.C2V_5 (C2V_168_223),
	.C2V_6 (C2V_168_254),
	.C2V_7 (C2V_168_307),
	.C2V_8 (C2V_168_459),
	.C2V_9 (C2V_168_556),
	.C2V_10 (C2V_168_589),
	.C2V_11 (C2V_168_793),
	.C2V_12 (C2V_168_821),
	.C2V_13 (C2V_168_902),
	.C2V_14 (C2V_168_916),
	.C2V_15 (C2V_168_999),
	.C2V_16 (C2V_168_1018),
	.C2V_17 (C2V_168_1082),
	.C2V_18 (C2V_168_1132),
	.C2V_19 (C2V_168_1319),
	.C2V_20 (C2V_168_1320),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU169 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_33_169),
	.V2C_2 (V2C_69_169),
	.V2C_3 (V2C_137_169),
	.V2C_4 (V2C_150_169),
	.V2C_5 (V2C_212_169),
	.V2C_6 (V2C_255_169),
	.V2C_7 (V2C_355_169),
	.V2C_8 (V2C_409_169),
	.V2C_9 (V2C_506_169),
	.V2C_10 (V2C_742_169),
	.V2C_11 (V2C_790_169),
	.V2C_12 (V2C_838_169),
	.V2C_13 (V2C_879_169),
	.V2C_14 (V2C_920_169),
	.V2C_15 (V2C_1002_169),
	.V2C_16 (V2C_1041_169),
	.V2C_17 (V2C_1067_169),
	.V2C_18 (V2C_1126_169),
	.V2C_19 (V2C_1320_169),
	.V2C_20 (V2C_1321_169),
	.C2V_1 (C2V_169_33),
	.C2V_2 (C2V_169_69),
	.C2V_3 (C2V_169_137),
	.C2V_4 (C2V_169_150),
	.C2V_5 (C2V_169_212),
	.C2V_6 (C2V_169_255),
	.C2V_7 (C2V_169_355),
	.C2V_8 (C2V_169_409),
	.C2V_9 (C2V_169_506),
	.C2V_10 (C2V_169_742),
	.C2V_11 (C2V_169_790),
	.C2V_12 (C2V_169_838),
	.C2V_13 (C2V_169_879),
	.C2V_14 (C2V_169_920),
	.C2V_15 (C2V_169_1002),
	.C2V_16 (C2V_169_1041),
	.C2V_17 (C2V_169_1067),
	.C2V_18 (C2V_169_1126),
	.C2V_19 (C2V_169_1320),
	.C2V_20 (C2V_169_1321),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU170 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_42_170),
	.V2C_2 (V2C_91_170),
	.V2C_3 (V2C_99_170),
	.V2C_4 (V2C_147_170),
	.V2C_5 (V2C_224_170),
	.V2C_6 (V2C_245_170),
	.V2C_7 (V2C_296_170),
	.V2C_8 (V2C_403_170),
	.V2C_9 (V2C_492_170),
	.V2C_10 (V2C_652_170),
	.V2C_11 (V2C_713_170),
	.V2C_12 (V2C_833_170),
	.V2C_13 (V2C_875_170),
	.V2C_14 (V2C_938_170),
	.V2C_15 (V2C_969_170),
	.V2C_16 (V2C_1049_170),
	.V2C_17 (V2C_1068_170),
	.V2C_18 (V2C_1147_170),
	.V2C_19 (V2C_1321_170),
	.V2C_20 (V2C_1322_170),
	.C2V_1 (C2V_170_42),
	.C2V_2 (C2V_170_91),
	.C2V_3 (C2V_170_99),
	.C2V_4 (C2V_170_147),
	.C2V_5 (C2V_170_224),
	.C2V_6 (C2V_170_245),
	.C2V_7 (C2V_170_296),
	.C2V_8 (C2V_170_403),
	.C2V_9 (C2V_170_492),
	.C2V_10 (C2V_170_652),
	.C2V_11 (C2V_170_713),
	.C2V_12 (C2V_170_833),
	.C2V_13 (C2V_170_875),
	.C2V_14 (C2V_170_938),
	.C2V_15 (C2V_170_969),
	.C2V_16 (C2V_170_1049),
	.C2V_17 (C2V_170_1068),
	.C2V_18 (C2V_170_1147),
	.C2V_19 (C2V_170_1321),
	.C2V_20 (C2V_170_1322),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU171 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_37_171),
	.V2C_2 (V2C_64_171),
	.V2C_3 (V2C_129_171),
	.V2C_4 (V2C_163_171),
	.V2C_5 (V2C_229_171),
	.V2C_6 (V2C_248_171),
	.V2C_7 (V2C_345_171),
	.V2C_8 (V2C_400_171),
	.V2C_9 (V2C_559_171),
	.V2C_10 (V2C_616_171),
	.V2C_11 (V2C_644_171),
	.V2C_12 (V2C_748_171),
	.V2C_13 (V2C_879_171),
	.V2C_14 (V2C_923_171),
	.V2C_15 (V2C_996_171),
	.V2C_16 (V2C_1056_171),
	.V2C_17 (V2C_1086_171),
	.V2C_18 (V2C_1131_171),
	.V2C_19 (V2C_1322_171),
	.V2C_20 (V2C_1323_171),
	.C2V_1 (C2V_171_37),
	.C2V_2 (C2V_171_64),
	.C2V_3 (C2V_171_129),
	.C2V_4 (C2V_171_163),
	.C2V_5 (C2V_171_229),
	.C2V_6 (C2V_171_248),
	.C2V_7 (C2V_171_345),
	.C2V_8 (C2V_171_400),
	.C2V_9 (C2V_171_559),
	.C2V_10 (C2V_171_616),
	.C2V_11 (C2V_171_644),
	.C2V_12 (C2V_171_748),
	.C2V_13 (C2V_171_879),
	.C2V_14 (C2V_171_923),
	.C2V_15 (C2V_171_996),
	.C2V_16 (C2V_171_1056),
	.C2V_17 (C2V_171_1086),
	.C2V_18 (C2V_171_1131),
	.C2V_19 (C2V_171_1322),
	.C2V_20 (C2V_171_1323),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU172 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_8_172),
	.V2C_2 (V2C_67_172),
	.V2C_3 (V2C_106_172),
	.V2C_4 (V2C_162_172),
	.V2C_5 (V2C_227_172),
	.V2C_6 (V2C_281_172),
	.V2C_7 (V2C_457_172),
	.V2C_8 (V2C_497_172),
	.V2C_9 (V2C_533_172),
	.V2C_10 (V2C_595_172),
	.V2C_11 (V2C_668_172),
	.V2C_12 (V2C_714_172),
	.V2C_13 (V2C_883_172),
	.V2C_14 (V2C_955_172),
	.V2C_15 (V2C_991_172),
	.V2C_16 (V2C_1021_172),
	.V2C_17 (V2C_1096_172),
	.V2C_18 (V2C_1112_172),
	.V2C_19 (V2C_1323_172),
	.V2C_20 (V2C_1324_172),
	.C2V_1 (C2V_172_8),
	.C2V_2 (C2V_172_67),
	.C2V_3 (C2V_172_106),
	.C2V_4 (C2V_172_162),
	.C2V_5 (C2V_172_227),
	.C2V_6 (C2V_172_281),
	.C2V_7 (C2V_172_457),
	.C2V_8 (C2V_172_497),
	.C2V_9 (C2V_172_533),
	.C2V_10 (C2V_172_595),
	.C2V_11 (C2V_172_668),
	.C2V_12 (C2V_172_714),
	.C2V_13 (C2V_172_883),
	.C2V_14 (C2V_172_955),
	.C2V_15 (C2V_172_991),
	.C2V_16 (C2V_172_1021),
	.C2V_17 (C2V_172_1096),
	.C2V_18 (C2V_172_1112),
	.C2V_19 (C2V_172_1323),
	.C2V_20 (C2V_172_1324),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU173 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_27_173),
	.V2C_2 (V2C_85_173),
	.V2C_3 (V2C_120_173),
	.V2C_4 (V2C_191_173),
	.V2C_5 (V2C_207_173),
	.V2C_6 (V2C_273_173),
	.V2C_7 (V2C_322_173),
	.V2C_8 (V2C_341_173),
	.V2C_9 (V2C_468_173),
	.V2C_10 (V2C_702_173),
	.V2C_11 (V2C_766_173),
	.V2C_12 (V2C_772_173),
	.V2C_13 (V2C_898_173),
	.V2C_14 (V2C_946_173),
	.V2C_15 (V2C_989_173),
	.V2C_16 (V2C_1041_173),
	.V2C_17 (V2C_1090_173),
	.V2C_18 (V2C_1138_173),
	.V2C_19 (V2C_1324_173),
	.V2C_20 (V2C_1325_173),
	.C2V_1 (C2V_173_27),
	.C2V_2 (C2V_173_85),
	.C2V_3 (C2V_173_120),
	.C2V_4 (C2V_173_191),
	.C2V_5 (C2V_173_207),
	.C2V_6 (C2V_173_273),
	.C2V_7 (C2V_173_322),
	.C2V_8 (C2V_173_341),
	.C2V_9 (C2V_173_468),
	.C2V_10 (C2V_173_702),
	.C2V_11 (C2V_173_766),
	.C2V_12 (C2V_173_772),
	.C2V_13 (C2V_173_898),
	.C2V_14 (C2V_173_946),
	.C2V_15 (C2V_173_989),
	.C2V_16 (C2V_173_1041),
	.C2V_17 (C2V_173_1090),
	.C2V_18 (C2V_173_1138),
	.C2V_19 (C2V_173_1324),
	.C2V_20 (C2V_173_1325),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU174 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_10_174),
	.V2C_2 (V2C_82_174),
	.V2C_3 (V2C_122_174),
	.V2C_4 (V2C_190_174),
	.V2C_5 (V2C_224_174),
	.V2C_6 (V2C_255_174),
	.V2C_7 (V2C_308_174),
	.V2C_8 (V2C_460_174),
	.V2C_9 (V2C_557_174),
	.V2C_10 (V2C_590_174),
	.V2C_11 (V2C_794_174),
	.V2C_12 (V2C_822_174),
	.V2C_13 (V2C_903_174),
	.V2C_14 (V2C_917_174),
	.V2C_15 (V2C_1000_174),
	.V2C_16 (V2C_1019_174),
	.V2C_17 (V2C_1083_174),
	.V2C_18 (V2C_1133_174),
	.V2C_19 (V2C_1325_174),
	.V2C_20 (V2C_1326_174),
	.C2V_1 (C2V_174_10),
	.C2V_2 (C2V_174_82),
	.C2V_3 (C2V_174_122),
	.C2V_4 (C2V_174_190),
	.C2V_5 (C2V_174_224),
	.C2V_6 (C2V_174_255),
	.C2V_7 (C2V_174_308),
	.C2V_8 (C2V_174_460),
	.C2V_9 (C2V_174_557),
	.C2V_10 (C2V_174_590),
	.C2V_11 (C2V_174_794),
	.C2V_12 (C2V_174_822),
	.C2V_13 (C2V_174_903),
	.C2V_14 (C2V_174_917),
	.C2V_15 (C2V_174_1000),
	.C2V_16 (C2V_174_1019),
	.C2V_17 (C2V_174_1083),
	.C2V_18 (C2V_174_1133),
	.C2V_19 (C2V_174_1325),
	.C2V_20 (C2V_174_1326),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU175 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_34_175),
	.V2C_2 (V2C_70_175),
	.V2C_3 (V2C_138_175),
	.V2C_4 (V2C_151_175),
	.V2C_5 (V2C_213_175),
	.V2C_6 (V2C_256_175),
	.V2C_7 (V2C_356_175),
	.V2C_8 (V2C_410_175),
	.V2C_9 (V2C_507_175),
	.V2C_10 (V2C_743_175),
	.V2C_11 (V2C_791_175),
	.V2C_12 (V2C_839_175),
	.V2C_13 (V2C_880_175),
	.V2C_14 (V2C_921_175),
	.V2C_15 (V2C_1003_175),
	.V2C_16 (V2C_1042_175),
	.V2C_17 (V2C_1068_175),
	.V2C_18 (V2C_1127_175),
	.V2C_19 (V2C_1326_175),
	.V2C_20 (V2C_1327_175),
	.C2V_1 (C2V_175_34),
	.C2V_2 (C2V_175_70),
	.C2V_3 (C2V_175_138),
	.C2V_4 (C2V_175_151),
	.C2V_5 (C2V_175_213),
	.C2V_6 (C2V_175_256),
	.C2V_7 (C2V_175_356),
	.C2V_8 (C2V_175_410),
	.C2V_9 (C2V_175_507),
	.C2V_10 (C2V_175_743),
	.C2V_11 (C2V_175_791),
	.C2V_12 (C2V_175_839),
	.C2V_13 (C2V_175_880),
	.C2V_14 (C2V_175_921),
	.C2V_15 (C2V_175_1003),
	.C2V_16 (C2V_175_1042),
	.C2V_17 (C2V_175_1068),
	.C2V_18 (C2V_175_1127),
	.C2V_19 (C2V_175_1326),
	.C2V_20 (C2V_175_1327),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU176 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_43_176),
	.V2C_2 (V2C_92_176),
	.V2C_3 (V2C_100_176),
	.V2C_4 (V2C_148_176),
	.V2C_5 (V2C_225_176),
	.V2C_6 (V2C_246_176),
	.V2C_7 (V2C_297_176),
	.V2C_8 (V2C_404_176),
	.V2C_9 (V2C_493_176),
	.V2C_10 (V2C_653_176),
	.V2C_11 (V2C_714_176),
	.V2C_12 (V2C_834_176),
	.V2C_13 (V2C_876_176),
	.V2C_14 (V2C_939_176),
	.V2C_15 (V2C_970_176),
	.V2C_16 (V2C_1050_176),
	.V2C_17 (V2C_1069_176),
	.V2C_18 (V2C_1148_176),
	.V2C_19 (V2C_1327_176),
	.V2C_20 (V2C_1328_176),
	.C2V_1 (C2V_176_43),
	.C2V_2 (C2V_176_92),
	.C2V_3 (C2V_176_100),
	.C2V_4 (C2V_176_148),
	.C2V_5 (C2V_176_225),
	.C2V_6 (C2V_176_246),
	.C2V_7 (C2V_176_297),
	.C2V_8 (C2V_176_404),
	.C2V_9 (C2V_176_493),
	.C2V_10 (C2V_176_653),
	.C2V_11 (C2V_176_714),
	.C2V_12 (C2V_176_834),
	.C2V_13 (C2V_176_876),
	.C2V_14 (C2V_176_939),
	.C2V_15 (C2V_176_970),
	.C2V_16 (C2V_176_1050),
	.C2V_17 (C2V_176_1069),
	.C2V_18 (C2V_176_1148),
	.C2V_19 (C2V_176_1327),
	.C2V_20 (C2V_176_1328),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU177 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_38_177),
	.V2C_2 (V2C_65_177),
	.V2C_3 (V2C_130_177),
	.V2C_4 (V2C_164_177),
	.V2C_5 (V2C_230_177),
	.V2C_6 (V2C_249_177),
	.V2C_7 (V2C_346_177),
	.V2C_8 (V2C_401_177),
	.V2C_9 (V2C_560_177),
	.V2C_10 (V2C_617_177),
	.V2C_11 (V2C_645_177),
	.V2C_12 (V2C_749_177),
	.V2C_13 (V2C_880_177),
	.V2C_14 (V2C_924_177),
	.V2C_15 (V2C_997_177),
	.V2C_16 (V2C_1009_177),
	.V2C_17 (V2C_1087_177),
	.V2C_18 (V2C_1132_177),
	.V2C_19 (V2C_1328_177),
	.V2C_20 (V2C_1329_177),
	.C2V_1 (C2V_177_38),
	.C2V_2 (C2V_177_65),
	.C2V_3 (C2V_177_130),
	.C2V_4 (C2V_177_164),
	.C2V_5 (C2V_177_230),
	.C2V_6 (C2V_177_249),
	.C2V_7 (C2V_177_346),
	.C2V_8 (C2V_177_401),
	.C2V_9 (C2V_177_560),
	.C2V_10 (C2V_177_617),
	.C2V_11 (C2V_177_645),
	.C2V_12 (C2V_177_749),
	.C2V_13 (C2V_177_880),
	.C2V_14 (C2V_177_924),
	.C2V_15 (C2V_177_997),
	.C2V_16 (C2V_177_1009),
	.C2V_17 (C2V_177_1087),
	.C2V_18 (C2V_177_1132),
	.C2V_19 (C2V_177_1328),
	.C2V_20 (C2V_177_1329),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU178 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_9_178),
	.V2C_2 (V2C_68_178),
	.V2C_3 (V2C_107_178),
	.V2C_4 (V2C_163_178),
	.V2C_5 (V2C_228_178),
	.V2C_6 (V2C_282_178),
	.V2C_7 (V2C_458_178),
	.V2C_8 (V2C_498_178),
	.V2C_9 (V2C_534_178),
	.V2C_10 (V2C_596_178),
	.V2C_11 (V2C_669_178),
	.V2C_12 (V2C_715_178),
	.V2C_13 (V2C_884_178),
	.V2C_14 (V2C_956_178),
	.V2C_15 (V2C_992_178),
	.V2C_16 (V2C_1022_178),
	.V2C_17 (V2C_1097_178),
	.V2C_18 (V2C_1113_178),
	.V2C_19 (V2C_1329_178),
	.V2C_20 (V2C_1330_178),
	.C2V_1 (C2V_178_9),
	.C2V_2 (C2V_178_68),
	.C2V_3 (C2V_178_107),
	.C2V_4 (C2V_178_163),
	.C2V_5 (C2V_178_228),
	.C2V_6 (C2V_178_282),
	.C2V_7 (C2V_178_458),
	.C2V_8 (C2V_178_498),
	.C2V_9 (C2V_178_534),
	.C2V_10 (C2V_178_596),
	.C2V_11 (C2V_178_669),
	.C2V_12 (C2V_178_715),
	.C2V_13 (C2V_178_884),
	.C2V_14 (C2V_178_956),
	.C2V_15 (C2V_178_992),
	.C2V_16 (C2V_178_1022),
	.C2V_17 (C2V_178_1097),
	.C2V_18 (C2V_178_1113),
	.C2V_19 (C2V_178_1329),
	.C2V_20 (C2V_178_1330),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU179 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_28_179),
	.V2C_2 (V2C_86_179),
	.V2C_3 (V2C_121_179),
	.V2C_4 (V2C_192_179),
	.V2C_5 (V2C_208_179),
	.V2C_6 (V2C_274_179),
	.V2C_7 (V2C_323_179),
	.V2C_8 (V2C_342_179),
	.V2C_9 (V2C_469_179),
	.V2C_10 (V2C_703_179),
	.V2C_11 (V2C_767_179),
	.V2C_12 (V2C_773_179),
	.V2C_13 (V2C_899_179),
	.V2C_14 (V2C_947_179),
	.V2C_15 (V2C_990_179),
	.V2C_16 (V2C_1042_179),
	.V2C_17 (V2C_1091_179),
	.V2C_18 (V2C_1139_179),
	.V2C_19 (V2C_1330_179),
	.V2C_20 (V2C_1331_179),
	.C2V_1 (C2V_179_28),
	.C2V_2 (C2V_179_86),
	.C2V_3 (C2V_179_121),
	.C2V_4 (C2V_179_192),
	.C2V_5 (C2V_179_208),
	.C2V_6 (C2V_179_274),
	.C2V_7 (C2V_179_323),
	.C2V_8 (C2V_179_342),
	.C2V_9 (C2V_179_469),
	.C2V_10 (C2V_179_703),
	.C2V_11 (C2V_179_767),
	.C2V_12 (C2V_179_773),
	.C2V_13 (C2V_179_899),
	.C2V_14 (C2V_179_947),
	.C2V_15 (C2V_179_990),
	.C2V_16 (C2V_179_1042),
	.C2V_17 (C2V_179_1091),
	.C2V_18 (C2V_179_1139),
	.C2V_19 (C2V_179_1330),
	.C2V_20 (C2V_179_1331),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU180 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_11_180),
	.V2C_2 (V2C_83_180),
	.V2C_3 (V2C_123_180),
	.V2C_4 (V2C_191_180),
	.V2C_5 (V2C_225_180),
	.V2C_6 (V2C_256_180),
	.V2C_7 (V2C_309_180),
	.V2C_8 (V2C_461_180),
	.V2C_9 (V2C_558_180),
	.V2C_10 (V2C_591_180),
	.V2C_11 (V2C_795_180),
	.V2C_12 (V2C_823_180),
	.V2C_13 (V2C_904_180),
	.V2C_14 (V2C_918_180),
	.V2C_15 (V2C_1001_180),
	.V2C_16 (V2C_1020_180),
	.V2C_17 (V2C_1084_180),
	.V2C_18 (V2C_1134_180),
	.V2C_19 (V2C_1331_180),
	.V2C_20 (V2C_1332_180),
	.C2V_1 (C2V_180_11),
	.C2V_2 (C2V_180_83),
	.C2V_3 (C2V_180_123),
	.C2V_4 (C2V_180_191),
	.C2V_5 (C2V_180_225),
	.C2V_6 (C2V_180_256),
	.C2V_7 (C2V_180_309),
	.C2V_8 (C2V_180_461),
	.C2V_9 (C2V_180_558),
	.C2V_10 (C2V_180_591),
	.C2V_11 (C2V_180_795),
	.C2V_12 (C2V_180_823),
	.C2V_13 (C2V_180_904),
	.C2V_14 (C2V_180_918),
	.C2V_15 (C2V_180_1001),
	.C2V_16 (C2V_180_1020),
	.C2V_17 (C2V_180_1084),
	.C2V_18 (C2V_180_1134),
	.C2V_19 (C2V_180_1331),
	.C2V_20 (C2V_180_1332),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU181 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_35_181),
	.V2C_2 (V2C_71_181),
	.V2C_3 (V2C_139_181),
	.V2C_4 (V2C_152_181),
	.V2C_5 (V2C_214_181),
	.V2C_6 (V2C_257_181),
	.V2C_7 (V2C_357_181),
	.V2C_8 (V2C_411_181),
	.V2C_9 (V2C_508_181),
	.V2C_10 (V2C_744_181),
	.V2C_11 (V2C_792_181),
	.V2C_12 (V2C_840_181),
	.V2C_13 (V2C_881_181),
	.V2C_14 (V2C_922_181),
	.V2C_15 (V2C_1004_181),
	.V2C_16 (V2C_1043_181),
	.V2C_17 (V2C_1069_181),
	.V2C_18 (V2C_1128_181),
	.V2C_19 (V2C_1332_181),
	.V2C_20 (V2C_1333_181),
	.C2V_1 (C2V_181_35),
	.C2V_2 (C2V_181_71),
	.C2V_3 (C2V_181_139),
	.C2V_4 (C2V_181_152),
	.C2V_5 (C2V_181_214),
	.C2V_6 (C2V_181_257),
	.C2V_7 (C2V_181_357),
	.C2V_8 (C2V_181_411),
	.C2V_9 (C2V_181_508),
	.C2V_10 (C2V_181_744),
	.C2V_11 (C2V_181_792),
	.C2V_12 (C2V_181_840),
	.C2V_13 (C2V_181_881),
	.C2V_14 (C2V_181_922),
	.C2V_15 (C2V_181_1004),
	.C2V_16 (C2V_181_1043),
	.C2V_17 (C2V_181_1069),
	.C2V_18 (C2V_181_1128),
	.C2V_19 (C2V_181_1332),
	.C2V_20 (C2V_181_1333),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU182 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_44_182),
	.V2C_2 (V2C_93_182),
	.V2C_3 (V2C_101_182),
	.V2C_4 (V2C_149_182),
	.V2C_5 (V2C_226_182),
	.V2C_6 (V2C_247_182),
	.V2C_7 (V2C_298_182),
	.V2C_8 (V2C_405_182),
	.V2C_9 (V2C_494_182),
	.V2C_10 (V2C_654_182),
	.V2C_11 (V2C_715_182),
	.V2C_12 (V2C_835_182),
	.V2C_13 (V2C_877_182),
	.V2C_14 (V2C_940_182),
	.V2C_15 (V2C_971_182),
	.V2C_16 (V2C_1051_182),
	.V2C_17 (V2C_1070_182),
	.V2C_18 (V2C_1149_182),
	.V2C_19 (V2C_1333_182),
	.V2C_20 (V2C_1334_182),
	.C2V_1 (C2V_182_44),
	.C2V_2 (C2V_182_93),
	.C2V_3 (C2V_182_101),
	.C2V_4 (C2V_182_149),
	.C2V_5 (C2V_182_226),
	.C2V_6 (C2V_182_247),
	.C2V_7 (C2V_182_298),
	.C2V_8 (C2V_182_405),
	.C2V_9 (C2V_182_494),
	.C2V_10 (C2V_182_654),
	.C2V_11 (C2V_182_715),
	.C2V_12 (C2V_182_835),
	.C2V_13 (C2V_182_877),
	.C2V_14 (C2V_182_940),
	.C2V_15 (C2V_182_971),
	.C2V_16 (C2V_182_1051),
	.C2V_17 (C2V_182_1070),
	.C2V_18 (C2V_182_1149),
	.C2V_19 (C2V_182_1333),
	.C2V_20 (C2V_182_1334),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU183 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_39_183),
	.V2C_2 (V2C_66_183),
	.V2C_3 (V2C_131_183),
	.V2C_4 (V2C_165_183),
	.V2C_5 (V2C_231_183),
	.V2C_6 (V2C_250_183),
	.V2C_7 (V2C_347_183),
	.V2C_8 (V2C_402_183),
	.V2C_9 (V2C_561_183),
	.V2C_10 (V2C_618_183),
	.V2C_11 (V2C_646_183),
	.V2C_12 (V2C_750_183),
	.V2C_13 (V2C_881_183),
	.V2C_14 (V2C_925_183),
	.V2C_15 (V2C_998_183),
	.V2C_16 (V2C_1010_183),
	.V2C_17 (V2C_1088_183),
	.V2C_18 (V2C_1133_183),
	.V2C_19 (V2C_1334_183),
	.V2C_20 (V2C_1335_183),
	.C2V_1 (C2V_183_39),
	.C2V_2 (C2V_183_66),
	.C2V_3 (C2V_183_131),
	.C2V_4 (C2V_183_165),
	.C2V_5 (C2V_183_231),
	.C2V_6 (C2V_183_250),
	.C2V_7 (C2V_183_347),
	.C2V_8 (C2V_183_402),
	.C2V_9 (C2V_183_561),
	.C2V_10 (C2V_183_618),
	.C2V_11 (C2V_183_646),
	.C2V_12 (C2V_183_750),
	.C2V_13 (C2V_183_881),
	.C2V_14 (C2V_183_925),
	.C2V_15 (C2V_183_998),
	.C2V_16 (C2V_183_1010),
	.C2V_17 (C2V_183_1088),
	.C2V_18 (C2V_183_1133),
	.C2V_19 (C2V_183_1334),
	.C2V_20 (C2V_183_1335),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU184 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_10_184),
	.V2C_2 (V2C_69_184),
	.V2C_3 (V2C_108_184),
	.V2C_4 (V2C_164_184),
	.V2C_5 (V2C_229_184),
	.V2C_6 (V2C_283_184),
	.V2C_7 (V2C_459_184),
	.V2C_8 (V2C_499_184),
	.V2C_9 (V2C_535_184),
	.V2C_10 (V2C_597_184),
	.V2C_11 (V2C_670_184),
	.V2C_12 (V2C_716_184),
	.V2C_13 (V2C_885_184),
	.V2C_14 (V2C_957_184),
	.V2C_15 (V2C_993_184),
	.V2C_16 (V2C_1023_184),
	.V2C_17 (V2C_1098_184),
	.V2C_18 (V2C_1114_184),
	.V2C_19 (V2C_1335_184),
	.V2C_20 (V2C_1336_184),
	.C2V_1 (C2V_184_10),
	.C2V_2 (C2V_184_69),
	.C2V_3 (C2V_184_108),
	.C2V_4 (C2V_184_164),
	.C2V_5 (C2V_184_229),
	.C2V_6 (C2V_184_283),
	.C2V_7 (C2V_184_459),
	.C2V_8 (C2V_184_499),
	.C2V_9 (C2V_184_535),
	.C2V_10 (C2V_184_597),
	.C2V_11 (C2V_184_670),
	.C2V_12 (C2V_184_716),
	.C2V_13 (C2V_184_885),
	.C2V_14 (C2V_184_957),
	.C2V_15 (C2V_184_993),
	.C2V_16 (C2V_184_1023),
	.C2V_17 (C2V_184_1098),
	.C2V_18 (C2V_184_1114),
	.C2V_19 (C2V_184_1335),
	.C2V_20 (C2V_184_1336),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU185 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_29_185),
	.V2C_2 (V2C_87_185),
	.V2C_3 (V2C_122_185),
	.V2C_4 (V2C_145_185),
	.V2C_5 (V2C_209_185),
	.V2C_6 (V2C_275_185),
	.V2C_7 (V2C_324_185),
	.V2C_8 (V2C_343_185),
	.V2C_9 (V2C_470_185),
	.V2C_10 (V2C_704_185),
	.V2C_11 (V2C_768_185),
	.V2C_12 (V2C_774_185),
	.V2C_13 (V2C_900_185),
	.V2C_14 (V2C_948_185),
	.V2C_15 (V2C_991_185),
	.V2C_16 (V2C_1043_185),
	.V2C_17 (V2C_1092_185),
	.V2C_18 (V2C_1140_185),
	.V2C_19 (V2C_1336_185),
	.V2C_20 (V2C_1337_185),
	.C2V_1 (C2V_185_29),
	.C2V_2 (C2V_185_87),
	.C2V_3 (C2V_185_122),
	.C2V_4 (C2V_185_145),
	.C2V_5 (C2V_185_209),
	.C2V_6 (C2V_185_275),
	.C2V_7 (C2V_185_324),
	.C2V_8 (C2V_185_343),
	.C2V_9 (C2V_185_470),
	.C2V_10 (C2V_185_704),
	.C2V_11 (C2V_185_768),
	.C2V_12 (C2V_185_774),
	.C2V_13 (C2V_185_900),
	.C2V_14 (C2V_185_948),
	.C2V_15 (C2V_185_991),
	.C2V_16 (C2V_185_1043),
	.C2V_17 (C2V_185_1092),
	.C2V_18 (C2V_185_1140),
	.C2V_19 (C2V_185_1336),
	.C2V_20 (C2V_185_1337),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU186 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_12_186),
	.V2C_2 (V2C_84_186),
	.V2C_3 (V2C_124_186),
	.V2C_4 (V2C_192_186),
	.V2C_5 (V2C_226_186),
	.V2C_6 (V2C_257_186),
	.V2C_7 (V2C_310_186),
	.V2C_8 (V2C_462_186),
	.V2C_9 (V2C_559_186),
	.V2C_10 (V2C_592_186),
	.V2C_11 (V2C_796_186),
	.V2C_12 (V2C_824_186),
	.V2C_13 (V2C_905_186),
	.V2C_14 (V2C_919_186),
	.V2C_15 (V2C_1002_186),
	.V2C_16 (V2C_1021_186),
	.V2C_17 (V2C_1085_186),
	.V2C_18 (V2C_1135_186),
	.V2C_19 (V2C_1337_186),
	.V2C_20 (V2C_1338_186),
	.C2V_1 (C2V_186_12),
	.C2V_2 (C2V_186_84),
	.C2V_3 (C2V_186_124),
	.C2V_4 (C2V_186_192),
	.C2V_5 (C2V_186_226),
	.C2V_6 (C2V_186_257),
	.C2V_7 (C2V_186_310),
	.C2V_8 (C2V_186_462),
	.C2V_9 (C2V_186_559),
	.C2V_10 (C2V_186_592),
	.C2V_11 (C2V_186_796),
	.C2V_12 (C2V_186_824),
	.C2V_13 (C2V_186_905),
	.C2V_14 (C2V_186_919),
	.C2V_15 (C2V_186_1002),
	.C2V_16 (C2V_186_1021),
	.C2V_17 (C2V_186_1085),
	.C2V_18 (C2V_186_1135),
	.C2V_19 (C2V_186_1337),
	.C2V_20 (C2V_186_1338),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU187 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_36_187),
	.V2C_2 (V2C_72_187),
	.V2C_3 (V2C_140_187),
	.V2C_4 (V2C_153_187),
	.V2C_5 (V2C_215_187),
	.V2C_6 (V2C_258_187),
	.V2C_7 (V2C_358_187),
	.V2C_8 (V2C_412_187),
	.V2C_9 (V2C_509_187),
	.V2C_10 (V2C_745_187),
	.V2C_11 (V2C_793_187),
	.V2C_12 (V2C_841_187),
	.V2C_13 (V2C_882_187),
	.V2C_14 (V2C_923_187),
	.V2C_15 (V2C_1005_187),
	.V2C_16 (V2C_1044_187),
	.V2C_17 (V2C_1070_187),
	.V2C_18 (V2C_1129_187),
	.V2C_19 (V2C_1338_187),
	.V2C_20 (V2C_1339_187),
	.C2V_1 (C2V_187_36),
	.C2V_2 (C2V_187_72),
	.C2V_3 (C2V_187_140),
	.C2V_4 (C2V_187_153),
	.C2V_5 (C2V_187_215),
	.C2V_6 (C2V_187_258),
	.C2V_7 (C2V_187_358),
	.C2V_8 (C2V_187_412),
	.C2V_9 (C2V_187_509),
	.C2V_10 (C2V_187_745),
	.C2V_11 (C2V_187_793),
	.C2V_12 (C2V_187_841),
	.C2V_13 (C2V_187_882),
	.C2V_14 (C2V_187_923),
	.C2V_15 (C2V_187_1005),
	.C2V_16 (C2V_187_1044),
	.C2V_17 (C2V_187_1070),
	.C2V_18 (C2V_187_1129),
	.C2V_19 (C2V_187_1338),
	.C2V_20 (C2V_187_1339),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU188 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_45_188),
	.V2C_2 (V2C_94_188),
	.V2C_3 (V2C_102_188),
	.V2C_4 (V2C_150_188),
	.V2C_5 (V2C_227_188),
	.V2C_6 (V2C_248_188),
	.V2C_7 (V2C_299_188),
	.V2C_8 (V2C_406_188),
	.V2C_9 (V2C_495_188),
	.V2C_10 (V2C_655_188),
	.V2C_11 (V2C_716_188),
	.V2C_12 (V2C_836_188),
	.V2C_13 (V2C_878_188),
	.V2C_14 (V2C_941_188),
	.V2C_15 (V2C_972_188),
	.V2C_16 (V2C_1052_188),
	.V2C_17 (V2C_1071_188),
	.V2C_18 (V2C_1150_188),
	.V2C_19 (V2C_1339_188),
	.V2C_20 (V2C_1340_188),
	.C2V_1 (C2V_188_45),
	.C2V_2 (C2V_188_94),
	.C2V_3 (C2V_188_102),
	.C2V_4 (C2V_188_150),
	.C2V_5 (C2V_188_227),
	.C2V_6 (C2V_188_248),
	.C2V_7 (C2V_188_299),
	.C2V_8 (C2V_188_406),
	.C2V_9 (C2V_188_495),
	.C2V_10 (C2V_188_655),
	.C2V_11 (C2V_188_716),
	.C2V_12 (C2V_188_836),
	.C2V_13 (C2V_188_878),
	.C2V_14 (C2V_188_941),
	.C2V_15 (C2V_188_972),
	.C2V_16 (C2V_188_1052),
	.C2V_17 (C2V_188_1071),
	.C2V_18 (C2V_188_1150),
	.C2V_19 (C2V_188_1339),
	.C2V_20 (C2V_188_1340),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU189 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_40_189),
	.V2C_2 (V2C_67_189),
	.V2C_3 (V2C_132_189),
	.V2C_4 (V2C_166_189),
	.V2C_5 (V2C_232_189),
	.V2C_6 (V2C_251_189),
	.V2C_7 (V2C_348_189),
	.V2C_8 (V2C_403_189),
	.V2C_9 (V2C_562_189),
	.V2C_10 (V2C_619_189),
	.V2C_11 (V2C_647_189),
	.V2C_12 (V2C_751_189),
	.V2C_13 (V2C_882_189),
	.V2C_14 (V2C_926_189),
	.V2C_15 (V2C_999_189),
	.V2C_16 (V2C_1011_189),
	.V2C_17 (V2C_1089_189),
	.V2C_18 (V2C_1134_189),
	.V2C_19 (V2C_1340_189),
	.V2C_20 (V2C_1341_189),
	.C2V_1 (C2V_189_40),
	.C2V_2 (C2V_189_67),
	.C2V_3 (C2V_189_132),
	.C2V_4 (C2V_189_166),
	.C2V_5 (C2V_189_232),
	.C2V_6 (C2V_189_251),
	.C2V_7 (C2V_189_348),
	.C2V_8 (C2V_189_403),
	.C2V_9 (C2V_189_562),
	.C2V_10 (C2V_189_619),
	.C2V_11 (C2V_189_647),
	.C2V_12 (C2V_189_751),
	.C2V_13 (C2V_189_882),
	.C2V_14 (C2V_189_926),
	.C2V_15 (C2V_189_999),
	.C2V_16 (C2V_189_1011),
	.C2V_17 (C2V_189_1089),
	.C2V_18 (C2V_189_1134),
	.C2V_19 (C2V_189_1340),
	.C2V_20 (C2V_189_1341),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU190 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_11_190),
	.V2C_2 (V2C_70_190),
	.V2C_3 (V2C_109_190),
	.V2C_4 (V2C_165_190),
	.V2C_5 (V2C_230_190),
	.V2C_6 (V2C_284_190),
	.V2C_7 (V2C_460_190),
	.V2C_8 (V2C_500_190),
	.V2C_9 (V2C_536_190),
	.V2C_10 (V2C_598_190),
	.V2C_11 (V2C_671_190),
	.V2C_12 (V2C_717_190),
	.V2C_13 (V2C_886_190),
	.V2C_14 (V2C_958_190),
	.V2C_15 (V2C_994_190),
	.V2C_16 (V2C_1024_190),
	.V2C_17 (V2C_1099_190),
	.V2C_18 (V2C_1115_190),
	.V2C_19 (V2C_1341_190),
	.V2C_20 (V2C_1342_190),
	.C2V_1 (C2V_190_11),
	.C2V_2 (C2V_190_70),
	.C2V_3 (C2V_190_109),
	.C2V_4 (C2V_190_165),
	.C2V_5 (C2V_190_230),
	.C2V_6 (C2V_190_284),
	.C2V_7 (C2V_190_460),
	.C2V_8 (C2V_190_500),
	.C2V_9 (C2V_190_536),
	.C2V_10 (C2V_190_598),
	.C2V_11 (C2V_190_671),
	.C2V_12 (C2V_190_717),
	.C2V_13 (C2V_190_886),
	.C2V_14 (C2V_190_958),
	.C2V_15 (C2V_190_994),
	.C2V_16 (C2V_190_1024),
	.C2V_17 (C2V_190_1099),
	.C2V_18 (C2V_190_1115),
	.C2V_19 (C2V_190_1341),
	.C2V_20 (C2V_190_1342),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU191 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_30_191),
	.V2C_2 (V2C_88_191),
	.V2C_3 (V2C_123_191),
	.V2C_4 (V2C_146_191),
	.V2C_5 (V2C_210_191),
	.V2C_6 (V2C_276_191),
	.V2C_7 (V2C_325_191),
	.V2C_8 (V2C_344_191),
	.V2C_9 (V2C_471_191),
	.V2C_10 (V2C_705_191),
	.V2C_11 (V2C_721_191),
	.V2C_12 (V2C_775_191),
	.V2C_13 (V2C_901_191),
	.V2C_14 (V2C_949_191),
	.V2C_15 (V2C_992_191),
	.V2C_16 (V2C_1044_191),
	.V2C_17 (V2C_1093_191),
	.V2C_18 (V2C_1141_191),
	.V2C_19 (V2C_1342_191),
	.V2C_20 (V2C_1343_191),
	.C2V_1 (C2V_191_30),
	.C2V_2 (C2V_191_88),
	.C2V_3 (C2V_191_123),
	.C2V_4 (C2V_191_146),
	.C2V_5 (C2V_191_210),
	.C2V_6 (C2V_191_276),
	.C2V_7 (C2V_191_325),
	.C2V_8 (C2V_191_344),
	.C2V_9 (C2V_191_471),
	.C2V_10 (C2V_191_705),
	.C2V_11 (C2V_191_721),
	.C2V_12 (C2V_191_775),
	.C2V_13 (C2V_191_901),
	.C2V_14 (C2V_191_949),
	.C2V_15 (C2V_191_992),
	.C2V_16 (C2V_191_1044),
	.C2V_17 (C2V_191_1093),
	.C2V_18 (C2V_191_1141),
	.C2V_19 (C2V_191_1342),
	.C2V_20 (C2V_191_1343),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU192 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_13_192),
	.V2C_2 (V2C_85_192),
	.V2C_3 (V2C_125_192),
	.V2C_4 (V2C_145_192),
	.V2C_5 (V2C_227_192),
	.V2C_6 (V2C_258_192),
	.V2C_7 (V2C_311_192),
	.V2C_8 (V2C_463_192),
	.V2C_9 (V2C_560_192),
	.V2C_10 (V2C_593_192),
	.V2C_11 (V2C_797_192),
	.V2C_12 (V2C_825_192),
	.V2C_13 (V2C_906_192),
	.V2C_14 (V2C_920_192),
	.V2C_15 (V2C_1003_192),
	.V2C_16 (V2C_1022_192),
	.V2C_17 (V2C_1086_192),
	.V2C_18 (V2C_1136_192),
	.V2C_19 (V2C_1343_192),
	.V2C_20 (V2C_1344_192),
	.C2V_1 (C2V_192_13),
	.C2V_2 (C2V_192_85),
	.C2V_3 (C2V_192_125),
	.C2V_4 (C2V_192_145),
	.C2V_5 (C2V_192_227),
	.C2V_6 (C2V_192_258),
	.C2V_7 (C2V_192_311),
	.C2V_8 (C2V_192_463),
	.C2V_9 (C2V_192_560),
	.C2V_10 (C2V_192_593),
	.C2V_11 (C2V_192_797),
	.C2V_12 (C2V_192_825),
	.C2V_13 (C2V_192_906),
	.C2V_14 (C2V_192_920),
	.C2V_15 (C2V_192_1003),
	.C2V_16 (C2V_192_1022),
	.C2V_17 (C2V_192_1086),
	.C2V_18 (C2V_192_1136),
	.C2V_19 (C2V_192_1343),
	.C2V_20 (C2V_192_1344),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU193 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_37_193),
	.V2C_2 (V2C_73_193),
	.V2C_3 (V2C_141_193),
	.V2C_4 (V2C_154_193),
	.V2C_5 (V2C_216_193),
	.V2C_6 (V2C_259_193),
	.V2C_7 (V2C_359_193),
	.V2C_8 (V2C_413_193),
	.V2C_9 (V2C_510_193),
	.V2C_10 (V2C_746_193),
	.V2C_11 (V2C_794_193),
	.V2C_12 (V2C_842_193),
	.V2C_13 (V2C_883_193),
	.V2C_14 (V2C_924_193),
	.V2C_15 (V2C_1006_193),
	.V2C_16 (V2C_1045_193),
	.V2C_17 (V2C_1071_193),
	.V2C_18 (V2C_1130_193),
	.V2C_19 (V2C_1344_193),
	.V2C_20 (V2C_1345_193),
	.C2V_1 (C2V_193_37),
	.C2V_2 (C2V_193_73),
	.C2V_3 (C2V_193_141),
	.C2V_4 (C2V_193_154),
	.C2V_5 (C2V_193_216),
	.C2V_6 (C2V_193_259),
	.C2V_7 (C2V_193_359),
	.C2V_8 (C2V_193_413),
	.C2V_9 (C2V_193_510),
	.C2V_10 (C2V_193_746),
	.C2V_11 (C2V_193_794),
	.C2V_12 (C2V_193_842),
	.C2V_13 (C2V_193_883),
	.C2V_14 (C2V_193_924),
	.C2V_15 (C2V_193_1006),
	.C2V_16 (C2V_193_1045),
	.C2V_17 (C2V_193_1071),
	.C2V_18 (C2V_193_1130),
	.C2V_19 (C2V_193_1344),
	.C2V_20 (C2V_193_1345),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU194 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_46_194),
	.V2C_2 (V2C_95_194),
	.V2C_3 (V2C_103_194),
	.V2C_4 (V2C_151_194),
	.V2C_5 (V2C_228_194),
	.V2C_6 (V2C_249_194),
	.V2C_7 (V2C_300_194),
	.V2C_8 (V2C_407_194),
	.V2C_9 (V2C_496_194),
	.V2C_10 (V2C_656_194),
	.V2C_11 (V2C_717_194),
	.V2C_12 (V2C_837_194),
	.V2C_13 (V2C_879_194),
	.V2C_14 (V2C_942_194),
	.V2C_15 (V2C_973_194),
	.V2C_16 (V2C_1053_194),
	.V2C_17 (V2C_1072_194),
	.V2C_18 (V2C_1151_194),
	.V2C_19 (V2C_1345_194),
	.V2C_20 (V2C_1346_194),
	.C2V_1 (C2V_194_46),
	.C2V_2 (C2V_194_95),
	.C2V_3 (C2V_194_103),
	.C2V_4 (C2V_194_151),
	.C2V_5 (C2V_194_228),
	.C2V_6 (C2V_194_249),
	.C2V_7 (C2V_194_300),
	.C2V_8 (C2V_194_407),
	.C2V_9 (C2V_194_496),
	.C2V_10 (C2V_194_656),
	.C2V_11 (C2V_194_717),
	.C2V_12 (C2V_194_837),
	.C2V_13 (C2V_194_879),
	.C2V_14 (C2V_194_942),
	.C2V_15 (C2V_194_973),
	.C2V_16 (C2V_194_1053),
	.C2V_17 (C2V_194_1072),
	.C2V_18 (C2V_194_1151),
	.C2V_19 (C2V_194_1345),
	.C2V_20 (C2V_194_1346),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU195 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_41_195),
	.V2C_2 (V2C_68_195),
	.V2C_3 (V2C_133_195),
	.V2C_4 (V2C_167_195),
	.V2C_5 (V2C_233_195),
	.V2C_6 (V2C_252_195),
	.V2C_7 (V2C_349_195),
	.V2C_8 (V2C_404_195),
	.V2C_9 (V2C_563_195),
	.V2C_10 (V2C_620_195),
	.V2C_11 (V2C_648_195),
	.V2C_12 (V2C_752_195),
	.V2C_13 (V2C_883_195),
	.V2C_14 (V2C_927_195),
	.V2C_15 (V2C_1000_195),
	.V2C_16 (V2C_1012_195),
	.V2C_17 (V2C_1090_195),
	.V2C_18 (V2C_1135_195),
	.V2C_19 (V2C_1346_195),
	.V2C_20 (V2C_1347_195),
	.C2V_1 (C2V_195_41),
	.C2V_2 (C2V_195_68),
	.C2V_3 (C2V_195_133),
	.C2V_4 (C2V_195_167),
	.C2V_5 (C2V_195_233),
	.C2V_6 (C2V_195_252),
	.C2V_7 (C2V_195_349),
	.C2V_8 (C2V_195_404),
	.C2V_9 (C2V_195_563),
	.C2V_10 (C2V_195_620),
	.C2V_11 (C2V_195_648),
	.C2V_12 (C2V_195_752),
	.C2V_13 (C2V_195_883),
	.C2V_14 (C2V_195_927),
	.C2V_15 (C2V_195_1000),
	.C2V_16 (C2V_195_1012),
	.C2V_17 (C2V_195_1090),
	.C2V_18 (C2V_195_1135),
	.C2V_19 (C2V_195_1346),
	.C2V_20 (C2V_195_1347),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU196 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_12_196),
	.V2C_2 (V2C_71_196),
	.V2C_3 (V2C_110_196),
	.V2C_4 (V2C_166_196),
	.V2C_5 (V2C_231_196),
	.V2C_6 (V2C_285_196),
	.V2C_7 (V2C_461_196),
	.V2C_8 (V2C_501_196),
	.V2C_9 (V2C_537_196),
	.V2C_10 (V2C_599_196),
	.V2C_11 (V2C_672_196),
	.V2C_12 (V2C_718_196),
	.V2C_13 (V2C_887_196),
	.V2C_14 (V2C_959_196),
	.V2C_15 (V2C_995_196),
	.V2C_16 (V2C_1025_196),
	.V2C_17 (V2C_1100_196),
	.V2C_18 (V2C_1116_196),
	.V2C_19 (V2C_1347_196),
	.V2C_20 (V2C_1348_196),
	.C2V_1 (C2V_196_12),
	.C2V_2 (C2V_196_71),
	.C2V_3 (C2V_196_110),
	.C2V_4 (C2V_196_166),
	.C2V_5 (C2V_196_231),
	.C2V_6 (C2V_196_285),
	.C2V_7 (C2V_196_461),
	.C2V_8 (C2V_196_501),
	.C2V_9 (C2V_196_537),
	.C2V_10 (C2V_196_599),
	.C2V_11 (C2V_196_672),
	.C2V_12 (C2V_196_718),
	.C2V_13 (C2V_196_887),
	.C2V_14 (C2V_196_959),
	.C2V_15 (C2V_196_995),
	.C2V_16 (C2V_196_1025),
	.C2V_17 (C2V_196_1100),
	.C2V_18 (C2V_196_1116),
	.C2V_19 (C2V_196_1347),
	.C2V_20 (C2V_196_1348),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU197 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_31_197),
	.V2C_2 (V2C_89_197),
	.V2C_3 (V2C_124_197),
	.V2C_4 (V2C_147_197),
	.V2C_5 (V2C_211_197),
	.V2C_6 (V2C_277_197),
	.V2C_7 (V2C_326_197),
	.V2C_8 (V2C_345_197),
	.V2C_9 (V2C_472_197),
	.V2C_10 (V2C_706_197),
	.V2C_11 (V2C_722_197),
	.V2C_12 (V2C_776_197),
	.V2C_13 (V2C_902_197),
	.V2C_14 (V2C_950_197),
	.V2C_15 (V2C_993_197),
	.V2C_16 (V2C_1045_197),
	.V2C_17 (V2C_1094_197),
	.V2C_18 (V2C_1142_197),
	.V2C_19 (V2C_1348_197),
	.V2C_20 (V2C_1349_197),
	.C2V_1 (C2V_197_31),
	.C2V_2 (C2V_197_89),
	.C2V_3 (C2V_197_124),
	.C2V_4 (C2V_197_147),
	.C2V_5 (C2V_197_211),
	.C2V_6 (C2V_197_277),
	.C2V_7 (C2V_197_326),
	.C2V_8 (C2V_197_345),
	.C2V_9 (C2V_197_472),
	.C2V_10 (C2V_197_706),
	.C2V_11 (C2V_197_722),
	.C2V_12 (C2V_197_776),
	.C2V_13 (C2V_197_902),
	.C2V_14 (C2V_197_950),
	.C2V_15 (C2V_197_993),
	.C2V_16 (C2V_197_1045),
	.C2V_17 (C2V_197_1094),
	.C2V_18 (C2V_197_1142),
	.C2V_19 (C2V_197_1348),
	.C2V_20 (C2V_197_1349),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU198 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_14_198),
	.V2C_2 (V2C_86_198),
	.V2C_3 (V2C_126_198),
	.V2C_4 (V2C_146_198),
	.V2C_5 (V2C_228_198),
	.V2C_6 (V2C_259_198),
	.V2C_7 (V2C_312_198),
	.V2C_8 (V2C_464_198),
	.V2C_9 (V2C_561_198),
	.V2C_10 (V2C_594_198),
	.V2C_11 (V2C_798_198),
	.V2C_12 (V2C_826_198),
	.V2C_13 (V2C_907_198),
	.V2C_14 (V2C_921_198),
	.V2C_15 (V2C_1004_198),
	.V2C_16 (V2C_1023_198),
	.V2C_17 (V2C_1087_198),
	.V2C_18 (V2C_1137_198),
	.V2C_19 (V2C_1349_198),
	.V2C_20 (V2C_1350_198),
	.C2V_1 (C2V_198_14),
	.C2V_2 (C2V_198_86),
	.C2V_3 (C2V_198_126),
	.C2V_4 (C2V_198_146),
	.C2V_5 (C2V_198_228),
	.C2V_6 (C2V_198_259),
	.C2V_7 (C2V_198_312),
	.C2V_8 (C2V_198_464),
	.C2V_9 (C2V_198_561),
	.C2V_10 (C2V_198_594),
	.C2V_11 (C2V_198_798),
	.C2V_12 (C2V_198_826),
	.C2V_13 (C2V_198_907),
	.C2V_14 (C2V_198_921),
	.C2V_15 (C2V_198_1004),
	.C2V_16 (C2V_198_1023),
	.C2V_17 (C2V_198_1087),
	.C2V_18 (C2V_198_1137),
	.C2V_19 (C2V_198_1349),
	.C2V_20 (C2V_198_1350),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU199 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_38_199),
	.V2C_2 (V2C_74_199),
	.V2C_3 (V2C_142_199),
	.V2C_4 (V2C_155_199),
	.V2C_5 (V2C_217_199),
	.V2C_6 (V2C_260_199),
	.V2C_7 (V2C_360_199),
	.V2C_8 (V2C_414_199),
	.V2C_9 (V2C_511_199),
	.V2C_10 (V2C_747_199),
	.V2C_11 (V2C_795_199),
	.V2C_12 (V2C_843_199),
	.V2C_13 (V2C_884_199),
	.V2C_14 (V2C_925_199),
	.V2C_15 (V2C_1007_199),
	.V2C_16 (V2C_1046_199),
	.V2C_17 (V2C_1072_199),
	.V2C_18 (V2C_1131_199),
	.V2C_19 (V2C_1350_199),
	.V2C_20 (V2C_1351_199),
	.C2V_1 (C2V_199_38),
	.C2V_2 (C2V_199_74),
	.C2V_3 (C2V_199_142),
	.C2V_4 (C2V_199_155),
	.C2V_5 (C2V_199_217),
	.C2V_6 (C2V_199_260),
	.C2V_7 (C2V_199_360),
	.C2V_8 (C2V_199_414),
	.C2V_9 (C2V_199_511),
	.C2V_10 (C2V_199_747),
	.C2V_11 (C2V_199_795),
	.C2V_12 (C2V_199_843),
	.C2V_13 (C2V_199_884),
	.C2V_14 (C2V_199_925),
	.C2V_15 (C2V_199_1007),
	.C2V_16 (C2V_199_1046),
	.C2V_17 (C2V_199_1072),
	.C2V_18 (C2V_199_1131),
	.C2V_19 (C2V_199_1350),
	.C2V_20 (C2V_199_1351),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU200 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_47_200),
	.V2C_2 (V2C_96_200),
	.V2C_3 (V2C_104_200),
	.V2C_4 (V2C_152_200),
	.V2C_5 (V2C_229_200),
	.V2C_6 (V2C_250_200),
	.V2C_7 (V2C_301_200),
	.V2C_8 (V2C_408_200),
	.V2C_9 (V2C_497_200),
	.V2C_10 (V2C_657_200),
	.V2C_11 (V2C_718_200),
	.V2C_12 (V2C_838_200),
	.V2C_13 (V2C_880_200),
	.V2C_14 (V2C_943_200),
	.V2C_15 (V2C_974_200),
	.V2C_16 (V2C_1054_200),
	.V2C_17 (V2C_1073_200),
	.V2C_18 (V2C_1152_200),
	.V2C_19 (V2C_1351_200),
	.V2C_20 (V2C_1352_200),
	.C2V_1 (C2V_200_47),
	.C2V_2 (C2V_200_96),
	.C2V_3 (C2V_200_104),
	.C2V_4 (C2V_200_152),
	.C2V_5 (C2V_200_229),
	.C2V_6 (C2V_200_250),
	.C2V_7 (C2V_200_301),
	.C2V_8 (C2V_200_408),
	.C2V_9 (C2V_200_497),
	.C2V_10 (C2V_200_657),
	.C2V_11 (C2V_200_718),
	.C2V_12 (C2V_200_838),
	.C2V_13 (C2V_200_880),
	.C2V_14 (C2V_200_943),
	.C2V_15 (C2V_200_974),
	.C2V_16 (C2V_200_1054),
	.C2V_17 (C2V_200_1073),
	.C2V_18 (C2V_200_1152),
	.C2V_19 (C2V_200_1351),
	.C2V_20 (C2V_200_1352),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU201 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_42_201),
	.V2C_2 (V2C_69_201),
	.V2C_3 (V2C_134_201),
	.V2C_4 (V2C_168_201),
	.V2C_5 (V2C_234_201),
	.V2C_6 (V2C_253_201),
	.V2C_7 (V2C_350_201),
	.V2C_8 (V2C_405_201),
	.V2C_9 (V2C_564_201),
	.V2C_10 (V2C_621_201),
	.V2C_11 (V2C_649_201),
	.V2C_12 (V2C_753_201),
	.V2C_13 (V2C_884_201),
	.V2C_14 (V2C_928_201),
	.V2C_15 (V2C_1001_201),
	.V2C_16 (V2C_1013_201),
	.V2C_17 (V2C_1091_201),
	.V2C_18 (V2C_1136_201),
	.V2C_19 (V2C_1352_201),
	.V2C_20 (V2C_1353_201),
	.C2V_1 (C2V_201_42),
	.C2V_2 (C2V_201_69),
	.C2V_3 (C2V_201_134),
	.C2V_4 (C2V_201_168),
	.C2V_5 (C2V_201_234),
	.C2V_6 (C2V_201_253),
	.C2V_7 (C2V_201_350),
	.C2V_8 (C2V_201_405),
	.C2V_9 (C2V_201_564),
	.C2V_10 (C2V_201_621),
	.C2V_11 (C2V_201_649),
	.C2V_12 (C2V_201_753),
	.C2V_13 (C2V_201_884),
	.C2V_14 (C2V_201_928),
	.C2V_15 (C2V_201_1001),
	.C2V_16 (C2V_201_1013),
	.C2V_17 (C2V_201_1091),
	.C2V_18 (C2V_201_1136),
	.C2V_19 (C2V_201_1352),
	.C2V_20 (C2V_201_1353),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU202 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_13_202),
	.V2C_2 (V2C_72_202),
	.V2C_3 (V2C_111_202),
	.V2C_4 (V2C_167_202),
	.V2C_5 (V2C_232_202),
	.V2C_6 (V2C_286_202),
	.V2C_7 (V2C_462_202),
	.V2C_8 (V2C_502_202),
	.V2C_9 (V2C_538_202),
	.V2C_10 (V2C_600_202),
	.V2C_11 (V2C_625_202),
	.V2C_12 (V2C_719_202),
	.V2C_13 (V2C_888_202),
	.V2C_14 (V2C_960_202),
	.V2C_15 (V2C_996_202),
	.V2C_16 (V2C_1026_202),
	.V2C_17 (V2C_1101_202),
	.V2C_18 (V2C_1117_202),
	.V2C_19 (V2C_1353_202),
	.V2C_20 (V2C_1354_202),
	.C2V_1 (C2V_202_13),
	.C2V_2 (C2V_202_72),
	.C2V_3 (C2V_202_111),
	.C2V_4 (C2V_202_167),
	.C2V_5 (C2V_202_232),
	.C2V_6 (C2V_202_286),
	.C2V_7 (C2V_202_462),
	.C2V_8 (C2V_202_502),
	.C2V_9 (C2V_202_538),
	.C2V_10 (C2V_202_600),
	.C2V_11 (C2V_202_625),
	.C2V_12 (C2V_202_719),
	.C2V_13 (C2V_202_888),
	.C2V_14 (C2V_202_960),
	.C2V_15 (C2V_202_996),
	.C2V_16 (C2V_202_1026),
	.C2V_17 (C2V_202_1101),
	.C2V_18 (C2V_202_1117),
	.C2V_19 (C2V_202_1353),
	.C2V_20 (C2V_202_1354),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU203 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_32_203),
	.V2C_2 (V2C_90_203),
	.V2C_3 (V2C_125_203),
	.V2C_4 (V2C_148_203),
	.V2C_5 (V2C_212_203),
	.V2C_6 (V2C_278_203),
	.V2C_7 (V2C_327_203),
	.V2C_8 (V2C_346_203),
	.V2C_9 (V2C_473_203),
	.V2C_10 (V2C_707_203),
	.V2C_11 (V2C_723_203),
	.V2C_12 (V2C_777_203),
	.V2C_13 (V2C_903_203),
	.V2C_14 (V2C_951_203),
	.V2C_15 (V2C_994_203),
	.V2C_16 (V2C_1046_203),
	.V2C_17 (V2C_1095_203),
	.V2C_18 (V2C_1143_203),
	.V2C_19 (V2C_1354_203),
	.V2C_20 (V2C_1355_203),
	.C2V_1 (C2V_203_32),
	.C2V_2 (C2V_203_90),
	.C2V_3 (C2V_203_125),
	.C2V_4 (C2V_203_148),
	.C2V_5 (C2V_203_212),
	.C2V_6 (C2V_203_278),
	.C2V_7 (C2V_203_327),
	.C2V_8 (C2V_203_346),
	.C2V_9 (C2V_203_473),
	.C2V_10 (C2V_203_707),
	.C2V_11 (C2V_203_723),
	.C2V_12 (C2V_203_777),
	.C2V_13 (C2V_203_903),
	.C2V_14 (C2V_203_951),
	.C2V_15 (C2V_203_994),
	.C2V_16 (C2V_203_1046),
	.C2V_17 (C2V_203_1095),
	.C2V_18 (C2V_203_1143),
	.C2V_19 (C2V_203_1354),
	.C2V_20 (C2V_203_1355),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU204 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_15_204),
	.V2C_2 (V2C_87_204),
	.V2C_3 (V2C_127_204),
	.V2C_4 (V2C_147_204),
	.V2C_5 (V2C_229_204),
	.V2C_6 (V2C_260_204),
	.V2C_7 (V2C_313_204),
	.V2C_8 (V2C_465_204),
	.V2C_9 (V2C_562_204),
	.V2C_10 (V2C_595_204),
	.V2C_11 (V2C_799_204),
	.V2C_12 (V2C_827_204),
	.V2C_13 (V2C_908_204),
	.V2C_14 (V2C_922_204),
	.V2C_15 (V2C_1005_204),
	.V2C_16 (V2C_1024_204),
	.V2C_17 (V2C_1088_204),
	.V2C_18 (V2C_1138_204),
	.V2C_19 (V2C_1355_204),
	.V2C_20 (V2C_1356_204),
	.C2V_1 (C2V_204_15),
	.C2V_2 (C2V_204_87),
	.C2V_3 (C2V_204_127),
	.C2V_4 (C2V_204_147),
	.C2V_5 (C2V_204_229),
	.C2V_6 (C2V_204_260),
	.C2V_7 (C2V_204_313),
	.C2V_8 (C2V_204_465),
	.C2V_9 (C2V_204_562),
	.C2V_10 (C2V_204_595),
	.C2V_11 (C2V_204_799),
	.C2V_12 (C2V_204_827),
	.C2V_13 (C2V_204_908),
	.C2V_14 (C2V_204_922),
	.C2V_15 (C2V_204_1005),
	.C2V_16 (C2V_204_1024),
	.C2V_17 (C2V_204_1088),
	.C2V_18 (C2V_204_1138),
	.C2V_19 (C2V_204_1355),
	.C2V_20 (C2V_204_1356),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU205 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_39_205),
	.V2C_2 (V2C_75_205),
	.V2C_3 (V2C_143_205),
	.V2C_4 (V2C_156_205),
	.V2C_5 (V2C_218_205),
	.V2C_6 (V2C_261_205),
	.V2C_7 (V2C_361_205),
	.V2C_8 (V2C_415_205),
	.V2C_9 (V2C_512_205),
	.V2C_10 (V2C_748_205),
	.V2C_11 (V2C_796_205),
	.V2C_12 (V2C_844_205),
	.V2C_13 (V2C_885_205),
	.V2C_14 (V2C_926_205),
	.V2C_15 (V2C_1008_205),
	.V2C_16 (V2C_1047_205),
	.V2C_17 (V2C_1073_205),
	.V2C_18 (V2C_1132_205),
	.V2C_19 (V2C_1356_205),
	.V2C_20 (V2C_1357_205),
	.C2V_1 (C2V_205_39),
	.C2V_2 (C2V_205_75),
	.C2V_3 (C2V_205_143),
	.C2V_4 (C2V_205_156),
	.C2V_5 (C2V_205_218),
	.C2V_6 (C2V_205_261),
	.C2V_7 (C2V_205_361),
	.C2V_8 (C2V_205_415),
	.C2V_9 (C2V_205_512),
	.C2V_10 (C2V_205_748),
	.C2V_11 (C2V_205_796),
	.C2V_12 (C2V_205_844),
	.C2V_13 (C2V_205_885),
	.C2V_14 (C2V_205_926),
	.C2V_15 (C2V_205_1008),
	.C2V_16 (C2V_205_1047),
	.C2V_17 (C2V_205_1073),
	.C2V_18 (C2V_205_1132),
	.C2V_19 (C2V_205_1356),
	.C2V_20 (C2V_205_1357),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU206 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_48_206),
	.V2C_2 (V2C_49_206),
	.V2C_3 (V2C_105_206),
	.V2C_4 (V2C_153_206),
	.V2C_5 (V2C_230_206),
	.V2C_6 (V2C_251_206),
	.V2C_7 (V2C_302_206),
	.V2C_8 (V2C_409_206),
	.V2C_9 (V2C_498_206),
	.V2C_10 (V2C_658_206),
	.V2C_11 (V2C_719_206),
	.V2C_12 (V2C_839_206),
	.V2C_13 (V2C_881_206),
	.V2C_14 (V2C_944_206),
	.V2C_15 (V2C_975_206),
	.V2C_16 (V2C_1055_206),
	.V2C_17 (V2C_1074_206),
	.V2C_18 (V2C_1105_206),
	.V2C_19 (V2C_1357_206),
	.V2C_20 (V2C_1358_206),
	.C2V_1 (C2V_206_48),
	.C2V_2 (C2V_206_49),
	.C2V_3 (C2V_206_105),
	.C2V_4 (C2V_206_153),
	.C2V_5 (C2V_206_230),
	.C2V_6 (C2V_206_251),
	.C2V_7 (C2V_206_302),
	.C2V_8 (C2V_206_409),
	.C2V_9 (C2V_206_498),
	.C2V_10 (C2V_206_658),
	.C2V_11 (C2V_206_719),
	.C2V_12 (C2V_206_839),
	.C2V_13 (C2V_206_881),
	.C2V_14 (C2V_206_944),
	.C2V_15 (C2V_206_975),
	.C2V_16 (C2V_206_1055),
	.C2V_17 (C2V_206_1074),
	.C2V_18 (C2V_206_1105),
	.C2V_19 (C2V_206_1357),
	.C2V_20 (C2V_206_1358),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU207 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_43_207),
	.V2C_2 (V2C_70_207),
	.V2C_3 (V2C_135_207),
	.V2C_4 (V2C_169_207),
	.V2C_5 (V2C_235_207),
	.V2C_6 (V2C_254_207),
	.V2C_7 (V2C_351_207),
	.V2C_8 (V2C_406_207),
	.V2C_9 (V2C_565_207),
	.V2C_10 (V2C_622_207),
	.V2C_11 (V2C_650_207),
	.V2C_12 (V2C_754_207),
	.V2C_13 (V2C_885_207),
	.V2C_14 (V2C_929_207),
	.V2C_15 (V2C_1002_207),
	.V2C_16 (V2C_1014_207),
	.V2C_17 (V2C_1092_207),
	.V2C_18 (V2C_1137_207),
	.V2C_19 (V2C_1358_207),
	.V2C_20 (V2C_1359_207),
	.C2V_1 (C2V_207_43),
	.C2V_2 (C2V_207_70),
	.C2V_3 (C2V_207_135),
	.C2V_4 (C2V_207_169),
	.C2V_5 (C2V_207_235),
	.C2V_6 (C2V_207_254),
	.C2V_7 (C2V_207_351),
	.C2V_8 (C2V_207_406),
	.C2V_9 (C2V_207_565),
	.C2V_10 (C2V_207_622),
	.C2V_11 (C2V_207_650),
	.C2V_12 (C2V_207_754),
	.C2V_13 (C2V_207_885),
	.C2V_14 (C2V_207_929),
	.C2V_15 (C2V_207_1002),
	.C2V_16 (C2V_207_1014),
	.C2V_17 (C2V_207_1092),
	.C2V_18 (C2V_207_1137),
	.C2V_19 (C2V_207_1358),
	.C2V_20 (C2V_207_1359),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU208 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_14_208),
	.V2C_2 (V2C_73_208),
	.V2C_3 (V2C_112_208),
	.V2C_4 (V2C_168_208),
	.V2C_5 (V2C_233_208),
	.V2C_6 (V2C_287_208),
	.V2C_7 (V2C_463_208),
	.V2C_8 (V2C_503_208),
	.V2C_9 (V2C_539_208),
	.V2C_10 (V2C_601_208),
	.V2C_11 (V2C_626_208),
	.V2C_12 (V2C_720_208),
	.V2C_13 (V2C_889_208),
	.V2C_14 (V2C_913_208),
	.V2C_15 (V2C_997_208),
	.V2C_16 (V2C_1027_208),
	.V2C_17 (V2C_1102_208),
	.V2C_18 (V2C_1118_208),
	.V2C_19 (V2C_1359_208),
	.V2C_20 (V2C_1360_208),
	.C2V_1 (C2V_208_14),
	.C2V_2 (C2V_208_73),
	.C2V_3 (C2V_208_112),
	.C2V_4 (C2V_208_168),
	.C2V_5 (C2V_208_233),
	.C2V_6 (C2V_208_287),
	.C2V_7 (C2V_208_463),
	.C2V_8 (C2V_208_503),
	.C2V_9 (C2V_208_539),
	.C2V_10 (C2V_208_601),
	.C2V_11 (C2V_208_626),
	.C2V_12 (C2V_208_720),
	.C2V_13 (C2V_208_889),
	.C2V_14 (C2V_208_913),
	.C2V_15 (C2V_208_997),
	.C2V_16 (C2V_208_1027),
	.C2V_17 (C2V_208_1102),
	.C2V_18 (C2V_208_1118),
	.C2V_19 (C2V_208_1359),
	.C2V_20 (C2V_208_1360),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU209 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_33_209),
	.V2C_2 (V2C_91_209),
	.V2C_3 (V2C_126_209),
	.V2C_4 (V2C_149_209),
	.V2C_5 (V2C_213_209),
	.V2C_6 (V2C_279_209),
	.V2C_7 (V2C_328_209),
	.V2C_8 (V2C_347_209),
	.V2C_9 (V2C_474_209),
	.V2C_10 (V2C_708_209),
	.V2C_11 (V2C_724_209),
	.V2C_12 (V2C_778_209),
	.V2C_13 (V2C_904_209),
	.V2C_14 (V2C_952_209),
	.V2C_15 (V2C_995_209),
	.V2C_16 (V2C_1047_209),
	.V2C_17 (V2C_1096_209),
	.V2C_18 (V2C_1144_209),
	.V2C_19 (V2C_1360_209),
	.V2C_20 (V2C_1361_209),
	.C2V_1 (C2V_209_33),
	.C2V_2 (C2V_209_91),
	.C2V_3 (C2V_209_126),
	.C2V_4 (C2V_209_149),
	.C2V_5 (C2V_209_213),
	.C2V_6 (C2V_209_279),
	.C2V_7 (C2V_209_328),
	.C2V_8 (C2V_209_347),
	.C2V_9 (C2V_209_474),
	.C2V_10 (C2V_209_708),
	.C2V_11 (C2V_209_724),
	.C2V_12 (C2V_209_778),
	.C2V_13 (C2V_209_904),
	.C2V_14 (C2V_209_952),
	.C2V_15 (C2V_209_995),
	.C2V_16 (C2V_209_1047),
	.C2V_17 (C2V_209_1096),
	.C2V_18 (C2V_209_1144),
	.C2V_19 (C2V_209_1360),
	.C2V_20 (C2V_209_1361),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU210 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_16_210),
	.V2C_2 (V2C_88_210),
	.V2C_3 (V2C_128_210),
	.V2C_4 (V2C_148_210),
	.V2C_5 (V2C_230_210),
	.V2C_6 (V2C_261_210),
	.V2C_7 (V2C_314_210),
	.V2C_8 (V2C_466_210),
	.V2C_9 (V2C_563_210),
	.V2C_10 (V2C_596_210),
	.V2C_11 (V2C_800_210),
	.V2C_12 (V2C_828_210),
	.V2C_13 (V2C_909_210),
	.V2C_14 (V2C_923_210),
	.V2C_15 (V2C_1006_210),
	.V2C_16 (V2C_1025_210),
	.V2C_17 (V2C_1089_210),
	.V2C_18 (V2C_1139_210),
	.V2C_19 (V2C_1361_210),
	.V2C_20 (V2C_1362_210),
	.C2V_1 (C2V_210_16),
	.C2V_2 (C2V_210_88),
	.C2V_3 (C2V_210_128),
	.C2V_4 (C2V_210_148),
	.C2V_5 (C2V_210_230),
	.C2V_6 (C2V_210_261),
	.C2V_7 (C2V_210_314),
	.C2V_8 (C2V_210_466),
	.C2V_9 (C2V_210_563),
	.C2V_10 (C2V_210_596),
	.C2V_11 (C2V_210_800),
	.C2V_12 (C2V_210_828),
	.C2V_13 (C2V_210_909),
	.C2V_14 (C2V_210_923),
	.C2V_15 (C2V_210_1006),
	.C2V_16 (C2V_210_1025),
	.C2V_17 (C2V_210_1089),
	.C2V_18 (C2V_210_1139),
	.C2V_19 (C2V_210_1361),
	.C2V_20 (C2V_210_1362),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU211 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_40_211),
	.V2C_2 (V2C_76_211),
	.V2C_3 (V2C_144_211),
	.V2C_4 (V2C_157_211),
	.V2C_5 (V2C_219_211),
	.V2C_6 (V2C_262_211),
	.V2C_7 (V2C_362_211),
	.V2C_8 (V2C_416_211),
	.V2C_9 (V2C_513_211),
	.V2C_10 (V2C_749_211),
	.V2C_11 (V2C_797_211),
	.V2C_12 (V2C_845_211),
	.V2C_13 (V2C_886_211),
	.V2C_14 (V2C_927_211),
	.V2C_15 (V2C_961_211),
	.V2C_16 (V2C_1048_211),
	.V2C_17 (V2C_1074_211),
	.V2C_18 (V2C_1133_211),
	.V2C_19 (V2C_1362_211),
	.V2C_20 (V2C_1363_211),
	.C2V_1 (C2V_211_40),
	.C2V_2 (C2V_211_76),
	.C2V_3 (C2V_211_144),
	.C2V_4 (C2V_211_157),
	.C2V_5 (C2V_211_219),
	.C2V_6 (C2V_211_262),
	.C2V_7 (C2V_211_362),
	.C2V_8 (C2V_211_416),
	.C2V_9 (C2V_211_513),
	.C2V_10 (C2V_211_749),
	.C2V_11 (C2V_211_797),
	.C2V_12 (C2V_211_845),
	.C2V_13 (C2V_211_886),
	.C2V_14 (C2V_211_927),
	.C2V_15 (C2V_211_961),
	.C2V_16 (C2V_211_1048),
	.C2V_17 (C2V_211_1074),
	.C2V_18 (C2V_211_1133),
	.C2V_19 (C2V_211_1362),
	.C2V_20 (C2V_211_1363),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU212 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_1_212),
	.V2C_2 (V2C_50_212),
	.V2C_3 (V2C_106_212),
	.V2C_4 (V2C_154_212),
	.V2C_5 (V2C_231_212),
	.V2C_6 (V2C_252_212),
	.V2C_7 (V2C_303_212),
	.V2C_8 (V2C_410_212),
	.V2C_9 (V2C_499_212),
	.V2C_10 (V2C_659_212),
	.V2C_11 (V2C_720_212),
	.V2C_12 (V2C_840_212),
	.V2C_13 (V2C_882_212),
	.V2C_14 (V2C_945_212),
	.V2C_15 (V2C_976_212),
	.V2C_16 (V2C_1056_212),
	.V2C_17 (V2C_1075_212),
	.V2C_18 (V2C_1106_212),
	.V2C_19 (V2C_1363_212),
	.V2C_20 (V2C_1364_212),
	.C2V_1 (C2V_212_1),
	.C2V_2 (C2V_212_50),
	.C2V_3 (C2V_212_106),
	.C2V_4 (C2V_212_154),
	.C2V_5 (C2V_212_231),
	.C2V_6 (C2V_212_252),
	.C2V_7 (C2V_212_303),
	.C2V_8 (C2V_212_410),
	.C2V_9 (C2V_212_499),
	.C2V_10 (C2V_212_659),
	.C2V_11 (C2V_212_720),
	.C2V_12 (C2V_212_840),
	.C2V_13 (C2V_212_882),
	.C2V_14 (C2V_212_945),
	.C2V_15 (C2V_212_976),
	.C2V_16 (C2V_212_1056),
	.C2V_17 (C2V_212_1075),
	.C2V_18 (C2V_212_1106),
	.C2V_19 (C2V_212_1363),
	.C2V_20 (C2V_212_1364),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU213 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_44_213),
	.V2C_2 (V2C_71_213),
	.V2C_3 (V2C_136_213),
	.V2C_4 (V2C_170_213),
	.V2C_5 (V2C_236_213),
	.V2C_6 (V2C_255_213),
	.V2C_7 (V2C_352_213),
	.V2C_8 (V2C_407_213),
	.V2C_9 (V2C_566_213),
	.V2C_10 (V2C_623_213),
	.V2C_11 (V2C_651_213),
	.V2C_12 (V2C_755_213),
	.V2C_13 (V2C_886_213),
	.V2C_14 (V2C_930_213),
	.V2C_15 (V2C_1003_213),
	.V2C_16 (V2C_1015_213),
	.V2C_17 (V2C_1093_213),
	.V2C_18 (V2C_1138_213),
	.V2C_19 (V2C_1364_213),
	.V2C_20 (V2C_1365_213),
	.C2V_1 (C2V_213_44),
	.C2V_2 (C2V_213_71),
	.C2V_3 (C2V_213_136),
	.C2V_4 (C2V_213_170),
	.C2V_5 (C2V_213_236),
	.C2V_6 (C2V_213_255),
	.C2V_7 (C2V_213_352),
	.C2V_8 (C2V_213_407),
	.C2V_9 (C2V_213_566),
	.C2V_10 (C2V_213_623),
	.C2V_11 (C2V_213_651),
	.C2V_12 (C2V_213_755),
	.C2V_13 (C2V_213_886),
	.C2V_14 (C2V_213_930),
	.C2V_15 (C2V_213_1003),
	.C2V_16 (C2V_213_1015),
	.C2V_17 (C2V_213_1093),
	.C2V_18 (C2V_213_1138),
	.C2V_19 (C2V_213_1364),
	.C2V_20 (C2V_213_1365),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU214 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_15_214),
	.V2C_2 (V2C_74_214),
	.V2C_3 (V2C_113_214),
	.V2C_4 (V2C_169_214),
	.V2C_5 (V2C_234_214),
	.V2C_6 (V2C_288_214),
	.V2C_7 (V2C_464_214),
	.V2C_8 (V2C_504_214),
	.V2C_9 (V2C_540_214),
	.V2C_10 (V2C_602_214),
	.V2C_11 (V2C_627_214),
	.V2C_12 (V2C_673_214),
	.V2C_13 (V2C_890_214),
	.V2C_14 (V2C_914_214),
	.V2C_15 (V2C_998_214),
	.V2C_16 (V2C_1028_214),
	.V2C_17 (V2C_1103_214),
	.V2C_18 (V2C_1119_214),
	.V2C_19 (V2C_1365_214),
	.V2C_20 (V2C_1366_214),
	.C2V_1 (C2V_214_15),
	.C2V_2 (C2V_214_74),
	.C2V_3 (C2V_214_113),
	.C2V_4 (C2V_214_169),
	.C2V_5 (C2V_214_234),
	.C2V_6 (C2V_214_288),
	.C2V_7 (C2V_214_464),
	.C2V_8 (C2V_214_504),
	.C2V_9 (C2V_214_540),
	.C2V_10 (C2V_214_602),
	.C2V_11 (C2V_214_627),
	.C2V_12 (C2V_214_673),
	.C2V_13 (C2V_214_890),
	.C2V_14 (C2V_214_914),
	.C2V_15 (C2V_214_998),
	.C2V_16 (C2V_214_1028),
	.C2V_17 (C2V_214_1103),
	.C2V_18 (C2V_214_1119),
	.C2V_19 (C2V_214_1365),
	.C2V_20 (C2V_214_1366),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU215 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_34_215),
	.V2C_2 (V2C_92_215),
	.V2C_3 (V2C_127_215),
	.V2C_4 (V2C_150_215),
	.V2C_5 (V2C_214_215),
	.V2C_6 (V2C_280_215),
	.V2C_7 (V2C_329_215),
	.V2C_8 (V2C_348_215),
	.V2C_9 (V2C_475_215),
	.V2C_10 (V2C_709_215),
	.V2C_11 (V2C_725_215),
	.V2C_12 (V2C_779_215),
	.V2C_13 (V2C_905_215),
	.V2C_14 (V2C_953_215),
	.V2C_15 (V2C_996_215),
	.V2C_16 (V2C_1048_215),
	.V2C_17 (V2C_1097_215),
	.V2C_18 (V2C_1145_215),
	.V2C_19 (V2C_1366_215),
	.V2C_20 (V2C_1367_215),
	.C2V_1 (C2V_215_34),
	.C2V_2 (C2V_215_92),
	.C2V_3 (C2V_215_127),
	.C2V_4 (C2V_215_150),
	.C2V_5 (C2V_215_214),
	.C2V_6 (C2V_215_280),
	.C2V_7 (C2V_215_329),
	.C2V_8 (C2V_215_348),
	.C2V_9 (C2V_215_475),
	.C2V_10 (C2V_215_709),
	.C2V_11 (C2V_215_725),
	.C2V_12 (C2V_215_779),
	.C2V_13 (C2V_215_905),
	.C2V_14 (C2V_215_953),
	.C2V_15 (C2V_215_996),
	.C2V_16 (C2V_215_1048),
	.C2V_17 (C2V_215_1097),
	.C2V_18 (C2V_215_1145),
	.C2V_19 (C2V_215_1366),
	.C2V_20 (C2V_215_1367),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU216 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_17_216),
	.V2C_2 (V2C_89_216),
	.V2C_3 (V2C_129_216),
	.V2C_4 (V2C_149_216),
	.V2C_5 (V2C_231_216),
	.V2C_6 (V2C_262_216),
	.V2C_7 (V2C_315_216),
	.V2C_8 (V2C_467_216),
	.V2C_9 (V2C_564_216),
	.V2C_10 (V2C_597_216),
	.V2C_11 (V2C_801_216),
	.V2C_12 (V2C_829_216),
	.V2C_13 (V2C_910_216),
	.V2C_14 (V2C_924_216),
	.V2C_15 (V2C_1007_216),
	.V2C_16 (V2C_1026_216),
	.V2C_17 (V2C_1090_216),
	.V2C_18 (V2C_1140_216),
	.V2C_19 (V2C_1367_216),
	.V2C_20 (V2C_1368_216),
	.C2V_1 (C2V_216_17),
	.C2V_2 (C2V_216_89),
	.C2V_3 (C2V_216_129),
	.C2V_4 (C2V_216_149),
	.C2V_5 (C2V_216_231),
	.C2V_6 (C2V_216_262),
	.C2V_7 (C2V_216_315),
	.C2V_8 (C2V_216_467),
	.C2V_9 (C2V_216_564),
	.C2V_10 (C2V_216_597),
	.C2V_11 (C2V_216_801),
	.C2V_12 (C2V_216_829),
	.C2V_13 (C2V_216_910),
	.C2V_14 (C2V_216_924),
	.C2V_15 (C2V_216_1007),
	.C2V_16 (C2V_216_1026),
	.C2V_17 (C2V_216_1090),
	.C2V_18 (C2V_216_1140),
	.C2V_19 (C2V_216_1367),
	.C2V_20 (C2V_216_1368),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU217 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_41_217),
	.V2C_2 (V2C_77_217),
	.V2C_3 (V2C_97_217),
	.V2C_4 (V2C_158_217),
	.V2C_5 (V2C_220_217),
	.V2C_6 (V2C_263_217),
	.V2C_7 (V2C_363_217),
	.V2C_8 (V2C_417_217),
	.V2C_9 (V2C_514_217),
	.V2C_10 (V2C_750_217),
	.V2C_11 (V2C_798_217),
	.V2C_12 (V2C_846_217),
	.V2C_13 (V2C_887_217),
	.V2C_14 (V2C_928_217),
	.V2C_15 (V2C_962_217),
	.V2C_16 (V2C_1049_217),
	.V2C_17 (V2C_1075_217),
	.V2C_18 (V2C_1134_217),
	.V2C_19 (V2C_1368_217),
	.V2C_20 (V2C_1369_217),
	.C2V_1 (C2V_217_41),
	.C2V_2 (C2V_217_77),
	.C2V_3 (C2V_217_97),
	.C2V_4 (C2V_217_158),
	.C2V_5 (C2V_217_220),
	.C2V_6 (C2V_217_263),
	.C2V_7 (C2V_217_363),
	.C2V_8 (C2V_217_417),
	.C2V_9 (C2V_217_514),
	.C2V_10 (C2V_217_750),
	.C2V_11 (C2V_217_798),
	.C2V_12 (C2V_217_846),
	.C2V_13 (C2V_217_887),
	.C2V_14 (C2V_217_928),
	.C2V_15 (C2V_217_962),
	.C2V_16 (C2V_217_1049),
	.C2V_17 (C2V_217_1075),
	.C2V_18 (C2V_217_1134),
	.C2V_19 (C2V_217_1368),
	.C2V_20 (C2V_217_1369),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU218 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_2_218),
	.V2C_2 (V2C_51_218),
	.V2C_3 (V2C_107_218),
	.V2C_4 (V2C_155_218),
	.V2C_5 (V2C_232_218),
	.V2C_6 (V2C_253_218),
	.V2C_7 (V2C_304_218),
	.V2C_8 (V2C_411_218),
	.V2C_9 (V2C_500_218),
	.V2C_10 (V2C_660_218),
	.V2C_11 (V2C_673_218),
	.V2C_12 (V2C_841_218),
	.V2C_13 (V2C_883_218),
	.V2C_14 (V2C_946_218),
	.V2C_15 (V2C_977_218),
	.V2C_16 (V2C_1009_218),
	.V2C_17 (V2C_1076_218),
	.V2C_18 (V2C_1107_218),
	.V2C_19 (V2C_1369_218),
	.V2C_20 (V2C_1370_218),
	.C2V_1 (C2V_218_2),
	.C2V_2 (C2V_218_51),
	.C2V_3 (C2V_218_107),
	.C2V_4 (C2V_218_155),
	.C2V_5 (C2V_218_232),
	.C2V_6 (C2V_218_253),
	.C2V_7 (C2V_218_304),
	.C2V_8 (C2V_218_411),
	.C2V_9 (C2V_218_500),
	.C2V_10 (C2V_218_660),
	.C2V_11 (C2V_218_673),
	.C2V_12 (C2V_218_841),
	.C2V_13 (C2V_218_883),
	.C2V_14 (C2V_218_946),
	.C2V_15 (C2V_218_977),
	.C2V_16 (C2V_218_1009),
	.C2V_17 (C2V_218_1076),
	.C2V_18 (C2V_218_1107),
	.C2V_19 (C2V_218_1369),
	.C2V_20 (C2V_218_1370),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU219 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_45_219),
	.V2C_2 (V2C_72_219),
	.V2C_3 (V2C_137_219),
	.V2C_4 (V2C_171_219),
	.V2C_5 (V2C_237_219),
	.V2C_6 (V2C_256_219),
	.V2C_7 (V2C_353_219),
	.V2C_8 (V2C_408_219),
	.V2C_9 (V2C_567_219),
	.V2C_10 (V2C_624_219),
	.V2C_11 (V2C_652_219),
	.V2C_12 (V2C_756_219),
	.V2C_13 (V2C_887_219),
	.V2C_14 (V2C_931_219),
	.V2C_15 (V2C_1004_219),
	.V2C_16 (V2C_1016_219),
	.V2C_17 (V2C_1094_219),
	.V2C_18 (V2C_1139_219),
	.V2C_19 (V2C_1370_219),
	.V2C_20 (V2C_1371_219),
	.C2V_1 (C2V_219_45),
	.C2V_2 (C2V_219_72),
	.C2V_3 (C2V_219_137),
	.C2V_4 (C2V_219_171),
	.C2V_5 (C2V_219_237),
	.C2V_6 (C2V_219_256),
	.C2V_7 (C2V_219_353),
	.C2V_8 (C2V_219_408),
	.C2V_9 (C2V_219_567),
	.C2V_10 (C2V_219_624),
	.C2V_11 (C2V_219_652),
	.C2V_12 (C2V_219_756),
	.C2V_13 (C2V_219_887),
	.C2V_14 (C2V_219_931),
	.C2V_15 (C2V_219_1004),
	.C2V_16 (C2V_219_1016),
	.C2V_17 (C2V_219_1094),
	.C2V_18 (C2V_219_1139),
	.C2V_19 (C2V_219_1370),
	.C2V_20 (C2V_219_1371),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU220 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_16_220),
	.V2C_2 (V2C_75_220),
	.V2C_3 (V2C_114_220),
	.V2C_4 (V2C_170_220),
	.V2C_5 (V2C_235_220),
	.V2C_6 (V2C_241_220),
	.V2C_7 (V2C_465_220),
	.V2C_8 (V2C_505_220),
	.V2C_9 (V2C_541_220),
	.V2C_10 (V2C_603_220),
	.V2C_11 (V2C_628_220),
	.V2C_12 (V2C_674_220),
	.V2C_13 (V2C_891_220),
	.V2C_14 (V2C_915_220),
	.V2C_15 (V2C_999_220),
	.V2C_16 (V2C_1029_220),
	.V2C_17 (V2C_1104_220),
	.V2C_18 (V2C_1120_220),
	.V2C_19 (V2C_1371_220),
	.V2C_20 (V2C_1372_220),
	.C2V_1 (C2V_220_16),
	.C2V_2 (C2V_220_75),
	.C2V_3 (C2V_220_114),
	.C2V_4 (C2V_220_170),
	.C2V_5 (C2V_220_235),
	.C2V_6 (C2V_220_241),
	.C2V_7 (C2V_220_465),
	.C2V_8 (C2V_220_505),
	.C2V_9 (C2V_220_541),
	.C2V_10 (C2V_220_603),
	.C2V_11 (C2V_220_628),
	.C2V_12 (C2V_220_674),
	.C2V_13 (C2V_220_891),
	.C2V_14 (C2V_220_915),
	.C2V_15 (C2V_220_999),
	.C2V_16 (C2V_220_1029),
	.C2V_17 (C2V_220_1104),
	.C2V_18 (C2V_220_1120),
	.C2V_19 (C2V_220_1371),
	.C2V_20 (C2V_220_1372),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU221 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_35_221),
	.V2C_2 (V2C_93_221),
	.V2C_3 (V2C_128_221),
	.V2C_4 (V2C_151_221),
	.V2C_5 (V2C_215_221),
	.V2C_6 (V2C_281_221),
	.V2C_7 (V2C_330_221),
	.V2C_8 (V2C_349_221),
	.V2C_9 (V2C_476_221),
	.V2C_10 (V2C_710_221),
	.V2C_11 (V2C_726_221),
	.V2C_12 (V2C_780_221),
	.V2C_13 (V2C_906_221),
	.V2C_14 (V2C_954_221),
	.V2C_15 (V2C_997_221),
	.V2C_16 (V2C_1049_221),
	.V2C_17 (V2C_1098_221),
	.V2C_18 (V2C_1146_221),
	.V2C_19 (V2C_1372_221),
	.V2C_20 (V2C_1373_221),
	.C2V_1 (C2V_221_35),
	.C2V_2 (C2V_221_93),
	.C2V_3 (C2V_221_128),
	.C2V_4 (C2V_221_151),
	.C2V_5 (C2V_221_215),
	.C2V_6 (C2V_221_281),
	.C2V_7 (C2V_221_330),
	.C2V_8 (C2V_221_349),
	.C2V_9 (C2V_221_476),
	.C2V_10 (C2V_221_710),
	.C2V_11 (C2V_221_726),
	.C2V_12 (C2V_221_780),
	.C2V_13 (C2V_221_906),
	.C2V_14 (C2V_221_954),
	.C2V_15 (C2V_221_997),
	.C2V_16 (C2V_221_1049),
	.C2V_17 (C2V_221_1098),
	.C2V_18 (C2V_221_1146),
	.C2V_19 (C2V_221_1372),
	.C2V_20 (C2V_221_1373),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU222 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_18_222),
	.V2C_2 (V2C_90_222),
	.V2C_3 (V2C_130_222),
	.V2C_4 (V2C_150_222),
	.V2C_5 (V2C_232_222),
	.V2C_6 (V2C_263_222),
	.V2C_7 (V2C_316_222),
	.V2C_8 (V2C_468_222),
	.V2C_9 (V2C_565_222),
	.V2C_10 (V2C_598_222),
	.V2C_11 (V2C_802_222),
	.V2C_12 (V2C_830_222),
	.V2C_13 (V2C_911_222),
	.V2C_14 (V2C_925_222),
	.V2C_15 (V2C_1008_222),
	.V2C_16 (V2C_1027_222),
	.V2C_17 (V2C_1091_222),
	.V2C_18 (V2C_1141_222),
	.V2C_19 (V2C_1373_222),
	.V2C_20 (V2C_1374_222),
	.C2V_1 (C2V_222_18),
	.C2V_2 (C2V_222_90),
	.C2V_3 (C2V_222_130),
	.C2V_4 (C2V_222_150),
	.C2V_5 (C2V_222_232),
	.C2V_6 (C2V_222_263),
	.C2V_7 (C2V_222_316),
	.C2V_8 (C2V_222_468),
	.C2V_9 (C2V_222_565),
	.C2V_10 (C2V_222_598),
	.C2V_11 (C2V_222_802),
	.C2V_12 (C2V_222_830),
	.C2V_13 (C2V_222_911),
	.C2V_14 (C2V_222_925),
	.C2V_15 (C2V_222_1008),
	.C2V_16 (C2V_222_1027),
	.C2V_17 (C2V_222_1091),
	.C2V_18 (C2V_222_1141),
	.C2V_19 (C2V_222_1373),
	.C2V_20 (C2V_222_1374),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU223 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_42_223),
	.V2C_2 (V2C_78_223),
	.V2C_3 (V2C_98_223),
	.V2C_4 (V2C_159_223),
	.V2C_5 (V2C_221_223),
	.V2C_6 (V2C_264_223),
	.V2C_7 (V2C_364_223),
	.V2C_8 (V2C_418_223),
	.V2C_9 (V2C_515_223),
	.V2C_10 (V2C_751_223),
	.V2C_11 (V2C_799_223),
	.V2C_12 (V2C_847_223),
	.V2C_13 (V2C_888_223),
	.V2C_14 (V2C_929_223),
	.V2C_15 (V2C_963_223),
	.V2C_16 (V2C_1050_223),
	.V2C_17 (V2C_1076_223),
	.V2C_18 (V2C_1135_223),
	.V2C_19 (V2C_1374_223),
	.V2C_20 (V2C_1375_223),
	.C2V_1 (C2V_223_42),
	.C2V_2 (C2V_223_78),
	.C2V_3 (C2V_223_98),
	.C2V_4 (C2V_223_159),
	.C2V_5 (C2V_223_221),
	.C2V_6 (C2V_223_264),
	.C2V_7 (C2V_223_364),
	.C2V_8 (C2V_223_418),
	.C2V_9 (C2V_223_515),
	.C2V_10 (C2V_223_751),
	.C2V_11 (C2V_223_799),
	.C2V_12 (C2V_223_847),
	.C2V_13 (C2V_223_888),
	.C2V_14 (C2V_223_929),
	.C2V_15 (C2V_223_963),
	.C2V_16 (C2V_223_1050),
	.C2V_17 (C2V_223_1076),
	.C2V_18 (C2V_223_1135),
	.C2V_19 (C2V_223_1374),
	.C2V_20 (C2V_223_1375),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU224 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_3_224),
	.V2C_2 (V2C_52_224),
	.V2C_3 (V2C_108_224),
	.V2C_4 (V2C_156_224),
	.V2C_5 (V2C_233_224),
	.V2C_6 (V2C_254_224),
	.V2C_7 (V2C_305_224),
	.V2C_8 (V2C_412_224),
	.V2C_9 (V2C_501_224),
	.V2C_10 (V2C_661_224),
	.V2C_11 (V2C_674_224),
	.V2C_12 (V2C_842_224),
	.V2C_13 (V2C_884_224),
	.V2C_14 (V2C_947_224),
	.V2C_15 (V2C_978_224),
	.V2C_16 (V2C_1010_224),
	.V2C_17 (V2C_1077_224),
	.V2C_18 (V2C_1108_224),
	.V2C_19 (V2C_1375_224),
	.V2C_20 (V2C_1376_224),
	.C2V_1 (C2V_224_3),
	.C2V_2 (C2V_224_52),
	.C2V_3 (C2V_224_108),
	.C2V_4 (C2V_224_156),
	.C2V_5 (C2V_224_233),
	.C2V_6 (C2V_224_254),
	.C2V_7 (C2V_224_305),
	.C2V_8 (C2V_224_412),
	.C2V_9 (C2V_224_501),
	.C2V_10 (C2V_224_661),
	.C2V_11 (C2V_224_674),
	.C2V_12 (C2V_224_842),
	.C2V_13 (C2V_224_884),
	.C2V_14 (C2V_224_947),
	.C2V_15 (C2V_224_978),
	.C2V_16 (C2V_224_1010),
	.C2V_17 (C2V_224_1077),
	.C2V_18 (C2V_224_1108),
	.C2V_19 (C2V_224_1375),
	.C2V_20 (C2V_224_1376),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU225 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_46_225),
	.V2C_2 (V2C_73_225),
	.V2C_3 (V2C_138_225),
	.V2C_4 (V2C_172_225),
	.V2C_5 (V2C_238_225),
	.V2C_6 (V2C_257_225),
	.V2C_7 (V2C_354_225),
	.V2C_8 (V2C_409_225),
	.V2C_9 (V2C_568_225),
	.V2C_10 (V2C_577_225),
	.V2C_11 (V2C_653_225),
	.V2C_12 (V2C_757_225),
	.V2C_13 (V2C_888_225),
	.V2C_14 (V2C_932_225),
	.V2C_15 (V2C_1005_225),
	.V2C_16 (V2C_1017_225),
	.V2C_17 (V2C_1095_225),
	.V2C_18 (V2C_1140_225),
	.V2C_19 (V2C_1376_225),
	.V2C_20 (V2C_1377_225),
	.C2V_1 (C2V_225_46),
	.C2V_2 (C2V_225_73),
	.C2V_3 (C2V_225_138),
	.C2V_4 (C2V_225_172),
	.C2V_5 (C2V_225_238),
	.C2V_6 (C2V_225_257),
	.C2V_7 (C2V_225_354),
	.C2V_8 (C2V_225_409),
	.C2V_9 (C2V_225_568),
	.C2V_10 (C2V_225_577),
	.C2V_11 (C2V_225_653),
	.C2V_12 (C2V_225_757),
	.C2V_13 (C2V_225_888),
	.C2V_14 (C2V_225_932),
	.C2V_15 (C2V_225_1005),
	.C2V_16 (C2V_225_1017),
	.C2V_17 (C2V_225_1095),
	.C2V_18 (C2V_225_1140),
	.C2V_19 (C2V_225_1376),
	.C2V_20 (C2V_225_1377),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU226 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_17_226),
	.V2C_2 (V2C_76_226),
	.V2C_3 (V2C_115_226),
	.V2C_4 (V2C_171_226),
	.V2C_5 (V2C_236_226),
	.V2C_6 (V2C_242_226),
	.V2C_7 (V2C_466_226),
	.V2C_8 (V2C_506_226),
	.V2C_9 (V2C_542_226),
	.V2C_10 (V2C_604_226),
	.V2C_11 (V2C_629_226),
	.V2C_12 (V2C_675_226),
	.V2C_13 (V2C_892_226),
	.V2C_14 (V2C_916_226),
	.V2C_15 (V2C_1000_226),
	.V2C_16 (V2C_1030_226),
	.V2C_17 (V2C_1057_226),
	.V2C_18 (V2C_1121_226),
	.V2C_19 (V2C_1377_226),
	.V2C_20 (V2C_1378_226),
	.C2V_1 (C2V_226_17),
	.C2V_2 (C2V_226_76),
	.C2V_3 (C2V_226_115),
	.C2V_4 (C2V_226_171),
	.C2V_5 (C2V_226_236),
	.C2V_6 (C2V_226_242),
	.C2V_7 (C2V_226_466),
	.C2V_8 (C2V_226_506),
	.C2V_9 (C2V_226_542),
	.C2V_10 (C2V_226_604),
	.C2V_11 (C2V_226_629),
	.C2V_12 (C2V_226_675),
	.C2V_13 (C2V_226_892),
	.C2V_14 (C2V_226_916),
	.C2V_15 (C2V_226_1000),
	.C2V_16 (C2V_226_1030),
	.C2V_17 (C2V_226_1057),
	.C2V_18 (C2V_226_1121),
	.C2V_19 (C2V_226_1377),
	.C2V_20 (C2V_226_1378),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU227 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_36_227),
	.V2C_2 (V2C_94_227),
	.V2C_3 (V2C_129_227),
	.V2C_4 (V2C_152_227),
	.V2C_5 (V2C_216_227),
	.V2C_6 (V2C_282_227),
	.V2C_7 (V2C_331_227),
	.V2C_8 (V2C_350_227),
	.V2C_9 (V2C_477_227),
	.V2C_10 (V2C_711_227),
	.V2C_11 (V2C_727_227),
	.V2C_12 (V2C_781_227),
	.V2C_13 (V2C_907_227),
	.V2C_14 (V2C_955_227),
	.V2C_15 (V2C_998_227),
	.V2C_16 (V2C_1050_227),
	.V2C_17 (V2C_1099_227),
	.V2C_18 (V2C_1147_227),
	.V2C_19 (V2C_1378_227),
	.V2C_20 (V2C_1379_227),
	.C2V_1 (C2V_227_36),
	.C2V_2 (C2V_227_94),
	.C2V_3 (C2V_227_129),
	.C2V_4 (C2V_227_152),
	.C2V_5 (C2V_227_216),
	.C2V_6 (C2V_227_282),
	.C2V_7 (C2V_227_331),
	.C2V_8 (C2V_227_350),
	.C2V_9 (C2V_227_477),
	.C2V_10 (C2V_227_711),
	.C2V_11 (C2V_227_727),
	.C2V_12 (C2V_227_781),
	.C2V_13 (C2V_227_907),
	.C2V_14 (C2V_227_955),
	.C2V_15 (C2V_227_998),
	.C2V_16 (C2V_227_1050),
	.C2V_17 (C2V_227_1099),
	.C2V_18 (C2V_227_1147),
	.C2V_19 (C2V_227_1378),
	.C2V_20 (C2V_227_1379),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU228 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_19_228),
	.V2C_2 (V2C_91_228),
	.V2C_3 (V2C_131_228),
	.V2C_4 (V2C_151_228),
	.V2C_5 (V2C_233_228),
	.V2C_6 (V2C_264_228),
	.V2C_7 (V2C_317_228),
	.V2C_8 (V2C_469_228),
	.V2C_9 (V2C_566_228),
	.V2C_10 (V2C_599_228),
	.V2C_11 (V2C_803_228),
	.V2C_12 (V2C_831_228),
	.V2C_13 (V2C_912_228),
	.V2C_14 (V2C_926_228),
	.V2C_15 (V2C_961_228),
	.V2C_16 (V2C_1028_228),
	.V2C_17 (V2C_1092_228),
	.V2C_18 (V2C_1142_228),
	.V2C_19 (V2C_1379_228),
	.V2C_20 (V2C_1380_228),
	.C2V_1 (C2V_228_19),
	.C2V_2 (C2V_228_91),
	.C2V_3 (C2V_228_131),
	.C2V_4 (C2V_228_151),
	.C2V_5 (C2V_228_233),
	.C2V_6 (C2V_228_264),
	.C2V_7 (C2V_228_317),
	.C2V_8 (C2V_228_469),
	.C2V_9 (C2V_228_566),
	.C2V_10 (C2V_228_599),
	.C2V_11 (C2V_228_803),
	.C2V_12 (C2V_228_831),
	.C2V_13 (C2V_228_912),
	.C2V_14 (C2V_228_926),
	.C2V_15 (C2V_228_961),
	.C2V_16 (C2V_228_1028),
	.C2V_17 (C2V_228_1092),
	.C2V_18 (C2V_228_1142),
	.C2V_19 (C2V_228_1379),
	.C2V_20 (C2V_228_1380),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU229 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_43_229),
	.V2C_2 (V2C_79_229),
	.V2C_3 (V2C_99_229),
	.V2C_4 (V2C_160_229),
	.V2C_5 (V2C_222_229),
	.V2C_6 (V2C_265_229),
	.V2C_7 (V2C_365_229),
	.V2C_8 (V2C_419_229),
	.V2C_9 (V2C_516_229),
	.V2C_10 (V2C_752_229),
	.V2C_11 (V2C_800_229),
	.V2C_12 (V2C_848_229),
	.V2C_13 (V2C_889_229),
	.V2C_14 (V2C_930_229),
	.V2C_15 (V2C_964_229),
	.V2C_16 (V2C_1051_229),
	.V2C_17 (V2C_1077_229),
	.V2C_18 (V2C_1136_229),
	.V2C_19 (V2C_1380_229),
	.V2C_20 (V2C_1381_229),
	.C2V_1 (C2V_229_43),
	.C2V_2 (C2V_229_79),
	.C2V_3 (C2V_229_99),
	.C2V_4 (C2V_229_160),
	.C2V_5 (C2V_229_222),
	.C2V_6 (C2V_229_265),
	.C2V_7 (C2V_229_365),
	.C2V_8 (C2V_229_419),
	.C2V_9 (C2V_229_516),
	.C2V_10 (C2V_229_752),
	.C2V_11 (C2V_229_800),
	.C2V_12 (C2V_229_848),
	.C2V_13 (C2V_229_889),
	.C2V_14 (C2V_229_930),
	.C2V_15 (C2V_229_964),
	.C2V_16 (C2V_229_1051),
	.C2V_17 (C2V_229_1077),
	.C2V_18 (C2V_229_1136),
	.C2V_19 (C2V_229_1380),
	.C2V_20 (C2V_229_1381),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU230 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_4_230),
	.V2C_2 (V2C_53_230),
	.V2C_3 (V2C_109_230),
	.V2C_4 (V2C_157_230),
	.V2C_5 (V2C_234_230),
	.V2C_6 (V2C_255_230),
	.V2C_7 (V2C_306_230),
	.V2C_8 (V2C_413_230),
	.V2C_9 (V2C_502_230),
	.V2C_10 (V2C_662_230),
	.V2C_11 (V2C_675_230),
	.V2C_12 (V2C_843_230),
	.V2C_13 (V2C_885_230),
	.V2C_14 (V2C_948_230),
	.V2C_15 (V2C_979_230),
	.V2C_16 (V2C_1011_230),
	.V2C_17 (V2C_1078_230),
	.V2C_18 (V2C_1109_230),
	.V2C_19 (V2C_1381_230),
	.V2C_20 (V2C_1382_230),
	.C2V_1 (C2V_230_4),
	.C2V_2 (C2V_230_53),
	.C2V_3 (C2V_230_109),
	.C2V_4 (C2V_230_157),
	.C2V_5 (C2V_230_234),
	.C2V_6 (C2V_230_255),
	.C2V_7 (C2V_230_306),
	.C2V_8 (C2V_230_413),
	.C2V_9 (C2V_230_502),
	.C2V_10 (C2V_230_662),
	.C2V_11 (C2V_230_675),
	.C2V_12 (C2V_230_843),
	.C2V_13 (C2V_230_885),
	.C2V_14 (C2V_230_948),
	.C2V_15 (C2V_230_979),
	.C2V_16 (C2V_230_1011),
	.C2V_17 (C2V_230_1078),
	.C2V_18 (C2V_230_1109),
	.C2V_19 (C2V_230_1381),
	.C2V_20 (C2V_230_1382),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU231 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_47_231),
	.V2C_2 (V2C_74_231),
	.V2C_3 (V2C_139_231),
	.V2C_4 (V2C_173_231),
	.V2C_5 (V2C_239_231),
	.V2C_6 (V2C_258_231),
	.V2C_7 (V2C_355_231),
	.V2C_8 (V2C_410_231),
	.V2C_9 (V2C_569_231),
	.V2C_10 (V2C_578_231),
	.V2C_11 (V2C_654_231),
	.V2C_12 (V2C_758_231),
	.V2C_13 (V2C_889_231),
	.V2C_14 (V2C_933_231),
	.V2C_15 (V2C_1006_231),
	.V2C_16 (V2C_1018_231),
	.V2C_17 (V2C_1096_231),
	.V2C_18 (V2C_1141_231),
	.V2C_19 (V2C_1382_231),
	.V2C_20 (V2C_1383_231),
	.C2V_1 (C2V_231_47),
	.C2V_2 (C2V_231_74),
	.C2V_3 (C2V_231_139),
	.C2V_4 (C2V_231_173),
	.C2V_5 (C2V_231_239),
	.C2V_6 (C2V_231_258),
	.C2V_7 (C2V_231_355),
	.C2V_8 (C2V_231_410),
	.C2V_9 (C2V_231_569),
	.C2V_10 (C2V_231_578),
	.C2V_11 (C2V_231_654),
	.C2V_12 (C2V_231_758),
	.C2V_13 (C2V_231_889),
	.C2V_14 (C2V_231_933),
	.C2V_15 (C2V_231_1006),
	.C2V_16 (C2V_231_1018),
	.C2V_17 (C2V_231_1096),
	.C2V_18 (C2V_231_1141),
	.C2V_19 (C2V_231_1382),
	.C2V_20 (C2V_231_1383),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU232 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_18_232),
	.V2C_2 (V2C_77_232),
	.V2C_3 (V2C_116_232),
	.V2C_4 (V2C_172_232),
	.V2C_5 (V2C_237_232),
	.V2C_6 (V2C_243_232),
	.V2C_7 (V2C_467_232),
	.V2C_8 (V2C_507_232),
	.V2C_9 (V2C_543_232),
	.V2C_10 (V2C_605_232),
	.V2C_11 (V2C_630_232),
	.V2C_12 (V2C_676_232),
	.V2C_13 (V2C_893_232),
	.V2C_14 (V2C_917_232),
	.V2C_15 (V2C_1001_232),
	.V2C_16 (V2C_1031_232),
	.V2C_17 (V2C_1058_232),
	.V2C_18 (V2C_1122_232),
	.V2C_19 (V2C_1383_232),
	.V2C_20 (V2C_1384_232),
	.C2V_1 (C2V_232_18),
	.C2V_2 (C2V_232_77),
	.C2V_3 (C2V_232_116),
	.C2V_4 (C2V_232_172),
	.C2V_5 (C2V_232_237),
	.C2V_6 (C2V_232_243),
	.C2V_7 (C2V_232_467),
	.C2V_8 (C2V_232_507),
	.C2V_9 (C2V_232_543),
	.C2V_10 (C2V_232_605),
	.C2V_11 (C2V_232_630),
	.C2V_12 (C2V_232_676),
	.C2V_13 (C2V_232_893),
	.C2V_14 (C2V_232_917),
	.C2V_15 (C2V_232_1001),
	.C2V_16 (C2V_232_1031),
	.C2V_17 (C2V_232_1058),
	.C2V_18 (C2V_232_1122),
	.C2V_19 (C2V_232_1383),
	.C2V_20 (C2V_232_1384),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU233 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_37_233),
	.V2C_2 (V2C_95_233),
	.V2C_3 (V2C_130_233),
	.V2C_4 (V2C_153_233),
	.V2C_5 (V2C_217_233),
	.V2C_6 (V2C_283_233),
	.V2C_7 (V2C_332_233),
	.V2C_8 (V2C_351_233),
	.V2C_9 (V2C_478_233),
	.V2C_10 (V2C_712_233),
	.V2C_11 (V2C_728_233),
	.V2C_12 (V2C_782_233),
	.V2C_13 (V2C_908_233),
	.V2C_14 (V2C_956_233),
	.V2C_15 (V2C_999_233),
	.V2C_16 (V2C_1051_233),
	.V2C_17 (V2C_1100_233),
	.V2C_18 (V2C_1148_233),
	.V2C_19 (V2C_1384_233),
	.V2C_20 (V2C_1385_233),
	.C2V_1 (C2V_233_37),
	.C2V_2 (C2V_233_95),
	.C2V_3 (C2V_233_130),
	.C2V_4 (C2V_233_153),
	.C2V_5 (C2V_233_217),
	.C2V_6 (C2V_233_283),
	.C2V_7 (C2V_233_332),
	.C2V_8 (C2V_233_351),
	.C2V_9 (C2V_233_478),
	.C2V_10 (C2V_233_712),
	.C2V_11 (C2V_233_728),
	.C2V_12 (C2V_233_782),
	.C2V_13 (C2V_233_908),
	.C2V_14 (C2V_233_956),
	.C2V_15 (C2V_233_999),
	.C2V_16 (C2V_233_1051),
	.C2V_17 (C2V_233_1100),
	.C2V_18 (C2V_233_1148),
	.C2V_19 (C2V_233_1384),
	.C2V_20 (C2V_233_1385),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU234 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_20_234),
	.V2C_2 (V2C_92_234),
	.V2C_3 (V2C_132_234),
	.V2C_4 (V2C_152_234),
	.V2C_5 (V2C_234_234),
	.V2C_6 (V2C_265_234),
	.V2C_7 (V2C_318_234),
	.V2C_8 (V2C_470_234),
	.V2C_9 (V2C_567_234),
	.V2C_10 (V2C_600_234),
	.V2C_11 (V2C_804_234),
	.V2C_12 (V2C_832_234),
	.V2C_13 (V2C_865_234),
	.V2C_14 (V2C_927_234),
	.V2C_15 (V2C_962_234),
	.V2C_16 (V2C_1029_234),
	.V2C_17 (V2C_1093_234),
	.V2C_18 (V2C_1143_234),
	.V2C_19 (V2C_1385_234),
	.V2C_20 (V2C_1386_234),
	.C2V_1 (C2V_234_20),
	.C2V_2 (C2V_234_92),
	.C2V_3 (C2V_234_132),
	.C2V_4 (C2V_234_152),
	.C2V_5 (C2V_234_234),
	.C2V_6 (C2V_234_265),
	.C2V_7 (C2V_234_318),
	.C2V_8 (C2V_234_470),
	.C2V_9 (C2V_234_567),
	.C2V_10 (C2V_234_600),
	.C2V_11 (C2V_234_804),
	.C2V_12 (C2V_234_832),
	.C2V_13 (C2V_234_865),
	.C2V_14 (C2V_234_927),
	.C2V_15 (C2V_234_962),
	.C2V_16 (C2V_234_1029),
	.C2V_17 (C2V_234_1093),
	.C2V_18 (C2V_234_1143),
	.C2V_19 (C2V_234_1385),
	.C2V_20 (C2V_234_1386),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU235 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_44_235),
	.V2C_2 (V2C_80_235),
	.V2C_3 (V2C_100_235),
	.V2C_4 (V2C_161_235),
	.V2C_5 (V2C_223_235),
	.V2C_6 (V2C_266_235),
	.V2C_7 (V2C_366_235),
	.V2C_8 (V2C_420_235),
	.V2C_9 (V2C_517_235),
	.V2C_10 (V2C_753_235),
	.V2C_11 (V2C_801_235),
	.V2C_12 (V2C_849_235),
	.V2C_13 (V2C_890_235),
	.V2C_14 (V2C_931_235),
	.V2C_15 (V2C_965_235),
	.V2C_16 (V2C_1052_235),
	.V2C_17 (V2C_1078_235),
	.V2C_18 (V2C_1137_235),
	.V2C_19 (V2C_1386_235),
	.V2C_20 (V2C_1387_235),
	.C2V_1 (C2V_235_44),
	.C2V_2 (C2V_235_80),
	.C2V_3 (C2V_235_100),
	.C2V_4 (C2V_235_161),
	.C2V_5 (C2V_235_223),
	.C2V_6 (C2V_235_266),
	.C2V_7 (C2V_235_366),
	.C2V_8 (C2V_235_420),
	.C2V_9 (C2V_235_517),
	.C2V_10 (C2V_235_753),
	.C2V_11 (C2V_235_801),
	.C2V_12 (C2V_235_849),
	.C2V_13 (C2V_235_890),
	.C2V_14 (C2V_235_931),
	.C2V_15 (C2V_235_965),
	.C2V_16 (C2V_235_1052),
	.C2V_17 (C2V_235_1078),
	.C2V_18 (C2V_235_1137),
	.C2V_19 (C2V_235_1386),
	.C2V_20 (C2V_235_1387),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU236 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_5_236),
	.V2C_2 (V2C_54_236),
	.V2C_3 (V2C_110_236),
	.V2C_4 (V2C_158_236),
	.V2C_5 (V2C_235_236),
	.V2C_6 (V2C_256_236),
	.V2C_7 (V2C_307_236),
	.V2C_8 (V2C_414_236),
	.V2C_9 (V2C_503_236),
	.V2C_10 (V2C_663_236),
	.V2C_11 (V2C_676_236),
	.V2C_12 (V2C_844_236),
	.V2C_13 (V2C_886_236),
	.V2C_14 (V2C_949_236),
	.V2C_15 (V2C_980_236),
	.V2C_16 (V2C_1012_236),
	.V2C_17 (V2C_1079_236),
	.V2C_18 (V2C_1110_236),
	.V2C_19 (V2C_1387_236),
	.V2C_20 (V2C_1388_236),
	.C2V_1 (C2V_236_5),
	.C2V_2 (C2V_236_54),
	.C2V_3 (C2V_236_110),
	.C2V_4 (C2V_236_158),
	.C2V_5 (C2V_236_235),
	.C2V_6 (C2V_236_256),
	.C2V_7 (C2V_236_307),
	.C2V_8 (C2V_236_414),
	.C2V_9 (C2V_236_503),
	.C2V_10 (C2V_236_663),
	.C2V_11 (C2V_236_676),
	.C2V_12 (C2V_236_844),
	.C2V_13 (C2V_236_886),
	.C2V_14 (C2V_236_949),
	.C2V_15 (C2V_236_980),
	.C2V_16 (C2V_236_1012),
	.C2V_17 (C2V_236_1079),
	.C2V_18 (C2V_236_1110),
	.C2V_19 (C2V_236_1387),
	.C2V_20 (C2V_236_1388),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU237 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_48_237),
	.V2C_2 (V2C_75_237),
	.V2C_3 (V2C_140_237),
	.V2C_4 (V2C_174_237),
	.V2C_5 (V2C_240_237),
	.V2C_6 (V2C_259_237),
	.V2C_7 (V2C_356_237),
	.V2C_8 (V2C_411_237),
	.V2C_9 (V2C_570_237),
	.V2C_10 (V2C_579_237),
	.V2C_11 (V2C_655_237),
	.V2C_12 (V2C_759_237),
	.V2C_13 (V2C_890_237),
	.V2C_14 (V2C_934_237),
	.V2C_15 (V2C_1007_237),
	.V2C_16 (V2C_1019_237),
	.V2C_17 (V2C_1097_237),
	.V2C_18 (V2C_1142_237),
	.V2C_19 (V2C_1388_237),
	.V2C_20 (V2C_1389_237),
	.C2V_1 (C2V_237_48),
	.C2V_2 (C2V_237_75),
	.C2V_3 (C2V_237_140),
	.C2V_4 (C2V_237_174),
	.C2V_5 (C2V_237_240),
	.C2V_6 (C2V_237_259),
	.C2V_7 (C2V_237_356),
	.C2V_8 (C2V_237_411),
	.C2V_9 (C2V_237_570),
	.C2V_10 (C2V_237_579),
	.C2V_11 (C2V_237_655),
	.C2V_12 (C2V_237_759),
	.C2V_13 (C2V_237_890),
	.C2V_14 (C2V_237_934),
	.C2V_15 (C2V_237_1007),
	.C2V_16 (C2V_237_1019),
	.C2V_17 (C2V_237_1097),
	.C2V_18 (C2V_237_1142),
	.C2V_19 (C2V_237_1388),
	.C2V_20 (C2V_237_1389),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU238 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_19_238),
	.V2C_2 (V2C_78_238),
	.V2C_3 (V2C_117_238),
	.V2C_4 (V2C_173_238),
	.V2C_5 (V2C_238_238),
	.V2C_6 (V2C_244_238),
	.V2C_7 (V2C_468_238),
	.V2C_8 (V2C_508_238),
	.V2C_9 (V2C_544_238),
	.V2C_10 (V2C_606_238),
	.V2C_11 (V2C_631_238),
	.V2C_12 (V2C_677_238),
	.V2C_13 (V2C_894_238),
	.V2C_14 (V2C_918_238),
	.V2C_15 (V2C_1002_238),
	.V2C_16 (V2C_1032_238),
	.V2C_17 (V2C_1059_238),
	.V2C_18 (V2C_1123_238),
	.V2C_19 (V2C_1389_238),
	.V2C_20 (V2C_1390_238),
	.C2V_1 (C2V_238_19),
	.C2V_2 (C2V_238_78),
	.C2V_3 (C2V_238_117),
	.C2V_4 (C2V_238_173),
	.C2V_5 (C2V_238_238),
	.C2V_6 (C2V_238_244),
	.C2V_7 (C2V_238_468),
	.C2V_8 (C2V_238_508),
	.C2V_9 (C2V_238_544),
	.C2V_10 (C2V_238_606),
	.C2V_11 (C2V_238_631),
	.C2V_12 (C2V_238_677),
	.C2V_13 (C2V_238_894),
	.C2V_14 (C2V_238_918),
	.C2V_15 (C2V_238_1002),
	.C2V_16 (C2V_238_1032),
	.C2V_17 (C2V_238_1059),
	.C2V_18 (C2V_238_1123),
	.C2V_19 (C2V_238_1389),
	.C2V_20 (C2V_238_1390),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU239 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_38_239),
	.V2C_2 (V2C_96_239),
	.V2C_3 (V2C_131_239),
	.V2C_4 (V2C_154_239),
	.V2C_5 (V2C_218_239),
	.V2C_6 (V2C_284_239),
	.V2C_7 (V2C_333_239),
	.V2C_8 (V2C_352_239),
	.V2C_9 (V2C_479_239),
	.V2C_10 (V2C_713_239),
	.V2C_11 (V2C_729_239),
	.V2C_12 (V2C_783_239),
	.V2C_13 (V2C_909_239),
	.V2C_14 (V2C_957_239),
	.V2C_15 (V2C_1000_239),
	.V2C_16 (V2C_1052_239),
	.V2C_17 (V2C_1101_239),
	.V2C_18 (V2C_1149_239),
	.V2C_19 (V2C_1390_239),
	.V2C_20 (V2C_1391_239),
	.C2V_1 (C2V_239_38),
	.C2V_2 (C2V_239_96),
	.C2V_3 (C2V_239_131),
	.C2V_4 (C2V_239_154),
	.C2V_5 (C2V_239_218),
	.C2V_6 (C2V_239_284),
	.C2V_7 (C2V_239_333),
	.C2V_8 (C2V_239_352),
	.C2V_9 (C2V_239_479),
	.C2V_10 (C2V_239_713),
	.C2V_11 (C2V_239_729),
	.C2V_12 (C2V_239_783),
	.C2V_13 (C2V_239_909),
	.C2V_14 (C2V_239_957),
	.C2V_15 (C2V_239_1000),
	.C2V_16 (C2V_239_1052),
	.C2V_17 (C2V_239_1101),
	.C2V_18 (C2V_239_1149),
	.C2V_19 (C2V_239_1390),
	.C2V_20 (C2V_239_1391),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU240 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_21_240),
	.V2C_2 (V2C_93_240),
	.V2C_3 (V2C_133_240),
	.V2C_4 (V2C_153_240),
	.V2C_5 (V2C_235_240),
	.V2C_6 (V2C_266_240),
	.V2C_7 (V2C_319_240),
	.V2C_8 (V2C_471_240),
	.V2C_9 (V2C_568_240),
	.V2C_10 (V2C_601_240),
	.V2C_11 (V2C_805_240),
	.V2C_12 (V2C_833_240),
	.V2C_13 (V2C_866_240),
	.V2C_14 (V2C_928_240),
	.V2C_15 (V2C_963_240),
	.V2C_16 (V2C_1030_240),
	.V2C_17 (V2C_1094_240),
	.V2C_18 (V2C_1144_240),
	.V2C_19 (V2C_1391_240),
	.V2C_20 (V2C_1392_240),
	.C2V_1 (C2V_240_21),
	.C2V_2 (C2V_240_93),
	.C2V_3 (C2V_240_133),
	.C2V_4 (C2V_240_153),
	.C2V_5 (C2V_240_235),
	.C2V_6 (C2V_240_266),
	.C2V_7 (C2V_240_319),
	.C2V_8 (C2V_240_471),
	.C2V_9 (C2V_240_568),
	.C2V_10 (C2V_240_601),
	.C2V_11 (C2V_240_805),
	.C2V_12 (C2V_240_833),
	.C2V_13 (C2V_240_866),
	.C2V_14 (C2V_240_928),
	.C2V_15 (C2V_240_963),
	.C2V_16 (C2V_240_1030),
	.C2V_17 (C2V_240_1094),
	.C2V_18 (C2V_240_1144),
	.C2V_19 (C2V_240_1391),
	.C2V_20 (C2V_240_1392),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU241 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_45_241),
	.V2C_2 (V2C_81_241),
	.V2C_3 (V2C_101_241),
	.V2C_4 (V2C_162_241),
	.V2C_5 (V2C_224_241),
	.V2C_6 (V2C_267_241),
	.V2C_7 (V2C_367_241),
	.V2C_8 (V2C_421_241),
	.V2C_9 (V2C_518_241),
	.V2C_10 (V2C_754_241),
	.V2C_11 (V2C_802_241),
	.V2C_12 (V2C_850_241),
	.V2C_13 (V2C_891_241),
	.V2C_14 (V2C_932_241),
	.V2C_15 (V2C_966_241),
	.V2C_16 (V2C_1053_241),
	.V2C_17 (V2C_1079_241),
	.V2C_18 (V2C_1138_241),
	.V2C_19 (V2C_1392_241),
	.V2C_20 (V2C_1393_241),
	.C2V_1 (C2V_241_45),
	.C2V_2 (C2V_241_81),
	.C2V_3 (C2V_241_101),
	.C2V_4 (C2V_241_162),
	.C2V_5 (C2V_241_224),
	.C2V_6 (C2V_241_267),
	.C2V_7 (C2V_241_367),
	.C2V_8 (C2V_241_421),
	.C2V_9 (C2V_241_518),
	.C2V_10 (C2V_241_754),
	.C2V_11 (C2V_241_802),
	.C2V_12 (C2V_241_850),
	.C2V_13 (C2V_241_891),
	.C2V_14 (C2V_241_932),
	.C2V_15 (C2V_241_966),
	.C2V_16 (C2V_241_1053),
	.C2V_17 (C2V_241_1079),
	.C2V_18 (C2V_241_1138),
	.C2V_19 (C2V_241_1392),
	.C2V_20 (C2V_241_1393),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU242 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_6_242),
	.V2C_2 (V2C_55_242),
	.V2C_3 (V2C_111_242),
	.V2C_4 (V2C_159_242),
	.V2C_5 (V2C_236_242),
	.V2C_6 (V2C_257_242),
	.V2C_7 (V2C_308_242),
	.V2C_8 (V2C_415_242),
	.V2C_9 (V2C_504_242),
	.V2C_10 (V2C_664_242),
	.V2C_11 (V2C_677_242),
	.V2C_12 (V2C_845_242),
	.V2C_13 (V2C_887_242),
	.V2C_14 (V2C_950_242),
	.V2C_15 (V2C_981_242),
	.V2C_16 (V2C_1013_242),
	.V2C_17 (V2C_1080_242),
	.V2C_18 (V2C_1111_242),
	.V2C_19 (V2C_1393_242),
	.V2C_20 (V2C_1394_242),
	.C2V_1 (C2V_242_6),
	.C2V_2 (C2V_242_55),
	.C2V_3 (C2V_242_111),
	.C2V_4 (C2V_242_159),
	.C2V_5 (C2V_242_236),
	.C2V_6 (C2V_242_257),
	.C2V_7 (C2V_242_308),
	.C2V_8 (C2V_242_415),
	.C2V_9 (C2V_242_504),
	.C2V_10 (C2V_242_664),
	.C2V_11 (C2V_242_677),
	.C2V_12 (C2V_242_845),
	.C2V_13 (C2V_242_887),
	.C2V_14 (C2V_242_950),
	.C2V_15 (C2V_242_981),
	.C2V_16 (C2V_242_1013),
	.C2V_17 (C2V_242_1080),
	.C2V_18 (C2V_242_1111),
	.C2V_19 (C2V_242_1393),
	.C2V_20 (C2V_242_1394),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU243 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_1_243),
	.V2C_2 (V2C_76_243),
	.V2C_3 (V2C_141_243),
	.V2C_4 (V2C_175_243),
	.V2C_5 (V2C_193_243),
	.V2C_6 (V2C_260_243),
	.V2C_7 (V2C_357_243),
	.V2C_8 (V2C_412_243),
	.V2C_9 (V2C_571_243),
	.V2C_10 (V2C_580_243),
	.V2C_11 (V2C_656_243),
	.V2C_12 (V2C_760_243),
	.V2C_13 (V2C_891_243),
	.V2C_14 (V2C_935_243),
	.V2C_15 (V2C_1008_243),
	.V2C_16 (V2C_1020_243),
	.V2C_17 (V2C_1098_243),
	.V2C_18 (V2C_1143_243),
	.V2C_19 (V2C_1394_243),
	.V2C_20 (V2C_1395_243),
	.C2V_1 (C2V_243_1),
	.C2V_2 (C2V_243_76),
	.C2V_3 (C2V_243_141),
	.C2V_4 (C2V_243_175),
	.C2V_5 (C2V_243_193),
	.C2V_6 (C2V_243_260),
	.C2V_7 (C2V_243_357),
	.C2V_8 (C2V_243_412),
	.C2V_9 (C2V_243_571),
	.C2V_10 (C2V_243_580),
	.C2V_11 (C2V_243_656),
	.C2V_12 (C2V_243_760),
	.C2V_13 (C2V_243_891),
	.C2V_14 (C2V_243_935),
	.C2V_15 (C2V_243_1008),
	.C2V_16 (C2V_243_1020),
	.C2V_17 (C2V_243_1098),
	.C2V_18 (C2V_243_1143),
	.C2V_19 (C2V_243_1394),
	.C2V_20 (C2V_243_1395),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU244 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_20_244),
	.V2C_2 (V2C_79_244),
	.V2C_3 (V2C_118_244),
	.V2C_4 (V2C_174_244),
	.V2C_5 (V2C_239_244),
	.V2C_6 (V2C_245_244),
	.V2C_7 (V2C_469_244),
	.V2C_8 (V2C_509_244),
	.V2C_9 (V2C_545_244),
	.V2C_10 (V2C_607_244),
	.V2C_11 (V2C_632_244),
	.V2C_12 (V2C_678_244),
	.V2C_13 (V2C_895_244),
	.V2C_14 (V2C_919_244),
	.V2C_15 (V2C_1003_244),
	.V2C_16 (V2C_1033_244),
	.V2C_17 (V2C_1060_244),
	.V2C_18 (V2C_1124_244),
	.V2C_19 (V2C_1395_244),
	.V2C_20 (V2C_1396_244),
	.C2V_1 (C2V_244_20),
	.C2V_2 (C2V_244_79),
	.C2V_3 (C2V_244_118),
	.C2V_4 (C2V_244_174),
	.C2V_5 (C2V_244_239),
	.C2V_6 (C2V_244_245),
	.C2V_7 (C2V_244_469),
	.C2V_8 (C2V_244_509),
	.C2V_9 (C2V_244_545),
	.C2V_10 (C2V_244_607),
	.C2V_11 (C2V_244_632),
	.C2V_12 (C2V_244_678),
	.C2V_13 (C2V_244_895),
	.C2V_14 (C2V_244_919),
	.C2V_15 (C2V_244_1003),
	.C2V_16 (C2V_244_1033),
	.C2V_17 (C2V_244_1060),
	.C2V_18 (C2V_244_1124),
	.C2V_19 (C2V_244_1395),
	.C2V_20 (C2V_244_1396),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU245 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_39_245),
	.V2C_2 (V2C_49_245),
	.V2C_3 (V2C_132_245),
	.V2C_4 (V2C_155_245),
	.V2C_5 (V2C_219_245),
	.V2C_6 (V2C_285_245),
	.V2C_7 (V2C_334_245),
	.V2C_8 (V2C_353_245),
	.V2C_9 (V2C_480_245),
	.V2C_10 (V2C_714_245),
	.V2C_11 (V2C_730_245),
	.V2C_12 (V2C_784_245),
	.V2C_13 (V2C_910_245),
	.V2C_14 (V2C_958_245),
	.V2C_15 (V2C_1001_245),
	.V2C_16 (V2C_1053_245),
	.V2C_17 (V2C_1102_245),
	.V2C_18 (V2C_1150_245),
	.V2C_19 (V2C_1396_245),
	.V2C_20 (V2C_1397_245),
	.C2V_1 (C2V_245_39),
	.C2V_2 (C2V_245_49),
	.C2V_3 (C2V_245_132),
	.C2V_4 (C2V_245_155),
	.C2V_5 (C2V_245_219),
	.C2V_6 (C2V_245_285),
	.C2V_7 (C2V_245_334),
	.C2V_8 (C2V_245_353),
	.C2V_9 (C2V_245_480),
	.C2V_10 (C2V_245_714),
	.C2V_11 (C2V_245_730),
	.C2V_12 (C2V_245_784),
	.C2V_13 (C2V_245_910),
	.C2V_14 (C2V_245_958),
	.C2V_15 (C2V_245_1001),
	.C2V_16 (C2V_245_1053),
	.C2V_17 (C2V_245_1102),
	.C2V_18 (C2V_245_1150),
	.C2V_19 (C2V_245_1396),
	.C2V_20 (C2V_245_1397),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU246 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_22_246),
	.V2C_2 (V2C_94_246),
	.V2C_3 (V2C_134_246),
	.V2C_4 (V2C_154_246),
	.V2C_5 (V2C_236_246),
	.V2C_6 (V2C_267_246),
	.V2C_7 (V2C_320_246),
	.V2C_8 (V2C_472_246),
	.V2C_9 (V2C_569_246),
	.V2C_10 (V2C_602_246),
	.V2C_11 (V2C_806_246),
	.V2C_12 (V2C_834_246),
	.V2C_13 (V2C_867_246),
	.V2C_14 (V2C_929_246),
	.V2C_15 (V2C_964_246),
	.V2C_16 (V2C_1031_246),
	.V2C_17 (V2C_1095_246),
	.V2C_18 (V2C_1145_246),
	.V2C_19 (V2C_1397_246),
	.V2C_20 (V2C_1398_246),
	.C2V_1 (C2V_246_22),
	.C2V_2 (C2V_246_94),
	.C2V_3 (C2V_246_134),
	.C2V_4 (C2V_246_154),
	.C2V_5 (C2V_246_236),
	.C2V_6 (C2V_246_267),
	.C2V_7 (C2V_246_320),
	.C2V_8 (C2V_246_472),
	.C2V_9 (C2V_246_569),
	.C2V_10 (C2V_246_602),
	.C2V_11 (C2V_246_806),
	.C2V_12 (C2V_246_834),
	.C2V_13 (C2V_246_867),
	.C2V_14 (C2V_246_929),
	.C2V_15 (C2V_246_964),
	.C2V_16 (C2V_246_1031),
	.C2V_17 (C2V_246_1095),
	.C2V_18 (C2V_246_1145),
	.C2V_19 (C2V_246_1397),
	.C2V_20 (C2V_246_1398),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU247 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_46_247),
	.V2C_2 (V2C_82_247),
	.V2C_3 (V2C_102_247),
	.V2C_4 (V2C_163_247),
	.V2C_5 (V2C_225_247),
	.V2C_6 (V2C_268_247),
	.V2C_7 (V2C_368_247),
	.V2C_8 (V2C_422_247),
	.V2C_9 (V2C_519_247),
	.V2C_10 (V2C_755_247),
	.V2C_11 (V2C_803_247),
	.V2C_12 (V2C_851_247),
	.V2C_13 (V2C_892_247),
	.V2C_14 (V2C_933_247),
	.V2C_15 (V2C_967_247),
	.V2C_16 (V2C_1054_247),
	.V2C_17 (V2C_1080_247),
	.V2C_18 (V2C_1139_247),
	.V2C_19 (V2C_1398_247),
	.V2C_20 (V2C_1399_247),
	.C2V_1 (C2V_247_46),
	.C2V_2 (C2V_247_82),
	.C2V_3 (C2V_247_102),
	.C2V_4 (C2V_247_163),
	.C2V_5 (C2V_247_225),
	.C2V_6 (C2V_247_268),
	.C2V_7 (C2V_247_368),
	.C2V_8 (C2V_247_422),
	.C2V_9 (C2V_247_519),
	.C2V_10 (C2V_247_755),
	.C2V_11 (C2V_247_803),
	.C2V_12 (C2V_247_851),
	.C2V_13 (C2V_247_892),
	.C2V_14 (C2V_247_933),
	.C2V_15 (C2V_247_967),
	.C2V_16 (C2V_247_1054),
	.C2V_17 (C2V_247_1080),
	.C2V_18 (C2V_247_1139),
	.C2V_19 (C2V_247_1398),
	.C2V_20 (C2V_247_1399),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU248 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_7_248),
	.V2C_2 (V2C_56_248),
	.V2C_3 (V2C_112_248),
	.V2C_4 (V2C_160_248),
	.V2C_5 (V2C_237_248),
	.V2C_6 (V2C_258_248),
	.V2C_7 (V2C_309_248),
	.V2C_8 (V2C_416_248),
	.V2C_9 (V2C_505_248),
	.V2C_10 (V2C_665_248),
	.V2C_11 (V2C_678_248),
	.V2C_12 (V2C_846_248),
	.V2C_13 (V2C_888_248),
	.V2C_14 (V2C_951_248),
	.V2C_15 (V2C_982_248),
	.V2C_16 (V2C_1014_248),
	.V2C_17 (V2C_1081_248),
	.V2C_18 (V2C_1112_248),
	.V2C_19 (V2C_1399_248),
	.V2C_20 (V2C_1400_248),
	.C2V_1 (C2V_248_7),
	.C2V_2 (C2V_248_56),
	.C2V_3 (C2V_248_112),
	.C2V_4 (C2V_248_160),
	.C2V_5 (C2V_248_237),
	.C2V_6 (C2V_248_258),
	.C2V_7 (C2V_248_309),
	.C2V_8 (C2V_248_416),
	.C2V_9 (C2V_248_505),
	.C2V_10 (C2V_248_665),
	.C2V_11 (C2V_248_678),
	.C2V_12 (C2V_248_846),
	.C2V_13 (C2V_248_888),
	.C2V_14 (C2V_248_951),
	.C2V_15 (C2V_248_982),
	.C2V_16 (C2V_248_1014),
	.C2V_17 (C2V_248_1081),
	.C2V_18 (C2V_248_1112),
	.C2V_19 (C2V_248_1399),
	.C2V_20 (C2V_248_1400),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU249 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_2_249),
	.V2C_2 (V2C_77_249),
	.V2C_3 (V2C_142_249),
	.V2C_4 (V2C_176_249),
	.V2C_5 (V2C_194_249),
	.V2C_6 (V2C_261_249),
	.V2C_7 (V2C_358_249),
	.V2C_8 (V2C_413_249),
	.V2C_9 (V2C_572_249),
	.V2C_10 (V2C_581_249),
	.V2C_11 (V2C_657_249),
	.V2C_12 (V2C_761_249),
	.V2C_13 (V2C_892_249),
	.V2C_14 (V2C_936_249),
	.V2C_15 (V2C_961_249),
	.V2C_16 (V2C_1021_249),
	.V2C_17 (V2C_1099_249),
	.V2C_18 (V2C_1144_249),
	.V2C_19 (V2C_1400_249),
	.V2C_20 (V2C_1401_249),
	.C2V_1 (C2V_249_2),
	.C2V_2 (C2V_249_77),
	.C2V_3 (C2V_249_142),
	.C2V_4 (C2V_249_176),
	.C2V_5 (C2V_249_194),
	.C2V_6 (C2V_249_261),
	.C2V_7 (C2V_249_358),
	.C2V_8 (C2V_249_413),
	.C2V_9 (C2V_249_572),
	.C2V_10 (C2V_249_581),
	.C2V_11 (C2V_249_657),
	.C2V_12 (C2V_249_761),
	.C2V_13 (C2V_249_892),
	.C2V_14 (C2V_249_936),
	.C2V_15 (C2V_249_961),
	.C2V_16 (C2V_249_1021),
	.C2V_17 (C2V_249_1099),
	.C2V_18 (C2V_249_1144),
	.C2V_19 (C2V_249_1400),
	.C2V_20 (C2V_249_1401),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU250 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_21_250),
	.V2C_2 (V2C_80_250),
	.V2C_3 (V2C_119_250),
	.V2C_4 (V2C_175_250),
	.V2C_5 (V2C_240_250),
	.V2C_6 (V2C_246_250),
	.V2C_7 (V2C_470_250),
	.V2C_8 (V2C_510_250),
	.V2C_9 (V2C_546_250),
	.V2C_10 (V2C_608_250),
	.V2C_11 (V2C_633_250),
	.V2C_12 (V2C_679_250),
	.V2C_13 (V2C_896_250),
	.V2C_14 (V2C_920_250),
	.V2C_15 (V2C_1004_250),
	.V2C_16 (V2C_1034_250),
	.V2C_17 (V2C_1061_250),
	.V2C_18 (V2C_1125_250),
	.V2C_19 (V2C_1401_250),
	.V2C_20 (V2C_1402_250),
	.C2V_1 (C2V_250_21),
	.C2V_2 (C2V_250_80),
	.C2V_3 (C2V_250_119),
	.C2V_4 (C2V_250_175),
	.C2V_5 (C2V_250_240),
	.C2V_6 (C2V_250_246),
	.C2V_7 (C2V_250_470),
	.C2V_8 (C2V_250_510),
	.C2V_9 (C2V_250_546),
	.C2V_10 (C2V_250_608),
	.C2V_11 (C2V_250_633),
	.C2V_12 (C2V_250_679),
	.C2V_13 (C2V_250_896),
	.C2V_14 (C2V_250_920),
	.C2V_15 (C2V_250_1004),
	.C2V_16 (C2V_250_1034),
	.C2V_17 (C2V_250_1061),
	.C2V_18 (C2V_250_1125),
	.C2V_19 (C2V_250_1401),
	.C2V_20 (C2V_250_1402),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU251 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_40_251),
	.V2C_2 (V2C_50_251),
	.V2C_3 (V2C_133_251),
	.V2C_4 (V2C_156_251),
	.V2C_5 (V2C_220_251),
	.V2C_6 (V2C_286_251),
	.V2C_7 (V2C_335_251),
	.V2C_8 (V2C_354_251),
	.V2C_9 (V2C_433_251),
	.V2C_10 (V2C_715_251),
	.V2C_11 (V2C_731_251),
	.V2C_12 (V2C_785_251),
	.V2C_13 (V2C_911_251),
	.V2C_14 (V2C_959_251),
	.V2C_15 (V2C_1002_251),
	.V2C_16 (V2C_1054_251),
	.V2C_17 (V2C_1103_251),
	.V2C_18 (V2C_1151_251),
	.V2C_19 (V2C_1402_251),
	.V2C_20 (V2C_1403_251),
	.C2V_1 (C2V_251_40),
	.C2V_2 (C2V_251_50),
	.C2V_3 (C2V_251_133),
	.C2V_4 (C2V_251_156),
	.C2V_5 (C2V_251_220),
	.C2V_6 (C2V_251_286),
	.C2V_7 (C2V_251_335),
	.C2V_8 (C2V_251_354),
	.C2V_9 (C2V_251_433),
	.C2V_10 (C2V_251_715),
	.C2V_11 (C2V_251_731),
	.C2V_12 (C2V_251_785),
	.C2V_13 (C2V_251_911),
	.C2V_14 (C2V_251_959),
	.C2V_15 (C2V_251_1002),
	.C2V_16 (C2V_251_1054),
	.C2V_17 (C2V_251_1103),
	.C2V_18 (C2V_251_1151),
	.C2V_19 (C2V_251_1402),
	.C2V_20 (C2V_251_1403),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU252 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_23_252),
	.V2C_2 (V2C_95_252),
	.V2C_3 (V2C_135_252),
	.V2C_4 (V2C_155_252),
	.V2C_5 (V2C_237_252),
	.V2C_6 (V2C_268_252),
	.V2C_7 (V2C_321_252),
	.V2C_8 (V2C_473_252),
	.V2C_9 (V2C_570_252),
	.V2C_10 (V2C_603_252),
	.V2C_11 (V2C_807_252),
	.V2C_12 (V2C_835_252),
	.V2C_13 (V2C_868_252),
	.V2C_14 (V2C_930_252),
	.V2C_15 (V2C_965_252),
	.V2C_16 (V2C_1032_252),
	.V2C_17 (V2C_1096_252),
	.V2C_18 (V2C_1146_252),
	.V2C_19 (V2C_1403_252),
	.V2C_20 (V2C_1404_252),
	.C2V_1 (C2V_252_23),
	.C2V_2 (C2V_252_95),
	.C2V_3 (C2V_252_135),
	.C2V_4 (C2V_252_155),
	.C2V_5 (C2V_252_237),
	.C2V_6 (C2V_252_268),
	.C2V_7 (C2V_252_321),
	.C2V_8 (C2V_252_473),
	.C2V_9 (C2V_252_570),
	.C2V_10 (C2V_252_603),
	.C2V_11 (C2V_252_807),
	.C2V_12 (C2V_252_835),
	.C2V_13 (C2V_252_868),
	.C2V_14 (C2V_252_930),
	.C2V_15 (C2V_252_965),
	.C2V_16 (C2V_252_1032),
	.C2V_17 (C2V_252_1096),
	.C2V_18 (C2V_252_1146),
	.C2V_19 (C2V_252_1403),
	.C2V_20 (C2V_252_1404),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU253 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_47_253),
	.V2C_2 (V2C_83_253),
	.V2C_3 (V2C_103_253),
	.V2C_4 (V2C_164_253),
	.V2C_5 (V2C_226_253),
	.V2C_6 (V2C_269_253),
	.V2C_7 (V2C_369_253),
	.V2C_8 (V2C_423_253),
	.V2C_9 (V2C_520_253),
	.V2C_10 (V2C_756_253),
	.V2C_11 (V2C_804_253),
	.V2C_12 (V2C_852_253),
	.V2C_13 (V2C_893_253),
	.V2C_14 (V2C_934_253),
	.V2C_15 (V2C_968_253),
	.V2C_16 (V2C_1055_253),
	.V2C_17 (V2C_1081_253),
	.V2C_18 (V2C_1140_253),
	.V2C_19 (V2C_1404_253),
	.V2C_20 (V2C_1405_253),
	.C2V_1 (C2V_253_47),
	.C2V_2 (C2V_253_83),
	.C2V_3 (C2V_253_103),
	.C2V_4 (C2V_253_164),
	.C2V_5 (C2V_253_226),
	.C2V_6 (C2V_253_269),
	.C2V_7 (C2V_253_369),
	.C2V_8 (C2V_253_423),
	.C2V_9 (C2V_253_520),
	.C2V_10 (C2V_253_756),
	.C2V_11 (C2V_253_804),
	.C2V_12 (C2V_253_852),
	.C2V_13 (C2V_253_893),
	.C2V_14 (C2V_253_934),
	.C2V_15 (C2V_253_968),
	.C2V_16 (C2V_253_1055),
	.C2V_17 (C2V_253_1081),
	.C2V_18 (C2V_253_1140),
	.C2V_19 (C2V_253_1404),
	.C2V_20 (C2V_253_1405),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU254 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_8_254),
	.V2C_2 (V2C_57_254),
	.V2C_3 (V2C_113_254),
	.V2C_4 (V2C_161_254),
	.V2C_5 (V2C_238_254),
	.V2C_6 (V2C_259_254),
	.V2C_7 (V2C_310_254),
	.V2C_8 (V2C_417_254),
	.V2C_9 (V2C_506_254),
	.V2C_10 (V2C_666_254),
	.V2C_11 (V2C_679_254),
	.V2C_12 (V2C_847_254),
	.V2C_13 (V2C_889_254),
	.V2C_14 (V2C_952_254),
	.V2C_15 (V2C_983_254),
	.V2C_16 (V2C_1015_254),
	.V2C_17 (V2C_1082_254),
	.V2C_18 (V2C_1113_254),
	.V2C_19 (V2C_1405_254),
	.V2C_20 (V2C_1406_254),
	.C2V_1 (C2V_254_8),
	.C2V_2 (C2V_254_57),
	.C2V_3 (C2V_254_113),
	.C2V_4 (C2V_254_161),
	.C2V_5 (C2V_254_238),
	.C2V_6 (C2V_254_259),
	.C2V_7 (C2V_254_310),
	.C2V_8 (C2V_254_417),
	.C2V_9 (C2V_254_506),
	.C2V_10 (C2V_254_666),
	.C2V_11 (C2V_254_679),
	.C2V_12 (C2V_254_847),
	.C2V_13 (C2V_254_889),
	.C2V_14 (C2V_254_952),
	.C2V_15 (C2V_254_983),
	.C2V_16 (C2V_254_1015),
	.C2V_17 (C2V_254_1082),
	.C2V_18 (C2V_254_1113),
	.C2V_19 (C2V_254_1405),
	.C2V_20 (C2V_254_1406),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU255 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_3_255),
	.V2C_2 (V2C_78_255),
	.V2C_3 (V2C_143_255),
	.V2C_4 (V2C_177_255),
	.V2C_5 (V2C_195_255),
	.V2C_6 (V2C_262_255),
	.V2C_7 (V2C_359_255),
	.V2C_8 (V2C_414_255),
	.V2C_9 (V2C_573_255),
	.V2C_10 (V2C_582_255),
	.V2C_11 (V2C_658_255),
	.V2C_12 (V2C_762_255),
	.V2C_13 (V2C_893_255),
	.V2C_14 (V2C_937_255),
	.V2C_15 (V2C_962_255),
	.V2C_16 (V2C_1022_255),
	.V2C_17 (V2C_1100_255),
	.V2C_18 (V2C_1145_255),
	.V2C_19 (V2C_1406_255),
	.V2C_20 (V2C_1407_255),
	.C2V_1 (C2V_255_3),
	.C2V_2 (C2V_255_78),
	.C2V_3 (C2V_255_143),
	.C2V_4 (C2V_255_177),
	.C2V_5 (C2V_255_195),
	.C2V_6 (C2V_255_262),
	.C2V_7 (C2V_255_359),
	.C2V_8 (C2V_255_414),
	.C2V_9 (C2V_255_573),
	.C2V_10 (C2V_255_582),
	.C2V_11 (C2V_255_658),
	.C2V_12 (C2V_255_762),
	.C2V_13 (C2V_255_893),
	.C2V_14 (C2V_255_937),
	.C2V_15 (C2V_255_962),
	.C2V_16 (C2V_255_1022),
	.C2V_17 (C2V_255_1100),
	.C2V_18 (C2V_255_1145),
	.C2V_19 (C2V_255_1406),
	.C2V_20 (C2V_255_1407),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU256 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_22_256),
	.V2C_2 (V2C_81_256),
	.V2C_3 (V2C_120_256),
	.V2C_4 (V2C_176_256),
	.V2C_5 (V2C_193_256),
	.V2C_6 (V2C_247_256),
	.V2C_7 (V2C_471_256),
	.V2C_8 (V2C_511_256),
	.V2C_9 (V2C_547_256),
	.V2C_10 (V2C_609_256),
	.V2C_11 (V2C_634_256),
	.V2C_12 (V2C_680_256),
	.V2C_13 (V2C_897_256),
	.V2C_14 (V2C_921_256),
	.V2C_15 (V2C_1005_256),
	.V2C_16 (V2C_1035_256),
	.V2C_17 (V2C_1062_256),
	.V2C_18 (V2C_1126_256),
	.V2C_19 (V2C_1407_256),
	.V2C_20 (V2C_1408_256),
	.C2V_1 (C2V_256_22),
	.C2V_2 (C2V_256_81),
	.C2V_3 (C2V_256_120),
	.C2V_4 (C2V_256_176),
	.C2V_5 (C2V_256_193),
	.C2V_6 (C2V_256_247),
	.C2V_7 (C2V_256_471),
	.C2V_8 (C2V_256_511),
	.C2V_9 (C2V_256_547),
	.C2V_10 (C2V_256_609),
	.C2V_11 (C2V_256_634),
	.C2V_12 (C2V_256_680),
	.C2V_13 (C2V_256_897),
	.C2V_14 (C2V_256_921),
	.C2V_15 (C2V_256_1005),
	.C2V_16 (C2V_256_1035),
	.C2V_17 (C2V_256_1062),
	.C2V_18 (C2V_256_1126),
	.C2V_19 (C2V_256_1407),
	.C2V_20 (C2V_256_1408),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU257 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_41_257),
	.V2C_2 (V2C_51_257),
	.V2C_3 (V2C_134_257),
	.V2C_4 (V2C_157_257),
	.V2C_5 (V2C_221_257),
	.V2C_6 (V2C_287_257),
	.V2C_7 (V2C_336_257),
	.V2C_8 (V2C_355_257),
	.V2C_9 (V2C_434_257),
	.V2C_10 (V2C_716_257),
	.V2C_11 (V2C_732_257),
	.V2C_12 (V2C_786_257),
	.V2C_13 (V2C_912_257),
	.V2C_14 (V2C_960_257),
	.V2C_15 (V2C_1003_257),
	.V2C_16 (V2C_1055_257),
	.V2C_17 (V2C_1104_257),
	.V2C_18 (V2C_1152_257),
	.V2C_19 (V2C_1408_257),
	.V2C_20 (V2C_1409_257),
	.C2V_1 (C2V_257_41),
	.C2V_2 (C2V_257_51),
	.C2V_3 (C2V_257_134),
	.C2V_4 (C2V_257_157),
	.C2V_5 (C2V_257_221),
	.C2V_6 (C2V_257_287),
	.C2V_7 (C2V_257_336),
	.C2V_8 (C2V_257_355),
	.C2V_9 (C2V_257_434),
	.C2V_10 (C2V_257_716),
	.C2V_11 (C2V_257_732),
	.C2V_12 (C2V_257_786),
	.C2V_13 (C2V_257_912),
	.C2V_14 (C2V_257_960),
	.C2V_15 (C2V_257_1003),
	.C2V_16 (C2V_257_1055),
	.C2V_17 (C2V_257_1104),
	.C2V_18 (C2V_257_1152),
	.C2V_19 (C2V_257_1408),
	.C2V_20 (C2V_257_1409),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU258 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_24_258),
	.V2C_2 (V2C_96_258),
	.V2C_3 (V2C_136_258),
	.V2C_4 (V2C_156_258),
	.V2C_5 (V2C_238_258),
	.V2C_6 (V2C_269_258),
	.V2C_7 (V2C_322_258),
	.V2C_8 (V2C_474_258),
	.V2C_9 (V2C_571_258),
	.V2C_10 (V2C_604_258),
	.V2C_11 (V2C_808_258),
	.V2C_12 (V2C_836_258),
	.V2C_13 (V2C_869_258),
	.V2C_14 (V2C_931_258),
	.V2C_15 (V2C_966_258),
	.V2C_16 (V2C_1033_258),
	.V2C_17 (V2C_1097_258),
	.V2C_18 (V2C_1147_258),
	.V2C_19 (V2C_1409_258),
	.V2C_20 (V2C_1410_258),
	.C2V_1 (C2V_258_24),
	.C2V_2 (C2V_258_96),
	.C2V_3 (C2V_258_136),
	.C2V_4 (C2V_258_156),
	.C2V_5 (C2V_258_238),
	.C2V_6 (C2V_258_269),
	.C2V_7 (C2V_258_322),
	.C2V_8 (C2V_258_474),
	.C2V_9 (C2V_258_571),
	.C2V_10 (C2V_258_604),
	.C2V_11 (C2V_258_808),
	.C2V_12 (C2V_258_836),
	.C2V_13 (C2V_258_869),
	.C2V_14 (C2V_258_931),
	.C2V_15 (C2V_258_966),
	.C2V_16 (C2V_258_1033),
	.C2V_17 (C2V_258_1097),
	.C2V_18 (C2V_258_1147),
	.C2V_19 (C2V_258_1409),
	.C2V_20 (C2V_258_1410),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU259 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_48_259),
	.V2C_2 (V2C_84_259),
	.V2C_3 (V2C_104_259),
	.V2C_4 (V2C_165_259),
	.V2C_5 (V2C_227_259),
	.V2C_6 (V2C_270_259),
	.V2C_7 (V2C_370_259),
	.V2C_8 (V2C_424_259),
	.V2C_9 (V2C_521_259),
	.V2C_10 (V2C_757_259),
	.V2C_11 (V2C_805_259),
	.V2C_12 (V2C_853_259),
	.V2C_13 (V2C_894_259),
	.V2C_14 (V2C_935_259),
	.V2C_15 (V2C_969_259),
	.V2C_16 (V2C_1056_259),
	.V2C_17 (V2C_1082_259),
	.V2C_18 (V2C_1141_259),
	.V2C_19 (V2C_1410_259),
	.V2C_20 (V2C_1411_259),
	.C2V_1 (C2V_259_48),
	.C2V_2 (C2V_259_84),
	.C2V_3 (C2V_259_104),
	.C2V_4 (C2V_259_165),
	.C2V_5 (C2V_259_227),
	.C2V_6 (C2V_259_270),
	.C2V_7 (C2V_259_370),
	.C2V_8 (C2V_259_424),
	.C2V_9 (C2V_259_521),
	.C2V_10 (C2V_259_757),
	.C2V_11 (C2V_259_805),
	.C2V_12 (C2V_259_853),
	.C2V_13 (C2V_259_894),
	.C2V_14 (C2V_259_935),
	.C2V_15 (C2V_259_969),
	.C2V_16 (C2V_259_1056),
	.C2V_17 (C2V_259_1082),
	.C2V_18 (C2V_259_1141),
	.C2V_19 (C2V_259_1410),
	.C2V_20 (C2V_259_1411),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU260 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_9_260),
	.V2C_2 (V2C_58_260),
	.V2C_3 (V2C_114_260),
	.V2C_4 (V2C_162_260),
	.V2C_5 (V2C_239_260),
	.V2C_6 (V2C_260_260),
	.V2C_7 (V2C_311_260),
	.V2C_8 (V2C_418_260),
	.V2C_9 (V2C_507_260),
	.V2C_10 (V2C_667_260),
	.V2C_11 (V2C_680_260),
	.V2C_12 (V2C_848_260),
	.V2C_13 (V2C_890_260),
	.V2C_14 (V2C_953_260),
	.V2C_15 (V2C_984_260),
	.V2C_16 (V2C_1016_260),
	.V2C_17 (V2C_1083_260),
	.V2C_18 (V2C_1114_260),
	.V2C_19 (V2C_1411_260),
	.V2C_20 (V2C_1412_260),
	.C2V_1 (C2V_260_9),
	.C2V_2 (C2V_260_58),
	.C2V_3 (C2V_260_114),
	.C2V_4 (C2V_260_162),
	.C2V_5 (C2V_260_239),
	.C2V_6 (C2V_260_260),
	.C2V_7 (C2V_260_311),
	.C2V_8 (C2V_260_418),
	.C2V_9 (C2V_260_507),
	.C2V_10 (C2V_260_667),
	.C2V_11 (C2V_260_680),
	.C2V_12 (C2V_260_848),
	.C2V_13 (C2V_260_890),
	.C2V_14 (C2V_260_953),
	.C2V_15 (C2V_260_984),
	.C2V_16 (C2V_260_1016),
	.C2V_17 (C2V_260_1083),
	.C2V_18 (C2V_260_1114),
	.C2V_19 (C2V_260_1411),
	.C2V_20 (C2V_260_1412),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU261 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_4_261),
	.V2C_2 (V2C_79_261),
	.V2C_3 (V2C_144_261),
	.V2C_4 (V2C_178_261),
	.V2C_5 (V2C_196_261),
	.V2C_6 (V2C_263_261),
	.V2C_7 (V2C_360_261),
	.V2C_8 (V2C_415_261),
	.V2C_9 (V2C_574_261),
	.V2C_10 (V2C_583_261),
	.V2C_11 (V2C_659_261),
	.V2C_12 (V2C_763_261),
	.V2C_13 (V2C_894_261),
	.V2C_14 (V2C_938_261),
	.V2C_15 (V2C_963_261),
	.V2C_16 (V2C_1023_261),
	.V2C_17 (V2C_1101_261),
	.V2C_18 (V2C_1146_261),
	.V2C_19 (V2C_1412_261),
	.V2C_20 (V2C_1413_261),
	.C2V_1 (C2V_261_4),
	.C2V_2 (C2V_261_79),
	.C2V_3 (C2V_261_144),
	.C2V_4 (C2V_261_178),
	.C2V_5 (C2V_261_196),
	.C2V_6 (C2V_261_263),
	.C2V_7 (C2V_261_360),
	.C2V_8 (C2V_261_415),
	.C2V_9 (C2V_261_574),
	.C2V_10 (C2V_261_583),
	.C2V_11 (C2V_261_659),
	.C2V_12 (C2V_261_763),
	.C2V_13 (C2V_261_894),
	.C2V_14 (C2V_261_938),
	.C2V_15 (C2V_261_963),
	.C2V_16 (C2V_261_1023),
	.C2V_17 (C2V_261_1101),
	.C2V_18 (C2V_261_1146),
	.C2V_19 (C2V_261_1412),
	.C2V_20 (C2V_261_1413),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU262 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_23_262),
	.V2C_2 (V2C_82_262),
	.V2C_3 (V2C_121_262),
	.V2C_4 (V2C_177_262),
	.V2C_5 (V2C_194_262),
	.V2C_6 (V2C_248_262),
	.V2C_7 (V2C_472_262),
	.V2C_8 (V2C_512_262),
	.V2C_9 (V2C_548_262),
	.V2C_10 (V2C_610_262),
	.V2C_11 (V2C_635_262),
	.V2C_12 (V2C_681_262),
	.V2C_13 (V2C_898_262),
	.V2C_14 (V2C_922_262),
	.V2C_15 (V2C_1006_262),
	.V2C_16 (V2C_1036_262),
	.V2C_17 (V2C_1063_262),
	.V2C_18 (V2C_1127_262),
	.V2C_19 (V2C_1413_262),
	.V2C_20 (V2C_1414_262),
	.C2V_1 (C2V_262_23),
	.C2V_2 (C2V_262_82),
	.C2V_3 (C2V_262_121),
	.C2V_4 (C2V_262_177),
	.C2V_5 (C2V_262_194),
	.C2V_6 (C2V_262_248),
	.C2V_7 (C2V_262_472),
	.C2V_8 (C2V_262_512),
	.C2V_9 (C2V_262_548),
	.C2V_10 (C2V_262_610),
	.C2V_11 (C2V_262_635),
	.C2V_12 (C2V_262_681),
	.C2V_13 (C2V_262_898),
	.C2V_14 (C2V_262_922),
	.C2V_15 (C2V_262_1006),
	.C2V_16 (C2V_262_1036),
	.C2V_17 (C2V_262_1063),
	.C2V_18 (C2V_262_1127),
	.C2V_19 (C2V_262_1413),
	.C2V_20 (C2V_262_1414),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU263 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_42_263),
	.V2C_2 (V2C_52_263),
	.V2C_3 (V2C_135_263),
	.V2C_4 (V2C_158_263),
	.V2C_5 (V2C_222_263),
	.V2C_6 (V2C_288_263),
	.V2C_7 (V2C_289_263),
	.V2C_8 (V2C_356_263),
	.V2C_9 (V2C_435_263),
	.V2C_10 (V2C_717_263),
	.V2C_11 (V2C_733_263),
	.V2C_12 (V2C_787_263),
	.V2C_13 (V2C_865_263),
	.V2C_14 (V2C_913_263),
	.V2C_15 (V2C_1004_263),
	.V2C_16 (V2C_1056_263),
	.V2C_17 (V2C_1057_263),
	.V2C_18 (V2C_1105_263),
	.V2C_19 (V2C_1414_263),
	.V2C_20 (V2C_1415_263),
	.C2V_1 (C2V_263_42),
	.C2V_2 (C2V_263_52),
	.C2V_3 (C2V_263_135),
	.C2V_4 (C2V_263_158),
	.C2V_5 (C2V_263_222),
	.C2V_6 (C2V_263_288),
	.C2V_7 (C2V_263_289),
	.C2V_8 (C2V_263_356),
	.C2V_9 (C2V_263_435),
	.C2V_10 (C2V_263_717),
	.C2V_11 (C2V_263_733),
	.C2V_12 (C2V_263_787),
	.C2V_13 (C2V_263_865),
	.C2V_14 (C2V_263_913),
	.C2V_15 (C2V_263_1004),
	.C2V_16 (C2V_263_1056),
	.C2V_17 (C2V_263_1057),
	.C2V_18 (C2V_263_1105),
	.C2V_19 (C2V_263_1414),
	.C2V_20 (C2V_263_1415),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU264 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_25_264),
	.V2C_2 (V2C_49_264),
	.V2C_3 (V2C_137_264),
	.V2C_4 (V2C_157_264),
	.V2C_5 (V2C_239_264),
	.V2C_6 (V2C_270_264),
	.V2C_7 (V2C_323_264),
	.V2C_8 (V2C_475_264),
	.V2C_9 (V2C_572_264),
	.V2C_10 (V2C_605_264),
	.V2C_11 (V2C_809_264),
	.V2C_12 (V2C_837_264),
	.V2C_13 (V2C_870_264),
	.V2C_14 (V2C_932_264),
	.V2C_15 (V2C_967_264),
	.V2C_16 (V2C_1034_264),
	.V2C_17 (V2C_1098_264),
	.V2C_18 (V2C_1148_264),
	.V2C_19 (V2C_1415_264),
	.V2C_20 (V2C_1416_264),
	.C2V_1 (C2V_264_25),
	.C2V_2 (C2V_264_49),
	.C2V_3 (C2V_264_137),
	.C2V_4 (C2V_264_157),
	.C2V_5 (C2V_264_239),
	.C2V_6 (C2V_264_270),
	.C2V_7 (C2V_264_323),
	.C2V_8 (C2V_264_475),
	.C2V_9 (C2V_264_572),
	.C2V_10 (C2V_264_605),
	.C2V_11 (C2V_264_809),
	.C2V_12 (C2V_264_837),
	.C2V_13 (C2V_264_870),
	.C2V_14 (C2V_264_932),
	.C2V_15 (C2V_264_967),
	.C2V_16 (C2V_264_1034),
	.C2V_17 (C2V_264_1098),
	.C2V_18 (C2V_264_1148),
	.C2V_19 (C2V_264_1415),
	.C2V_20 (C2V_264_1416),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU265 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_1_265),
	.V2C_2 (V2C_85_265),
	.V2C_3 (V2C_105_265),
	.V2C_4 (V2C_166_265),
	.V2C_5 (V2C_228_265),
	.V2C_6 (V2C_271_265),
	.V2C_7 (V2C_371_265),
	.V2C_8 (V2C_425_265),
	.V2C_9 (V2C_522_265),
	.V2C_10 (V2C_758_265),
	.V2C_11 (V2C_806_265),
	.V2C_12 (V2C_854_265),
	.V2C_13 (V2C_895_265),
	.V2C_14 (V2C_936_265),
	.V2C_15 (V2C_970_265),
	.V2C_16 (V2C_1009_265),
	.V2C_17 (V2C_1083_265),
	.V2C_18 (V2C_1142_265),
	.V2C_19 (V2C_1416_265),
	.V2C_20 (V2C_1417_265),
	.C2V_1 (C2V_265_1),
	.C2V_2 (C2V_265_85),
	.C2V_3 (C2V_265_105),
	.C2V_4 (C2V_265_166),
	.C2V_5 (C2V_265_228),
	.C2V_6 (C2V_265_271),
	.C2V_7 (C2V_265_371),
	.C2V_8 (C2V_265_425),
	.C2V_9 (C2V_265_522),
	.C2V_10 (C2V_265_758),
	.C2V_11 (C2V_265_806),
	.C2V_12 (C2V_265_854),
	.C2V_13 (C2V_265_895),
	.C2V_14 (C2V_265_936),
	.C2V_15 (C2V_265_970),
	.C2V_16 (C2V_265_1009),
	.C2V_17 (C2V_265_1083),
	.C2V_18 (C2V_265_1142),
	.C2V_19 (C2V_265_1416),
	.C2V_20 (C2V_265_1417),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU266 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_10_266),
	.V2C_2 (V2C_59_266),
	.V2C_3 (V2C_115_266),
	.V2C_4 (V2C_163_266),
	.V2C_5 (V2C_240_266),
	.V2C_6 (V2C_261_266),
	.V2C_7 (V2C_312_266),
	.V2C_8 (V2C_419_266),
	.V2C_9 (V2C_508_266),
	.V2C_10 (V2C_668_266),
	.V2C_11 (V2C_681_266),
	.V2C_12 (V2C_849_266),
	.V2C_13 (V2C_891_266),
	.V2C_14 (V2C_954_266),
	.V2C_15 (V2C_985_266),
	.V2C_16 (V2C_1017_266),
	.V2C_17 (V2C_1084_266),
	.V2C_18 (V2C_1115_266),
	.V2C_19 (V2C_1417_266),
	.V2C_20 (V2C_1418_266),
	.C2V_1 (C2V_266_10),
	.C2V_2 (C2V_266_59),
	.C2V_3 (C2V_266_115),
	.C2V_4 (C2V_266_163),
	.C2V_5 (C2V_266_240),
	.C2V_6 (C2V_266_261),
	.C2V_7 (C2V_266_312),
	.C2V_8 (C2V_266_419),
	.C2V_9 (C2V_266_508),
	.C2V_10 (C2V_266_668),
	.C2V_11 (C2V_266_681),
	.C2V_12 (C2V_266_849),
	.C2V_13 (C2V_266_891),
	.C2V_14 (C2V_266_954),
	.C2V_15 (C2V_266_985),
	.C2V_16 (C2V_266_1017),
	.C2V_17 (C2V_266_1084),
	.C2V_18 (C2V_266_1115),
	.C2V_19 (C2V_266_1417),
	.C2V_20 (C2V_266_1418),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU267 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_5_267),
	.V2C_2 (V2C_80_267),
	.V2C_3 (V2C_97_267),
	.V2C_4 (V2C_179_267),
	.V2C_5 (V2C_197_267),
	.V2C_6 (V2C_264_267),
	.V2C_7 (V2C_361_267),
	.V2C_8 (V2C_416_267),
	.V2C_9 (V2C_575_267),
	.V2C_10 (V2C_584_267),
	.V2C_11 (V2C_660_267),
	.V2C_12 (V2C_764_267),
	.V2C_13 (V2C_895_267),
	.V2C_14 (V2C_939_267),
	.V2C_15 (V2C_964_267),
	.V2C_16 (V2C_1024_267),
	.V2C_17 (V2C_1102_267),
	.V2C_18 (V2C_1147_267),
	.V2C_19 (V2C_1418_267),
	.V2C_20 (V2C_1419_267),
	.C2V_1 (C2V_267_5),
	.C2V_2 (C2V_267_80),
	.C2V_3 (C2V_267_97),
	.C2V_4 (C2V_267_179),
	.C2V_5 (C2V_267_197),
	.C2V_6 (C2V_267_264),
	.C2V_7 (C2V_267_361),
	.C2V_8 (C2V_267_416),
	.C2V_9 (C2V_267_575),
	.C2V_10 (C2V_267_584),
	.C2V_11 (C2V_267_660),
	.C2V_12 (C2V_267_764),
	.C2V_13 (C2V_267_895),
	.C2V_14 (C2V_267_939),
	.C2V_15 (C2V_267_964),
	.C2V_16 (C2V_267_1024),
	.C2V_17 (C2V_267_1102),
	.C2V_18 (C2V_267_1147),
	.C2V_19 (C2V_267_1418),
	.C2V_20 (C2V_267_1419),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU268 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_24_268),
	.V2C_2 (V2C_83_268),
	.V2C_3 (V2C_122_268),
	.V2C_4 (V2C_178_268),
	.V2C_5 (V2C_195_268),
	.V2C_6 (V2C_249_268),
	.V2C_7 (V2C_473_268),
	.V2C_8 (V2C_513_268),
	.V2C_9 (V2C_549_268),
	.V2C_10 (V2C_611_268),
	.V2C_11 (V2C_636_268),
	.V2C_12 (V2C_682_268),
	.V2C_13 (V2C_899_268),
	.V2C_14 (V2C_923_268),
	.V2C_15 (V2C_1007_268),
	.V2C_16 (V2C_1037_268),
	.V2C_17 (V2C_1064_268),
	.V2C_18 (V2C_1128_268),
	.V2C_19 (V2C_1419_268),
	.V2C_20 (V2C_1420_268),
	.C2V_1 (C2V_268_24),
	.C2V_2 (C2V_268_83),
	.C2V_3 (C2V_268_122),
	.C2V_4 (C2V_268_178),
	.C2V_5 (C2V_268_195),
	.C2V_6 (C2V_268_249),
	.C2V_7 (C2V_268_473),
	.C2V_8 (C2V_268_513),
	.C2V_9 (C2V_268_549),
	.C2V_10 (C2V_268_611),
	.C2V_11 (C2V_268_636),
	.C2V_12 (C2V_268_682),
	.C2V_13 (C2V_268_899),
	.C2V_14 (C2V_268_923),
	.C2V_15 (C2V_268_1007),
	.C2V_16 (C2V_268_1037),
	.C2V_17 (C2V_268_1064),
	.C2V_18 (C2V_268_1128),
	.C2V_19 (C2V_268_1419),
	.C2V_20 (C2V_268_1420),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU269 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_43_269),
	.V2C_2 (V2C_53_269),
	.V2C_3 (V2C_136_269),
	.V2C_4 (V2C_159_269),
	.V2C_5 (V2C_223_269),
	.V2C_6 (V2C_241_269),
	.V2C_7 (V2C_290_269),
	.V2C_8 (V2C_357_269),
	.V2C_9 (V2C_436_269),
	.V2C_10 (V2C_718_269),
	.V2C_11 (V2C_734_269),
	.V2C_12 (V2C_788_269),
	.V2C_13 (V2C_866_269),
	.V2C_14 (V2C_914_269),
	.V2C_15 (V2C_1005_269),
	.V2C_16 (V2C_1009_269),
	.V2C_17 (V2C_1058_269),
	.V2C_18 (V2C_1106_269),
	.V2C_19 (V2C_1420_269),
	.V2C_20 (V2C_1421_269),
	.C2V_1 (C2V_269_43),
	.C2V_2 (C2V_269_53),
	.C2V_3 (C2V_269_136),
	.C2V_4 (C2V_269_159),
	.C2V_5 (C2V_269_223),
	.C2V_6 (C2V_269_241),
	.C2V_7 (C2V_269_290),
	.C2V_8 (C2V_269_357),
	.C2V_9 (C2V_269_436),
	.C2V_10 (C2V_269_718),
	.C2V_11 (C2V_269_734),
	.C2V_12 (C2V_269_788),
	.C2V_13 (C2V_269_866),
	.C2V_14 (C2V_269_914),
	.C2V_15 (C2V_269_1005),
	.C2V_16 (C2V_269_1009),
	.C2V_17 (C2V_269_1058),
	.C2V_18 (C2V_269_1106),
	.C2V_19 (C2V_269_1420),
	.C2V_20 (C2V_269_1421),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU270 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_26_270),
	.V2C_2 (V2C_50_270),
	.V2C_3 (V2C_138_270),
	.V2C_4 (V2C_158_270),
	.V2C_5 (V2C_240_270),
	.V2C_6 (V2C_271_270),
	.V2C_7 (V2C_324_270),
	.V2C_8 (V2C_476_270),
	.V2C_9 (V2C_573_270),
	.V2C_10 (V2C_606_270),
	.V2C_11 (V2C_810_270),
	.V2C_12 (V2C_838_270),
	.V2C_13 (V2C_871_270),
	.V2C_14 (V2C_933_270),
	.V2C_15 (V2C_968_270),
	.V2C_16 (V2C_1035_270),
	.V2C_17 (V2C_1099_270),
	.V2C_18 (V2C_1149_270),
	.V2C_19 (V2C_1421_270),
	.V2C_20 (V2C_1422_270),
	.C2V_1 (C2V_270_26),
	.C2V_2 (C2V_270_50),
	.C2V_3 (C2V_270_138),
	.C2V_4 (C2V_270_158),
	.C2V_5 (C2V_270_240),
	.C2V_6 (C2V_270_271),
	.C2V_7 (C2V_270_324),
	.C2V_8 (C2V_270_476),
	.C2V_9 (C2V_270_573),
	.C2V_10 (C2V_270_606),
	.C2V_11 (C2V_270_810),
	.C2V_12 (C2V_270_838),
	.C2V_13 (C2V_270_871),
	.C2V_14 (C2V_270_933),
	.C2V_15 (C2V_270_968),
	.C2V_16 (C2V_270_1035),
	.C2V_17 (C2V_270_1099),
	.C2V_18 (C2V_270_1149),
	.C2V_19 (C2V_270_1421),
	.C2V_20 (C2V_270_1422),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU271 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_2_271),
	.V2C_2 (V2C_86_271),
	.V2C_3 (V2C_106_271),
	.V2C_4 (V2C_167_271),
	.V2C_5 (V2C_229_271),
	.V2C_6 (V2C_272_271),
	.V2C_7 (V2C_372_271),
	.V2C_8 (V2C_426_271),
	.V2C_9 (V2C_523_271),
	.V2C_10 (V2C_759_271),
	.V2C_11 (V2C_807_271),
	.V2C_12 (V2C_855_271),
	.V2C_13 (V2C_896_271),
	.V2C_14 (V2C_937_271),
	.V2C_15 (V2C_971_271),
	.V2C_16 (V2C_1010_271),
	.V2C_17 (V2C_1084_271),
	.V2C_18 (V2C_1143_271),
	.V2C_19 (V2C_1422_271),
	.V2C_20 (V2C_1423_271),
	.C2V_1 (C2V_271_2),
	.C2V_2 (C2V_271_86),
	.C2V_3 (C2V_271_106),
	.C2V_4 (C2V_271_167),
	.C2V_5 (C2V_271_229),
	.C2V_6 (C2V_271_272),
	.C2V_7 (C2V_271_372),
	.C2V_8 (C2V_271_426),
	.C2V_9 (C2V_271_523),
	.C2V_10 (C2V_271_759),
	.C2V_11 (C2V_271_807),
	.C2V_12 (C2V_271_855),
	.C2V_13 (C2V_271_896),
	.C2V_14 (C2V_271_937),
	.C2V_15 (C2V_271_971),
	.C2V_16 (C2V_271_1010),
	.C2V_17 (C2V_271_1084),
	.C2V_18 (C2V_271_1143),
	.C2V_19 (C2V_271_1422),
	.C2V_20 (C2V_271_1423),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU272 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_11_272),
	.V2C_2 (V2C_60_272),
	.V2C_3 (V2C_116_272),
	.V2C_4 (V2C_164_272),
	.V2C_5 (V2C_193_272),
	.V2C_6 (V2C_262_272),
	.V2C_7 (V2C_313_272),
	.V2C_8 (V2C_420_272),
	.V2C_9 (V2C_509_272),
	.V2C_10 (V2C_669_272),
	.V2C_11 (V2C_682_272),
	.V2C_12 (V2C_850_272),
	.V2C_13 (V2C_892_272),
	.V2C_14 (V2C_955_272),
	.V2C_15 (V2C_986_272),
	.V2C_16 (V2C_1018_272),
	.V2C_17 (V2C_1085_272),
	.V2C_18 (V2C_1116_272),
	.V2C_19 (V2C_1423_272),
	.V2C_20 (V2C_1424_272),
	.C2V_1 (C2V_272_11),
	.C2V_2 (C2V_272_60),
	.C2V_3 (C2V_272_116),
	.C2V_4 (C2V_272_164),
	.C2V_5 (C2V_272_193),
	.C2V_6 (C2V_272_262),
	.C2V_7 (C2V_272_313),
	.C2V_8 (C2V_272_420),
	.C2V_9 (C2V_272_509),
	.C2V_10 (C2V_272_669),
	.C2V_11 (C2V_272_682),
	.C2V_12 (C2V_272_850),
	.C2V_13 (C2V_272_892),
	.C2V_14 (C2V_272_955),
	.C2V_15 (C2V_272_986),
	.C2V_16 (C2V_272_1018),
	.C2V_17 (C2V_272_1085),
	.C2V_18 (C2V_272_1116),
	.C2V_19 (C2V_272_1423),
	.C2V_20 (C2V_272_1424),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU273 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_6_273),
	.V2C_2 (V2C_81_273),
	.V2C_3 (V2C_98_273),
	.V2C_4 (V2C_180_273),
	.V2C_5 (V2C_198_273),
	.V2C_6 (V2C_265_273),
	.V2C_7 (V2C_362_273),
	.V2C_8 (V2C_417_273),
	.V2C_9 (V2C_576_273),
	.V2C_10 (V2C_585_273),
	.V2C_11 (V2C_661_273),
	.V2C_12 (V2C_765_273),
	.V2C_13 (V2C_896_273),
	.V2C_14 (V2C_940_273),
	.V2C_15 (V2C_965_273),
	.V2C_16 (V2C_1025_273),
	.V2C_17 (V2C_1103_273),
	.V2C_18 (V2C_1148_273),
	.V2C_19 (V2C_1424_273),
	.V2C_20 (V2C_1425_273),
	.C2V_1 (C2V_273_6),
	.C2V_2 (C2V_273_81),
	.C2V_3 (C2V_273_98),
	.C2V_4 (C2V_273_180),
	.C2V_5 (C2V_273_198),
	.C2V_6 (C2V_273_265),
	.C2V_7 (C2V_273_362),
	.C2V_8 (C2V_273_417),
	.C2V_9 (C2V_273_576),
	.C2V_10 (C2V_273_585),
	.C2V_11 (C2V_273_661),
	.C2V_12 (C2V_273_765),
	.C2V_13 (C2V_273_896),
	.C2V_14 (C2V_273_940),
	.C2V_15 (C2V_273_965),
	.C2V_16 (C2V_273_1025),
	.C2V_17 (C2V_273_1103),
	.C2V_18 (C2V_273_1148),
	.C2V_19 (C2V_273_1424),
	.C2V_20 (C2V_273_1425),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU274 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_25_274),
	.V2C_2 (V2C_84_274),
	.V2C_3 (V2C_123_274),
	.V2C_4 (V2C_179_274),
	.V2C_5 (V2C_196_274),
	.V2C_6 (V2C_250_274),
	.V2C_7 (V2C_474_274),
	.V2C_8 (V2C_514_274),
	.V2C_9 (V2C_550_274),
	.V2C_10 (V2C_612_274),
	.V2C_11 (V2C_637_274),
	.V2C_12 (V2C_683_274),
	.V2C_13 (V2C_900_274),
	.V2C_14 (V2C_924_274),
	.V2C_15 (V2C_1008_274),
	.V2C_16 (V2C_1038_274),
	.V2C_17 (V2C_1065_274),
	.V2C_18 (V2C_1129_274),
	.V2C_19 (V2C_1425_274),
	.V2C_20 (V2C_1426_274),
	.C2V_1 (C2V_274_25),
	.C2V_2 (C2V_274_84),
	.C2V_3 (C2V_274_123),
	.C2V_4 (C2V_274_179),
	.C2V_5 (C2V_274_196),
	.C2V_6 (C2V_274_250),
	.C2V_7 (C2V_274_474),
	.C2V_8 (C2V_274_514),
	.C2V_9 (C2V_274_550),
	.C2V_10 (C2V_274_612),
	.C2V_11 (C2V_274_637),
	.C2V_12 (C2V_274_683),
	.C2V_13 (C2V_274_900),
	.C2V_14 (C2V_274_924),
	.C2V_15 (C2V_274_1008),
	.C2V_16 (C2V_274_1038),
	.C2V_17 (C2V_274_1065),
	.C2V_18 (C2V_274_1129),
	.C2V_19 (C2V_274_1425),
	.C2V_20 (C2V_274_1426),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU275 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_44_275),
	.V2C_2 (V2C_54_275),
	.V2C_3 (V2C_137_275),
	.V2C_4 (V2C_160_275),
	.V2C_5 (V2C_224_275),
	.V2C_6 (V2C_242_275),
	.V2C_7 (V2C_291_275),
	.V2C_8 (V2C_358_275),
	.V2C_9 (V2C_437_275),
	.V2C_10 (V2C_719_275),
	.V2C_11 (V2C_735_275),
	.V2C_12 (V2C_789_275),
	.V2C_13 (V2C_867_275),
	.V2C_14 (V2C_915_275),
	.V2C_15 (V2C_1006_275),
	.V2C_16 (V2C_1010_275),
	.V2C_17 (V2C_1059_275),
	.V2C_18 (V2C_1107_275),
	.V2C_19 (V2C_1426_275),
	.V2C_20 (V2C_1427_275),
	.C2V_1 (C2V_275_44),
	.C2V_2 (C2V_275_54),
	.C2V_3 (C2V_275_137),
	.C2V_4 (C2V_275_160),
	.C2V_5 (C2V_275_224),
	.C2V_6 (C2V_275_242),
	.C2V_7 (C2V_275_291),
	.C2V_8 (C2V_275_358),
	.C2V_9 (C2V_275_437),
	.C2V_10 (C2V_275_719),
	.C2V_11 (C2V_275_735),
	.C2V_12 (C2V_275_789),
	.C2V_13 (C2V_275_867),
	.C2V_14 (C2V_275_915),
	.C2V_15 (C2V_275_1006),
	.C2V_16 (C2V_275_1010),
	.C2V_17 (C2V_275_1059),
	.C2V_18 (C2V_275_1107),
	.C2V_19 (C2V_275_1426),
	.C2V_20 (C2V_275_1427),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU276 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_27_276),
	.V2C_2 (V2C_51_276),
	.V2C_3 (V2C_139_276),
	.V2C_4 (V2C_159_276),
	.V2C_5 (V2C_193_276),
	.V2C_6 (V2C_272_276),
	.V2C_7 (V2C_325_276),
	.V2C_8 (V2C_477_276),
	.V2C_9 (V2C_574_276),
	.V2C_10 (V2C_607_276),
	.V2C_11 (V2C_811_276),
	.V2C_12 (V2C_839_276),
	.V2C_13 (V2C_872_276),
	.V2C_14 (V2C_934_276),
	.V2C_15 (V2C_969_276),
	.V2C_16 (V2C_1036_276),
	.V2C_17 (V2C_1100_276),
	.V2C_18 (V2C_1150_276),
	.V2C_19 (V2C_1427_276),
	.V2C_20 (V2C_1428_276),
	.C2V_1 (C2V_276_27),
	.C2V_2 (C2V_276_51),
	.C2V_3 (C2V_276_139),
	.C2V_4 (C2V_276_159),
	.C2V_5 (C2V_276_193),
	.C2V_6 (C2V_276_272),
	.C2V_7 (C2V_276_325),
	.C2V_8 (C2V_276_477),
	.C2V_9 (C2V_276_574),
	.C2V_10 (C2V_276_607),
	.C2V_11 (C2V_276_811),
	.C2V_12 (C2V_276_839),
	.C2V_13 (C2V_276_872),
	.C2V_14 (C2V_276_934),
	.C2V_15 (C2V_276_969),
	.C2V_16 (C2V_276_1036),
	.C2V_17 (C2V_276_1100),
	.C2V_18 (C2V_276_1150),
	.C2V_19 (C2V_276_1427),
	.C2V_20 (C2V_276_1428),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU277 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_3_277),
	.V2C_2 (V2C_87_277),
	.V2C_3 (V2C_107_277),
	.V2C_4 (V2C_168_277),
	.V2C_5 (V2C_230_277),
	.V2C_6 (V2C_273_277),
	.V2C_7 (V2C_373_277),
	.V2C_8 (V2C_427_277),
	.V2C_9 (V2C_524_277),
	.V2C_10 (V2C_760_277),
	.V2C_11 (V2C_808_277),
	.V2C_12 (V2C_856_277),
	.V2C_13 (V2C_897_277),
	.V2C_14 (V2C_938_277),
	.V2C_15 (V2C_972_277),
	.V2C_16 (V2C_1011_277),
	.V2C_17 (V2C_1085_277),
	.V2C_18 (V2C_1144_277),
	.V2C_19 (V2C_1428_277),
	.V2C_20 (V2C_1429_277),
	.C2V_1 (C2V_277_3),
	.C2V_2 (C2V_277_87),
	.C2V_3 (C2V_277_107),
	.C2V_4 (C2V_277_168),
	.C2V_5 (C2V_277_230),
	.C2V_6 (C2V_277_273),
	.C2V_7 (C2V_277_373),
	.C2V_8 (C2V_277_427),
	.C2V_9 (C2V_277_524),
	.C2V_10 (C2V_277_760),
	.C2V_11 (C2V_277_808),
	.C2V_12 (C2V_277_856),
	.C2V_13 (C2V_277_897),
	.C2V_14 (C2V_277_938),
	.C2V_15 (C2V_277_972),
	.C2V_16 (C2V_277_1011),
	.C2V_17 (C2V_277_1085),
	.C2V_18 (C2V_277_1144),
	.C2V_19 (C2V_277_1428),
	.C2V_20 (C2V_277_1429),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU278 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_12_278),
	.V2C_2 (V2C_61_278),
	.V2C_3 (V2C_117_278),
	.V2C_4 (V2C_165_278),
	.V2C_5 (V2C_194_278),
	.V2C_6 (V2C_263_278),
	.V2C_7 (V2C_314_278),
	.V2C_8 (V2C_421_278),
	.V2C_9 (V2C_510_278),
	.V2C_10 (V2C_670_278),
	.V2C_11 (V2C_683_278),
	.V2C_12 (V2C_851_278),
	.V2C_13 (V2C_893_278),
	.V2C_14 (V2C_956_278),
	.V2C_15 (V2C_987_278),
	.V2C_16 (V2C_1019_278),
	.V2C_17 (V2C_1086_278),
	.V2C_18 (V2C_1117_278),
	.V2C_19 (V2C_1429_278),
	.V2C_20 (V2C_1430_278),
	.C2V_1 (C2V_278_12),
	.C2V_2 (C2V_278_61),
	.C2V_3 (C2V_278_117),
	.C2V_4 (C2V_278_165),
	.C2V_5 (C2V_278_194),
	.C2V_6 (C2V_278_263),
	.C2V_7 (C2V_278_314),
	.C2V_8 (C2V_278_421),
	.C2V_9 (C2V_278_510),
	.C2V_10 (C2V_278_670),
	.C2V_11 (C2V_278_683),
	.C2V_12 (C2V_278_851),
	.C2V_13 (C2V_278_893),
	.C2V_14 (C2V_278_956),
	.C2V_15 (C2V_278_987),
	.C2V_16 (C2V_278_1019),
	.C2V_17 (C2V_278_1086),
	.C2V_18 (C2V_278_1117),
	.C2V_19 (C2V_278_1429),
	.C2V_20 (C2V_278_1430),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU279 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_7_279),
	.V2C_2 (V2C_82_279),
	.V2C_3 (V2C_99_279),
	.V2C_4 (V2C_181_279),
	.V2C_5 (V2C_199_279),
	.V2C_6 (V2C_266_279),
	.V2C_7 (V2C_363_279),
	.V2C_8 (V2C_418_279),
	.V2C_9 (V2C_529_279),
	.V2C_10 (V2C_586_279),
	.V2C_11 (V2C_662_279),
	.V2C_12 (V2C_766_279),
	.V2C_13 (V2C_897_279),
	.V2C_14 (V2C_941_279),
	.V2C_15 (V2C_966_279),
	.V2C_16 (V2C_1026_279),
	.V2C_17 (V2C_1104_279),
	.V2C_18 (V2C_1149_279),
	.V2C_19 (V2C_1430_279),
	.V2C_20 (V2C_1431_279),
	.C2V_1 (C2V_279_7),
	.C2V_2 (C2V_279_82),
	.C2V_3 (C2V_279_99),
	.C2V_4 (C2V_279_181),
	.C2V_5 (C2V_279_199),
	.C2V_6 (C2V_279_266),
	.C2V_7 (C2V_279_363),
	.C2V_8 (C2V_279_418),
	.C2V_9 (C2V_279_529),
	.C2V_10 (C2V_279_586),
	.C2V_11 (C2V_279_662),
	.C2V_12 (C2V_279_766),
	.C2V_13 (C2V_279_897),
	.C2V_14 (C2V_279_941),
	.C2V_15 (C2V_279_966),
	.C2V_16 (C2V_279_1026),
	.C2V_17 (C2V_279_1104),
	.C2V_18 (C2V_279_1149),
	.C2V_19 (C2V_279_1430),
	.C2V_20 (C2V_279_1431),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU280 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_26_280),
	.V2C_2 (V2C_85_280),
	.V2C_3 (V2C_124_280),
	.V2C_4 (V2C_180_280),
	.V2C_5 (V2C_197_280),
	.V2C_6 (V2C_251_280),
	.V2C_7 (V2C_475_280),
	.V2C_8 (V2C_515_280),
	.V2C_9 (V2C_551_280),
	.V2C_10 (V2C_613_280),
	.V2C_11 (V2C_638_280),
	.V2C_12 (V2C_684_280),
	.V2C_13 (V2C_901_280),
	.V2C_14 (V2C_925_280),
	.V2C_15 (V2C_961_280),
	.V2C_16 (V2C_1039_280),
	.V2C_17 (V2C_1066_280),
	.V2C_18 (V2C_1130_280),
	.V2C_19 (V2C_1431_280),
	.V2C_20 (V2C_1432_280),
	.C2V_1 (C2V_280_26),
	.C2V_2 (C2V_280_85),
	.C2V_3 (C2V_280_124),
	.C2V_4 (C2V_280_180),
	.C2V_5 (C2V_280_197),
	.C2V_6 (C2V_280_251),
	.C2V_7 (C2V_280_475),
	.C2V_8 (C2V_280_515),
	.C2V_9 (C2V_280_551),
	.C2V_10 (C2V_280_613),
	.C2V_11 (C2V_280_638),
	.C2V_12 (C2V_280_684),
	.C2V_13 (C2V_280_901),
	.C2V_14 (C2V_280_925),
	.C2V_15 (C2V_280_961),
	.C2V_16 (C2V_280_1039),
	.C2V_17 (C2V_280_1066),
	.C2V_18 (C2V_280_1130),
	.C2V_19 (C2V_280_1431),
	.C2V_20 (C2V_280_1432),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU281 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_45_281),
	.V2C_2 (V2C_55_281),
	.V2C_3 (V2C_138_281),
	.V2C_4 (V2C_161_281),
	.V2C_5 (V2C_225_281),
	.V2C_6 (V2C_243_281),
	.V2C_7 (V2C_292_281),
	.V2C_8 (V2C_359_281),
	.V2C_9 (V2C_438_281),
	.V2C_10 (V2C_720_281),
	.V2C_11 (V2C_736_281),
	.V2C_12 (V2C_790_281),
	.V2C_13 (V2C_868_281),
	.V2C_14 (V2C_916_281),
	.V2C_15 (V2C_1007_281),
	.V2C_16 (V2C_1011_281),
	.V2C_17 (V2C_1060_281),
	.V2C_18 (V2C_1108_281),
	.V2C_19 (V2C_1432_281),
	.V2C_20 (V2C_1433_281),
	.C2V_1 (C2V_281_45),
	.C2V_2 (C2V_281_55),
	.C2V_3 (C2V_281_138),
	.C2V_4 (C2V_281_161),
	.C2V_5 (C2V_281_225),
	.C2V_6 (C2V_281_243),
	.C2V_7 (C2V_281_292),
	.C2V_8 (C2V_281_359),
	.C2V_9 (C2V_281_438),
	.C2V_10 (C2V_281_720),
	.C2V_11 (C2V_281_736),
	.C2V_12 (C2V_281_790),
	.C2V_13 (C2V_281_868),
	.C2V_14 (C2V_281_916),
	.C2V_15 (C2V_281_1007),
	.C2V_16 (C2V_281_1011),
	.C2V_17 (C2V_281_1060),
	.C2V_18 (C2V_281_1108),
	.C2V_19 (C2V_281_1432),
	.C2V_20 (C2V_281_1433),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU282 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_28_282),
	.V2C_2 (V2C_52_282),
	.V2C_3 (V2C_140_282),
	.V2C_4 (V2C_160_282),
	.V2C_5 (V2C_194_282),
	.V2C_6 (V2C_273_282),
	.V2C_7 (V2C_326_282),
	.V2C_8 (V2C_478_282),
	.V2C_9 (V2C_575_282),
	.V2C_10 (V2C_608_282),
	.V2C_11 (V2C_812_282),
	.V2C_12 (V2C_840_282),
	.V2C_13 (V2C_873_282),
	.V2C_14 (V2C_935_282),
	.V2C_15 (V2C_970_282),
	.V2C_16 (V2C_1037_282),
	.V2C_17 (V2C_1101_282),
	.V2C_18 (V2C_1151_282),
	.V2C_19 (V2C_1433_282),
	.V2C_20 (V2C_1434_282),
	.C2V_1 (C2V_282_28),
	.C2V_2 (C2V_282_52),
	.C2V_3 (C2V_282_140),
	.C2V_4 (C2V_282_160),
	.C2V_5 (C2V_282_194),
	.C2V_6 (C2V_282_273),
	.C2V_7 (C2V_282_326),
	.C2V_8 (C2V_282_478),
	.C2V_9 (C2V_282_575),
	.C2V_10 (C2V_282_608),
	.C2V_11 (C2V_282_812),
	.C2V_12 (C2V_282_840),
	.C2V_13 (C2V_282_873),
	.C2V_14 (C2V_282_935),
	.C2V_15 (C2V_282_970),
	.C2V_16 (C2V_282_1037),
	.C2V_17 (C2V_282_1101),
	.C2V_18 (C2V_282_1151),
	.C2V_19 (C2V_282_1433),
	.C2V_20 (C2V_282_1434),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU283 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_4_283),
	.V2C_2 (V2C_88_283),
	.V2C_3 (V2C_108_283),
	.V2C_4 (V2C_169_283),
	.V2C_5 (V2C_231_283),
	.V2C_6 (V2C_274_283),
	.V2C_7 (V2C_374_283),
	.V2C_8 (V2C_428_283),
	.V2C_9 (V2C_525_283),
	.V2C_10 (V2C_761_283),
	.V2C_11 (V2C_809_283),
	.V2C_12 (V2C_857_283),
	.V2C_13 (V2C_898_283),
	.V2C_14 (V2C_939_283),
	.V2C_15 (V2C_973_283),
	.V2C_16 (V2C_1012_283),
	.V2C_17 (V2C_1086_283),
	.V2C_18 (V2C_1145_283),
	.V2C_19 (V2C_1434_283),
	.V2C_20 (V2C_1435_283),
	.C2V_1 (C2V_283_4),
	.C2V_2 (C2V_283_88),
	.C2V_3 (C2V_283_108),
	.C2V_4 (C2V_283_169),
	.C2V_5 (C2V_283_231),
	.C2V_6 (C2V_283_274),
	.C2V_7 (C2V_283_374),
	.C2V_8 (C2V_283_428),
	.C2V_9 (C2V_283_525),
	.C2V_10 (C2V_283_761),
	.C2V_11 (C2V_283_809),
	.C2V_12 (C2V_283_857),
	.C2V_13 (C2V_283_898),
	.C2V_14 (C2V_283_939),
	.C2V_15 (C2V_283_973),
	.C2V_16 (C2V_283_1012),
	.C2V_17 (C2V_283_1086),
	.C2V_18 (C2V_283_1145),
	.C2V_19 (C2V_283_1434),
	.C2V_20 (C2V_283_1435),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU284 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_13_284),
	.V2C_2 (V2C_62_284),
	.V2C_3 (V2C_118_284),
	.V2C_4 (V2C_166_284),
	.V2C_5 (V2C_195_284),
	.V2C_6 (V2C_264_284),
	.V2C_7 (V2C_315_284),
	.V2C_8 (V2C_422_284),
	.V2C_9 (V2C_511_284),
	.V2C_10 (V2C_671_284),
	.V2C_11 (V2C_684_284),
	.V2C_12 (V2C_852_284),
	.V2C_13 (V2C_894_284),
	.V2C_14 (V2C_957_284),
	.V2C_15 (V2C_988_284),
	.V2C_16 (V2C_1020_284),
	.V2C_17 (V2C_1087_284),
	.V2C_18 (V2C_1118_284),
	.V2C_19 (V2C_1435_284),
	.V2C_20 (V2C_1436_284),
	.C2V_1 (C2V_284_13),
	.C2V_2 (C2V_284_62),
	.C2V_3 (C2V_284_118),
	.C2V_4 (C2V_284_166),
	.C2V_5 (C2V_284_195),
	.C2V_6 (C2V_284_264),
	.C2V_7 (C2V_284_315),
	.C2V_8 (C2V_284_422),
	.C2V_9 (C2V_284_511),
	.C2V_10 (C2V_284_671),
	.C2V_11 (C2V_284_684),
	.C2V_12 (C2V_284_852),
	.C2V_13 (C2V_284_894),
	.C2V_14 (C2V_284_957),
	.C2V_15 (C2V_284_988),
	.C2V_16 (C2V_284_1020),
	.C2V_17 (C2V_284_1087),
	.C2V_18 (C2V_284_1118),
	.C2V_19 (C2V_284_1435),
	.C2V_20 (C2V_284_1436),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU285 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_8_285),
	.V2C_2 (V2C_83_285),
	.V2C_3 (V2C_100_285),
	.V2C_4 (V2C_182_285),
	.V2C_5 (V2C_200_285),
	.V2C_6 (V2C_267_285),
	.V2C_7 (V2C_364_285),
	.V2C_8 (V2C_419_285),
	.V2C_9 (V2C_530_285),
	.V2C_10 (V2C_587_285),
	.V2C_11 (V2C_663_285),
	.V2C_12 (V2C_767_285),
	.V2C_13 (V2C_898_285),
	.V2C_14 (V2C_942_285),
	.V2C_15 (V2C_967_285),
	.V2C_16 (V2C_1027_285),
	.V2C_17 (V2C_1057_285),
	.V2C_18 (V2C_1150_285),
	.V2C_19 (V2C_1436_285),
	.V2C_20 (V2C_1437_285),
	.C2V_1 (C2V_285_8),
	.C2V_2 (C2V_285_83),
	.C2V_3 (C2V_285_100),
	.C2V_4 (C2V_285_182),
	.C2V_5 (C2V_285_200),
	.C2V_6 (C2V_285_267),
	.C2V_7 (C2V_285_364),
	.C2V_8 (C2V_285_419),
	.C2V_9 (C2V_285_530),
	.C2V_10 (C2V_285_587),
	.C2V_11 (C2V_285_663),
	.C2V_12 (C2V_285_767),
	.C2V_13 (C2V_285_898),
	.C2V_14 (C2V_285_942),
	.C2V_15 (C2V_285_967),
	.C2V_16 (C2V_285_1027),
	.C2V_17 (C2V_285_1057),
	.C2V_18 (C2V_285_1150),
	.C2V_19 (C2V_285_1436),
	.C2V_20 (C2V_285_1437),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU286 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_27_286),
	.V2C_2 (V2C_86_286),
	.V2C_3 (V2C_125_286),
	.V2C_4 (V2C_181_286),
	.V2C_5 (V2C_198_286),
	.V2C_6 (V2C_252_286),
	.V2C_7 (V2C_476_286),
	.V2C_8 (V2C_516_286),
	.V2C_9 (V2C_552_286),
	.V2C_10 (V2C_614_286),
	.V2C_11 (V2C_639_286),
	.V2C_12 (V2C_685_286),
	.V2C_13 (V2C_902_286),
	.V2C_14 (V2C_926_286),
	.V2C_15 (V2C_962_286),
	.V2C_16 (V2C_1040_286),
	.V2C_17 (V2C_1067_286),
	.V2C_18 (V2C_1131_286),
	.V2C_19 (V2C_1437_286),
	.V2C_20 (V2C_1438_286),
	.C2V_1 (C2V_286_27),
	.C2V_2 (C2V_286_86),
	.C2V_3 (C2V_286_125),
	.C2V_4 (C2V_286_181),
	.C2V_5 (C2V_286_198),
	.C2V_6 (C2V_286_252),
	.C2V_7 (C2V_286_476),
	.C2V_8 (C2V_286_516),
	.C2V_9 (C2V_286_552),
	.C2V_10 (C2V_286_614),
	.C2V_11 (C2V_286_639),
	.C2V_12 (C2V_286_685),
	.C2V_13 (C2V_286_902),
	.C2V_14 (C2V_286_926),
	.C2V_15 (C2V_286_962),
	.C2V_16 (C2V_286_1040),
	.C2V_17 (C2V_286_1067),
	.C2V_18 (C2V_286_1131),
	.C2V_19 (C2V_286_1437),
	.C2V_20 (C2V_286_1438),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU287 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_46_287),
	.V2C_2 (V2C_56_287),
	.V2C_3 (V2C_139_287),
	.V2C_4 (V2C_162_287),
	.V2C_5 (V2C_226_287),
	.V2C_6 (V2C_244_287),
	.V2C_7 (V2C_293_287),
	.V2C_8 (V2C_360_287),
	.V2C_9 (V2C_439_287),
	.V2C_10 (V2C_673_287),
	.V2C_11 (V2C_737_287),
	.V2C_12 (V2C_791_287),
	.V2C_13 (V2C_869_287),
	.V2C_14 (V2C_917_287),
	.V2C_15 (V2C_1008_287),
	.V2C_16 (V2C_1012_287),
	.V2C_17 (V2C_1061_287),
	.V2C_18 (V2C_1109_287),
	.V2C_19 (V2C_1438_287),
	.V2C_20 (V2C_1439_287),
	.C2V_1 (C2V_287_46),
	.C2V_2 (C2V_287_56),
	.C2V_3 (C2V_287_139),
	.C2V_4 (C2V_287_162),
	.C2V_5 (C2V_287_226),
	.C2V_6 (C2V_287_244),
	.C2V_7 (C2V_287_293),
	.C2V_8 (C2V_287_360),
	.C2V_9 (C2V_287_439),
	.C2V_10 (C2V_287_673),
	.C2V_11 (C2V_287_737),
	.C2V_12 (C2V_287_791),
	.C2V_13 (C2V_287_869),
	.C2V_14 (C2V_287_917),
	.C2V_15 (C2V_287_1008),
	.C2V_16 (C2V_287_1012),
	.C2V_17 (C2V_287_1061),
	.C2V_18 (C2V_287_1109),
	.C2V_19 (C2V_287_1438),
	.C2V_20 (C2V_287_1439),
	.init_cnt (8'd2)
);

CNU_20 #(quan_width) CNU288 (	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.V2C_1 (V2C_29_288),
	.V2C_2 (V2C_53_288),
	.V2C_3 (V2C_141_288),
	.V2C_4 (V2C_161_288),
	.V2C_5 (V2C_195_288),
	.V2C_6 (V2C_274_288),
	.V2C_7 (V2C_327_288),
	.V2C_8 (V2C_479_288),
	.V2C_9 (V2C_576_288),
	.V2C_10 (V2C_609_288),
	.V2C_11 (V2C_813_288),
	.V2C_12 (V2C_841_288),
	.V2C_13 (V2C_874_288),
	.V2C_14 (V2C_936_288),
	.V2C_15 (V2C_971_288),
	.V2C_16 (V2C_1038_288),
	.V2C_17 (V2C_1102_288),
	.V2C_18 (V2C_1152_288),
	.V2C_19 (V2C_1439_288),
	.V2C_20 (V2C_1440_288),
	.C2V_1 (C2V_288_29),
	.C2V_2 (C2V_288_53),
	.C2V_3 (C2V_288_141),
	.C2V_4 (C2V_288_161),
	.C2V_5 (C2V_288_195),
	.C2V_6 (C2V_288_274),
	.C2V_7 (C2V_288_327),
	.C2V_8 (C2V_288_479),
	.C2V_9 (C2V_288_576),
	.C2V_10 (C2V_288_609),
	.C2V_11 (C2V_288_813),
	.C2V_12 (C2V_288_841),
	.C2V_13 (C2V_288_874),
	.C2V_14 (C2V_288_936),
	.C2V_15 (C2V_288_971),
	.C2V_16 (C2V_288_1038),
	.C2V_17 (C2V_288_1102),
	.C2V_18 (C2V_288_1152),
	.C2V_19 (C2V_288_1439),
	.C2V_20 (C2V_288_1440),
	.init_cnt (8'd2)
);

VNU_6 #(quan_width) VNU1 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_1),
	.C2V_2 (C2V_120_1),
	.C2V_3 (C2V_130_1),
	.C2V_4 (C2V_212_1),
	.C2V_5 (C2V_243_1),
	.C2V_6 (C2V_265_1),
	.L (L_1),
	.V2C_1 (V2C_1_17),
	.V2C_2 (V2C_1_120),
	.V2C_3 (V2C_1_130),
	.V2C_4 (V2C_1_212),
	.V2C_5 (V2C_1_243),
	.V2C_6 (V2C_1_265),
	.V (V_1)
);

VNU_6 #(quan_width) VNU2 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_2),
	.C2V_2 (C2V_126_2),
	.C2V_3 (C2V_136_2),
	.C2V_4 (C2V_218_2),
	.C2V_5 (C2V_249_2),
	.C2V_6 (C2V_271_2),
	.L (L_2),
	.V2C_1 (V2C_2_23),
	.V2C_2 (V2C_2_126),
	.V2C_3 (V2C_2_136),
	.V2C_4 (V2C_2_218),
	.V2C_5 (V2C_2_249),
	.V2C_6 (V2C_2_271),
	.V (V_2)
);

VNU_6 #(quan_width) VNU3 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_3),
	.C2V_2 (C2V_132_3),
	.C2V_3 (C2V_142_3),
	.C2V_4 (C2V_224_3),
	.C2V_5 (C2V_255_3),
	.C2V_6 (C2V_277_3),
	.L (L_3),
	.V2C_1 (V2C_3_29),
	.V2C_2 (V2C_3_132),
	.V2C_3 (V2C_3_142),
	.V2C_4 (V2C_3_224),
	.V2C_5 (V2C_3_255),
	.V2C_6 (V2C_3_277),
	.V (V_3)
);

VNU_6 #(quan_width) VNU4 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_4),
	.C2V_2 (C2V_138_4),
	.C2V_3 (C2V_148_4),
	.C2V_4 (C2V_230_4),
	.C2V_5 (C2V_261_4),
	.C2V_6 (C2V_283_4),
	.L (L_4),
	.V2C_1 (V2C_4_35),
	.V2C_2 (V2C_4_138),
	.V2C_3 (V2C_4_148),
	.V2C_4 (V2C_4_230),
	.V2C_5 (V2C_4_261),
	.V2C_6 (V2C_4_283),
	.V (V_4)
);

VNU_6 #(quan_width) VNU5 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_5),
	.C2V_2 (C2V_41_5),
	.C2V_3 (C2V_144_5),
	.C2V_4 (C2V_154_5),
	.C2V_5 (C2V_236_5),
	.C2V_6 (C2V_267_5),
	.L (L_5),
	.V2C_1 (V2C_5_1),
	.V2C_2 (V2C_5_41),
	.V2C_3 (V2C_5_144),
	.V2C_4 (V2C_5_154),
	.V2C_5 (V2C_5_236),
	.V2C_6 (V2C_5_267),
	.V (V_5)
);

VNU_6 #(quan_width) VNU6 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_6),
	.C2V_2 (C2V_47_6),
	.C2V_3 (C2V_150_6),
	.C2V_4 (C2V_160_6),
	.C2V_5 (C2V_242_6),
	.C2V_6 (C2V_273_6),
	.L (L_6),
	.V2C_1 (V2C_6_7),
	.V2C_2 (V2C_6_47),
	.V2C_3 (V2C_6_150),
	.V2C_4 (V2C_6_160),
	.V2C_5 (V2C_6_242),
	.V2C_6 (V2C_6_273),
	.V (V_6)
);

VNU_6 #(quan_width) VNU7 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_7),
	.C2V_2 (C2V_53_7),
	.C2V_3 (C2V_156_7),
	.C2V_4 (C2V_166_7),
	.C2V_5 (C2V_248_7),
	.C2V_6 (C2V_279_7),
	.L (L_7),
	.V2C_1 (V2C_7_13),
	.V2C_2 (V2C_7_53),
	.V2C_3 (V2C_7_156),
	.V2C_4 (V2C_7_166),
	.V2C_5 (V2C_7_248),
	.V2C_6 (V2C_7_279),
	.V (V_7)
);

VNU_6 #(quan_width) VNU8 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_8),
	.C2V_2 (C2V_59_8),
	.C2V_3 (C2V_162_8),
	.C2V_4 (C2V_172_8),
	.C2V_5 (C2V_254_8),
	.C2V_6 (C2V_285_8),
	.L (L_8),
	.V2C_1 (V2C_8_19),
	.V2C_2 (V2C_8_59),
	.V2C_3 (V2C_8_162),
	.V2C_4 (V2C_8_172),
	.V2C_5 (V2C_8_254),
	.V2C_6 (V2C_8_285),
	.V (V_8)
);

VNU_6 #(quan_width) VNU9 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_9),
	.C2V_2 (C2V_25_9),
	.C2V_3 (C2V_65_9),
	.C2V_4 (C2V_168_9),
	.C2V_5 (C2V_178_9),
	.C2V_6 (C2V_260_9),
	.L (L_9),
	.V2C_1 (V2C_9_3),
	.V2C_2 (V2C_9_25),
	.V2C_3 (V2C_9_65),
	.V2C_4 (V2C_9_168),
	.V2C_5 (V2C_9_178),
	.V2C_6 (V2C_9_260),
	.V (V_9)
);

VNU_6 #(quan_width) VNU10 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_10),
	.C2V_2 (C2V_31_10),
	.C2V_3 (C2V_71_10),
	.C2V_4 (C2V_174_10),
	.C2V_5 (C2V_184_10),
	.C2V_6 (C2V_266_10),
	.L (L_10),
	.V2C_1 (V2C_10_9),
	.V2C_2 (V2C_10_31),
	.V2C_3 (V2C_10_71),
	.V2C_4 (V2C_10_174),
	.V2C_5 (V2C_10_184),
	.V2C_6 (V2C_10_266),
	.V (V_10)
);

VNU_6 #(quan_width) VNU11 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_11),
	.C2V_2 (C2V_37_11),
	.C2V_3 (C2V_77_11),
	.C2V_4 (C2V_180_11),
	.C2V_5 (C2V_190_11),
	.C2V_6 (C2V_272_11),
	.L (L_11),
	.V2C_1 (V2C_11_15),
	.V2C_2 (V2C_11_37),
	.V2C_3 (V2C_11_77),
	.V2C_4 (V2C_11_180),
	.V2C_5 (V2C_11_190),
	.V2C_6 (V2C_11_272),
	.V (V_11)
);

VNU_6 #(quan_width) VNU12 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_12),
	.C2V_2 (C2V_43_12),
	.C2V_3 (C2V_83_12),
	.C2V_4 (C2V_186_12),
	.C2V_5 (C2V_196_12),
	.C2V_6 (C2V_278_12),
	.L (L_12),
	.V2C_1 (V2C_12_21),
	.V2C_2 (V2C_12_43),
	.V2C_3 (V2C_12_83),
	.V2C_4 (V2C_12_186),
	.V2C_5 (V2C_12_196),
	.V2C_6 (V2C_12_278),
	.V (V_12)
);

VNU_6 #(quan_width) VNU13 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_13),
	.C2V_2 (C2V_49_13),
	.C2V_3 (C2V_89_13),
	.C2V_4 (C2V_192_13),
	.C2V_5 (C2V_202_13),
	.C2V_6 (C2V_284_13),
	.L (L_13),
	.V2C_1 (V2C_13_27),
	.V2C_2 (V2C_13_49),
	.V2C_3 (V2C_13_89),
	.V2C_4 (V2C_13_192),
	.V2C_5 (V2C_13_202),
	.V2C_6 (V2C_13_284),
	.V (V_13)
);

VNU_6 #(quan_width) VNU14 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_14),
	.C2V_2 (C2V_33_14),
	.C2V_3 (C2V_55_14),
	.C2V_4 (C2V_95_14),
	.C2V_5 (C2V_198_14),
	.C2V_6 (C2V_208_14),
	.L (L_14),
	.V2C_1 (V2C_14_2),
	.V2C_2 (V2C_14_33),
	.V2C_3 (V2C_14_55),
	.V2C_4 (V2C_14_95),
	.V2C_5 (V2C_14_198),
	.V2C_6 (V2C_14_208),
	.V (V_14)
);

VNU_6 #(quan_width) VNU15 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_15),
	.C2V_2 (C2V_39_15),
	.C2V_3 (C2V_61_15),
	.C2V_4 (C2V_101_15),
	.C2V_5 (C2V_204_15),
	.C2V_6 (C2V_214_15),
	.L (L_15),
	.V2C_1 (V2C_15_8),
	.V2C_2 (V2C_15_39),
	.V2C_3 (V2C_15_61),
	.V2C_4 (V2C_15_101),
	.V2C_5 (V2C_15_204),
	.V2C_6 (V2C_15_214),
	.V (V_15)
);

VNU_6 #(quan_width) VNU16 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_16),
	.C2V_2 (C2V_45_16),
	.C2V_3 (C2V_67_16),
	.C2V_4 (C2V_107_16),
	.C2V_5 (C2V_210_16),
	.C2V_6 (C2V_220_16),
	.L (L_16),
	.V2C_1 (V2C_16_14),
	.V2C_2 (V2C_16_45),
	.V2C_3 (V2C_16_67),
	.V2C_4 (V2C_16_107),
	.V2C_5 (V2C_16_210),
	.V2C_6 (V2C_16_220),
	.V (V_16)
);

VNU_6 #(quan_width) VNU17 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_17),
	.C2V_2 (C2V_51_17),
	.C2V_3 (C2V_73_17),
	.C2V_4 (C2V_113_17),
	.C2V_5 (C2V_216_17),
	.C2V_6 (C2V_226_17),
	.L (L_17),
	.V2C_1 (V2C_17_20),
	.V2C_2 (V2C_17_51),
	.V2C_3 (V2C_17_73),
	.V2C_4 (V2C_17_113),
	.V2C_5 (V2C_17_216),
	.V2C_6 (V2C_17_226),
	.V (V_17)
);

VNU_6 #(quan_width) VNU18 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_18),
	.C2V_2 (C2V_57_18),
	.C2V_3 (C2V_79_18),
	.C2V_4 (C2V_119_18),
	.C2V_5 (C2V_222_18),
	.C2V_6 (C2V_232_18),
	.L (L_18),
	.V2C_1 (V2C_18_26),
	.V2C_2 (V2C_18_57),
	.V2C_3 (V2C_18_79),
	.V2C_4 (V2C_18_119),
	.V2C_5 (V2C_18_222),
	.V2C_6 (V2C_18_232),
	.V (V_18)
);

VNU_6 #(quan_width) VNU19 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_19),
	.C2V_2 (C2V_63_19),
	.C2V_3 (C2V_85_19),
	.C2V_4 (C2V_125_19),
	.C2V_5 (C2V_228_19),
	.C2V_6 (C2V_238_19),
	.L (L_19),
	.V2C_1 (V2C_19_32),
	.V2C_2 (V2C_19_63),
	.V2C_3 (V2C_19_85),
	.V2C_4 (V2C_19_125),
	.V2C_5 (V2C_19_228),
	.V2C_6 (V2C_19_238),
	.V (V_19)
);

VNU_6 #(quan_width) VNU20 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_20),
	.C2V_2 (C2V_69_20),
	.C2V_3 (C2V_91_20),
	.C2V_4 (C2V_131_20),
	.C2V_5 (C2V_234_20),
	.C2V_6 (C2V_244_20),
	.L (L_20),
	.V2C_1 (V2C_20_38),
	.V2C_2 (V2C_20_69),
	.V2C_3 (V2C_20_91),
	.V2C_4 (V2C_20_131),
	.V2C_5 (V2C_20_234),
	.V2C_6 (V2C_20_244),
	.V (V_20)
);

VNU_6 #(quan_width) VNU21 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_21),
	.C2V_2 (C2V_75_21),
	.C2V_3 (C2V_97_21),
	.C2V_4 (C2V_137_21),
	.C2V_5 (C2V_240_21),
	.C2V_6 (C2V_250_21),
	.L (L_21),
	.V2C_1 (V2C_21_44),
	.V2C_2 (V2C_21_75),
	.V2C_3 (V2C_21_97),
	.V2C_4 (V2C_21_137),
	.V2C_5 (V2C_21_240),
	.V2C_6 (V2C_21_250),
	.V (V_21)
);

VNU_6 #(quan_width) VNU22 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_22),
	.C2V_2 (C2V_81_22),
	.C2V_3 (C2V_103_22),
	.C2V_4 (C2V_143_22),
	.C2V_5 (C2V_246_22),
	.C2V_6 (C2V_256_22),
	.L (L_22),
	.V2C_1 (V2C_22_50),
	.V2C_2 (V2C_22_81),
	.V2C_3 (V2C_22_103),
	.V2C_4 (V2C_22_143),
	.V2C_5 (V2C_22_246),
	.V2C_6 (V2C_22_256),
	.V (V_22)
);

VNU_6 #(quan_width) VNU23 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_23),
	.C2V_2 (C2V_87_23),
	.C2V_3 (C2V_109_23),
	.C2V_4 (C2V_149_23),
	.C2V_5 (C2V_252_23),
	.C2V_6 (C2V_262_23),
	.L (L_23),
	.V2C_1 (V2C_23_56),
	.V2C_2 (V2C_23_87),
	.V2C_3 (V2C_23_109),
	.V2C_4 (V2C_23_149),
	.V2C_5 (V2C_23_252),
	.V2C_6 (V2C_23_262),
	.V (V_23)
);

VNU_6 #(quan_width) VNU24 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_24),
	.C2V_2 (C2V_93_24),
	.C2V_3 (C2V_115_24),
	.C2V_4 (C2V_155_24),
	.C2V_5 (C2V_258_24),
	.C2V_6 (C2V_268_24),
	.L (L_24),
	.V2C_1 (V2C_24_62),
	.V2C_2 (V2C_24_93),
	.V2C_3 (V2C_24_115),
	.V2C_4 (V2C_24_155),
	.V2C_5 (V2C_24_258),
	.V2C_6 (V2C_24_268),
	.V (V_24)
);

VNU_6 #(quan_width) VNU25 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_25),
	.C2V_2 (C2V_99_25),
	.C2V_3 (C2V_121_25),
	.C2V_4 (C2V_161_25),
	.C2V_5 (C2V_264_25),
	.C2V_6 (C2V_274_25),
	.L (L_25),
	.V2C_1 (V2C_25_68),
	.V2C_2 (V2C_25_99),
	.V2C_3 (V2C_25_121),
	.V2C_4 (V2C_25_161),
	.V2C_5 (V2C_25_264),
	.V2C_6 (V2C_25_274),
	.V (V_25)
);

VNU_6 #(quan_width) VNU26 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_26),
	.C2V_2 (C2V_105_26),
	.C2V_3 (C2V_127_26),
	.C2V_4 (C2V_167_26),
	.C2V_5 (C2V_270_26),
	.C2V_6 (C2V_280_26),
	.L (L_26),
	.V2C_1 (V2C_26_74),
	.V2C_2 (V2C_26_105),
	.V2C_3 (V2C_26_127),
	.V2C_4 (V2C_26_167),
	.V2C_5 (V2C_26_270),
	.V2C_6 (V2C_26_280),
	.V (V_26)
);

VNU_6 #(quan_width) VNU27 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_80_27),
	.C2V_2 (C2V_111_27),
	.C2V_3 (C2V_133_27),
	.C2V_4 (C2V_173_27),
	.C2V_5 (C2V_276_27),
	.C2V_6 (C2V_286_27),
	.L (L_27),
	.V2C_1 (V2C_27_80),
	.V2C_2 (V2C_27_111),
	.V2C_3 (V2C_27_133),
	.V2C_4 (V2C_27_173),
	.V2C_5 (V2C_27_276),
	.V2C_6 (V2C_27_286),
	.V (V_27)
);

VNU_6 #(quan_width) VNU28 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_28),
	.C2V_2 (C2V_86_28),
	.C2V_3 (C2V_117_28),
	.C2V_4 (C2V_139_28),
	.C2V_5 (C2V_179_28),
	.C2V_6 (C2V_282_28),
	.L (L_28),
	.V2C_1 (V2C_28_4),
	.V2C_2 (V2C_28_86),
	.V2C_3 (V2C_28_117),
	.V2C_4 (V2C_28_139),
	.V2C_5 (V2C_28_179),
	.V2C_6 (V2C_28_282),
	.V (V_28)
);

VNU_6 #(quan_width) VNU29 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_29),
	.C2V_2 (C2V_92_29),
	.C2V_3 (C2V_123_29),
	.C2V_4 (C2V_145_29),
	.C2V_5 (C2V_185_29),
	.C2V_6 (C2V_288_29),
	.L (L_29),
	.V2C_1 (V2C_29_10),
	.V2C_2 (V2C_29_92),
	.V2C_3 (V2C_29_123),
	.V2C_4 (V2C_29_145),
	.V2C_5 (V2C_29_185),
	.V2C_6 (V2C_29_288),
	.V (V_29)
);

VNU_6 #(quan_width) VNU30 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_30),
	.C2V_2 (C2V_16_30),
	.C2V_3 (C2V_98_30),
	.C2V_4 (C2V_129_30),
	.C2V_5 (C2V_151_30),
	.C2V_6 (C2V_191_30),
	.L (L_30),
	.V2C_1 (V2C_30_6),
	.V2C_2 (V2C_30_16),
	.V2C_3 (V2C_30_98),
	.V2C_4 (V2C_30_129),
	.V2C_5 (V2C_30_151),
	.V2C_6 (V2C_30_191),
	.V (V_30)
);

VNU_6 #(quan_width) VNU31 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_31),
	.C2V_2 (C2V_22_31),
	.C2V_3 (C2V_104_31),
	.C2V_4 (C2V_135_31),
	.C2V_5 (C2V_157_31),
	.C2V_6 (C2V_197_31),
	.L (L_31),
	.V2C_1 (V2C_31_12),
	.V2C_2 (V2C_31_22),
	.V2C_3 (V2C_31_104),
	.V2C_4 (V2C_31_135),
	.V2C_5 (V2C_31_157),
	.V2C_6 (V2C_31_197),
	.V (V_31)
);

VNU_6 #(quan_width) VNU32 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_32),
	.C2V_2 (C2V_28_32),
	.C2V_3 (C2V_110_32),
	.C2V_4 (C2V_141_32),
	.C2V_5 (C2V_163_32),
	.C2V_6 (C2V_203_32),
	.L (L_32),
	.V2C_1 (V2C_32_18),
	.V2C_2 (V2C_32_28),
	.V2C_3 (V2C_32_110),
	.V2C_4 (V2C_32_141),
	.V2C_5 (V2C_32_163),
	.V2C_6 (V2C_32_203),
	.V (V_32)
);

VNU_6 #(quan_width) VNU33 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_33),
	.C2V_2 (C2V_34_33),
	.C2V_3 (C2V_116_33),
	.C2V_4 (C2V_147_33),
	.C2V_5 (C2V_169_33),
	.C2V_6 (C2V_209_33),
	.L (L_33),
	.V2C_1 (V2C_33_24),
	.V2C_2 (V2C_33_34),
	.V2C_3 (V2C_33_116),
	.V2C_4 (V2C_33_147),
	.V2C_5 (V2C_33_169),
	.V2C_6 (V2C_33_209),
	.V (V_33)
);

VNU_6 #(quan_width) VNU34 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_34),
	.C2V_2 (C2V_40_34),
	.C2V_3 (C2V_122_34),
	.C2V_4 (C2V_153_34),
	.C2V_5 (C2V_175_34),
	.C2V_6 (C2V_215_34),
	.L (L_34),
	.V2C_1 (V2C_34_30),
	.V2C_2 (V2C_34_40),
	.V2C_3 (V2C_34_122),
	.V2C_4 (V2C_34_153),
	.V2C_5 (V2C_34_175),
	.V2C_6 (V2C_34_215),
	.V (V_34)
);

VNU_6 #(quan_width) VNU35 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_35),
	.C2V_2 (C2V_46_35),
	.C2V_3 (C2V_128_35),
	.C2V_4 (C2V_159_35),
	.C2V_5 (C2V_181_35),
	.C2V_6 (C2V_221_35),
	.L (L_35),
	.V2C_1 (V2C_35_36),
	.V2C_2 (V2C_35_46),
	.V2C_3 (V2C_35_128),
	.V2C_4 (V2C_35_159),
	.V2C_5 (V2C_35_181),
	.V2C_6 (V2C_35_221),
	.V (V_35)
);

VNU_6 #(quan_width) VNU36 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_36),
	.C2V_2 (C2V_52_36),
	.C2V_3 (C2V_134_36),
	.C2V_4 (C2V_165_36),
	.C2V_5 (C2V_187_36),
	.C2V_6 (C2V_227_36),
	.L (L_36),
	.V2C_1 (V2C_36_42),
	.V2C_2 (V2C_36_52),
	.V2C_3 (V2C_36_134),
	.V2C_4 (V2C_36_165),
	.V2C_5 (V2C_36_187),
	.V2C_6 (V2C_36_227),
	.V (V_36)
);

VNU_6 #(quan_width) VNU37 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_37),
	.C2V_2 (C2V_58_37),
	.C2V_3 (C2V_140_37),
	.C2V_4 (C2V_171_37),
	.C2V_5 (C2V_193_37),
	.C2V_6 (C2V_233_37),
	.L (L_37),
	.V2C_1 (V2C_37_48),
	.V2C_2 (V2C_37_58),
	.V2C_3 (V2C_37_140),
	.V2C_4 (V2C_37_171),
	.V2C_5 (V2C_37_193),
	.V2C_6 (V2C_37_233),
	.V (V_37)
);

VNU_6 #(quan_width) VNU38 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_54_38),
	.C2V_2 (C2V_64_38),
	.C2V_3 (C2V_146_38),
	.C2V_4 (C2V_177_38),
	.C2V_5 (C2V_199_38),
	.C2V_6 (C2V_239_38),
	.L (L_38),
	.V2C_1 (V2C_38_54),
	.V2C_2 (V2C_38_64),
	.V2C_3 (V2C_38_146),
	.V2C_4 (V2C_38_177),
	.V2C_5 (V2C_38_199),
	.V2C_6 (V2C_38_239),
	.V (V_38)
);

VNU_6 #(quan_width) VNU39 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_60_39),
	.C2V_2 (C2V_70_39),
	.C2V_3 (C2V_152_39),
	.C2V_4 (C2V_183_39),
	.C2V_5 (C2V_205_39),
	.C2V_6 (C2V_245_39),
	.L (L_39),
	.V2C_1 (V2C_39_60),
	.V2C_2 (V2C_39_70),
	.V2C_3 (V2C_39_152),
	.V2C_4 (V2C_39_183),
	.V2C_5 (V2C_39_205),
	.V2C_6 (V2C_39_245),
	.V (V_39)
);

VNU_6 #(quan_width) VNU40 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_66_40),
	.C2V_2 (C2V_76_40),
	.C2V_3 (C2V_158_40),
	.C2V_4 (C2V_189_40),
	.C2V_5 (C2V_211_40),
	.C2V_6 (C2V_251_40),
	.L (L_40),
	.V2C_1 (V2C_40_66),
	.V2C_2 (V2C_40_76),
	.V2C_3 (V2C_40_158),
	.V2C_4 (V2C_40_189),
	.V2C_5 (V2C_40_211),
	.V2C_6 (V2C_40_251),
	.V (V_40)
);

VNU_6 #(quan_width) VNU41 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_72_41),
	.C2V_2 (C2V_82_41),
	.C2V_3 (C2V_164_41),
	.C2V_4 (C2V_195_41),
	.C2V_5 (C2V_217_41),
	.C2V_6 (C2V_257_41),
	.L (L_41),
	.V2C_1 (V2C_41_72),
	.V2C_2 (V2C_41_82),
	.V2C_3 (V2C_41_164),
	.V2C_4 (V2C_41_195),
	.V2C_5 (V2C_41_217),
	.V2C_6 (V2C_41_257),
	.V (V_41)
);

VNU_6 #(quan_width) VNU42 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_78_42),
	.C2V_2 (C2V_88_42),
	.C2V_3 (C2V_170_42),
	.C2V_4 (C2V_201_42),
	.C2V_5 (C2V_223_42),
	.C2V_6 (C2V_263_42),
	.L (L_42),
	.V2C_1 (V2C_42_78),
	.V2C_2 (V2C_42_88),
	.V2C_3 (V2C_42_170),
	.V2C_4 (V2C_42_201),
	.V2C_5 (V2C_42_223),
	.V2C_6 (V2C_42_263),
	.V (V_42)
);

VNU_6 #(quan_width) VNU43 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_84_43),
	.C2V_2 (C2V_94_43),
	.C2V_3 (C2V_176_43),
	.C2V_4 (C2V_207_43),
	.C2V_5 (C2V_229_43),
	.C2V_6 (C2V_269_43),
	.L (L_43),
	.V2C_1 (V2C_43_84),
	.V2C_2 (V2C_43_94),
	.V2C_3 (V2C_43_176),
	.V2C_4 (V2C_43_207),
	.V2C_5 (V2C_43_229),
	.V2C_6 (V2C_43_269),
	.V (V_43)
);

VNU_6 #(quan_width) VNU44 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_90_44),
	.C2V_2 (C2V_100_44),
	.C2V_3 (C2V_182_44),
	.C2V_4 (C2V_213_44),
	.C2V_5 (C2V_235_44),
	.C2V_6 (C2V_275_44),
	.L (L_44),
	.V2C_1 (V2C_44_90),
	.V2C_2 (V2C_44_100),
	.V2C_3 (V2C_44_182),
	.V2C_4 (V2C_44_213),
	.V2C_5 (V2C_44_235),
	.V2C_6 (V2C_44_275),
	.V (V_44)
);

VNU_6 #(quan_width) VNU45 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_96_45),
	.C2V_2 (C2V_106_45),
	.C2V_3 (C2V_188_45),
	.C2V_4 (C2V_219_45),
	.C2V_5 (C2V_241_45),
	.C2V_6 (C2V_281_45),
	.L (L_45),
	.V2C_1 (V2C_45_96),
	.V2C_2 (V2C_45_106),
	.V2C_3 (V2C_45_188),
	.V2C_4 (V2C_45_219),
	.V2C_5 (V2C_45_241),
	.V2C_6 (V2C_45_281),
	.V (V_45)
);

VNU_6 #(quan_width) VNU46 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_102_46),
	.C2V_2 (C2V_112_46),
	.C2V_3 (C2V_194_46),
	.C2V_4 (C2V_225_46),
	.C2V_5 (C2V_247_46),
	.C2V_6 (C2V_287_46),
	.L (L_46),
	.V2C_1 (V2C_46_102),
	.V2C_2 (V2C_46_112),
	.V2C_3 (V2C_46_194),
	.V2C_4 (V2C_46_225),
	.V2C_5 (V2C_46_247),
	.V2C_6 (V2C_46_287),
	.V (V_46)
);

VNU_6 #(quan_width) VNU47 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_47),
	.C2V_2 (C2V_108_47),
	.C2V_3 (C2V_118_47),
	.C2V_4 (C2V_200_47),
	.C2V_5 (C2V_231_47),
	.C2V_6 (C2V_253_47),
	.L (L_47),
	.V2C_1 (V2C_47_5),
	.V2C_2 (V2C_47_108),
	.V2C_3 (V2C_47_118),
	.V2C_4 (V2C_47_200),
	.V2C_5 (V2C_47_231),
	.V2C_6 (V2C_47_253),
	.V (V_47)
);

VNU_6 #(quan_width) VNU48 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_48),
	.C2V_2 (C2V_114_48),
	.C2V_3 (C2V_124_48),
	.C2V_4 (C2V_206_48),
	.C2V_5 (C2V_237_48),
	.C2V_6 (C2V_259_48),
	.L (L_48),
	.V2C_1 (V2C_48_11),
	.V2C_2 (V2C_48_114),
	.V2C_3 (V2C_48_124),
	.V2C_4 (V2C_48_206),
	.V2C_5 (V2C_48_237),
	.V2C_6 (V2C_48_259),
	.V (V_48)
);

VNU_6 #(quan_width) VNU49 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_49),
	.C2V_2 (C2V_64_49),
	.C2V_3 (C2V_81_49),
	.C2V_4 (C2V_206_49),
	.C2V_5 (C2V_245_49),
	.C2V_6 (C2V_264_49),
	.L (L_49),
	.V2C_1 (V2C_49_49),
	.V2C_2 (V2C_49_64),
	.V2C_3 (V2C_49_81),
	.V2C_4 (V2C_49_206),
	.V2C_5 (V2C_49_245),
	.V2C_6 (V2C_49_264),
	.V (V_49)
);

VNU_6 #(quan_width) VNU50 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_50),
	.C2V_2 (C2V_70_50),
	.C2V_3 (C2V_87_50),
	.C2V_4 (C2V_212_50),
	.C2V_5 (C2V_251_50),
	.C2V_6 (C2V_270_50),
	.L (L_50),
	.V2C_1 (V2C_50_55),
	.V2C_2 (V2C_50_70),
	.V2C_3 (V2C_50_87),
	.V2C_4 (V2C_50_212),
	.V2C_5 (V2C_50_251),
	.V2C_6 (V2C_50_270),
	.V (V_50)
);

VNU_6 #(quan_width) VNU51 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_51),
	.C2V_2 (C2V_76_51),
	.C2V_3 (C2V_93_51),
	.C2V_4 (C2V_218_51),
	.C2V_5 (C2V_257_51),
	.C2V_6 (C2V_276_51),
	.L (L_51),
	.V2C_1 (V2C_51_61),
	.V2C_2 (V2C_51_76),
	.V2C_3 (V2C_51_93),
	.V2C_4 (V2C_51_218),
	.V2C_5 (V2C_51_257),
	.V2C_6 (V2C_51_276),
	.V (V_51)
);

VNU_6 #(quan_width) VNU52 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_52),
	.C2V_2 (C2V_82_52),
	.C2V_3 (C2V_99_52),
	.C2V_4 (C2V_224_52),
	.C2V_5 (C2V_263_52),
	.C2V_6 (C2V_282_52),
	.L (L_52),
	.V2C_1 (V2C_52_67),
	.V2C_2 (V2C_52_82),
	.V2C_3 (V2C_52_99),
	.V2C_4 (V2C_52_224),
	.V2C_5 (V2C_52_263),
	.V2C_6 (V2C_52_282),
	.V (V_52)
);

VNU_6 #(quan_width) VNU53 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_53),
	.C2V_2 (C2V_88_53),
	.C2V_3 (C2V_105_53),
	.C2V_4 (C2V_230_53),
	.C2V_5 (C2V_269_53),
	.C2V_6 (C2V_288_53),
	.L (L_53),
	.V2C_1 (V2C_53_73),
	.V2C_2 (V2C_53_88),
	.V2C_3 (V2C_53_105),
	.V2C_4 (V2C_53_230),
	.V2C_5 (V2C_53_269),
	.V2C_6 (V2C_53_288),
	.V (V_53)
);

VNU_6 #(quan_width) VNU54 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_54),
	.C2V_2 (C2V_79_54),
	.C2V_3 (C2V_94_54),
	.C2V_4 (C2V_111_54),
	.C2V_5 (C2V_236_54),
	.C2V_6 (C2V_275_54),
	.L (L_54),
	.V2C_1 (V2C_54_6),
	.V2C_2 (V2C_54_79),
	.V2C_3 (V2C_54_94),
	.V2C_4 (V2C_54_111),
	.V2C_5 (V2C_54_236),
	.V2C_6 (V2C_54_275),
	.V (V_54)
);

VNU_6 #(quan_width) VNU55 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_55),
	.C2V_2 (C2V_85_55),
	.C2V_3 (C2V_100_55),
	.C2V_4 (C2V_117_55),
	.C2V_5 (C2V_242_55),
	.C2V_6 (C2V_281_55),
	.L (L_55),
	.V2C_1 (V2C_55_12),
	.V2C_2 (V2C_55_85),
	.V2C_3 (V2C_55_100),
	.V2C_4 (V2C_55_117),
	.V2C_5 (V2C_55_242),
	.V2C_6 (V2C_55_281),
	.V (V_55)
);

VNU_6 #(quan_width) VNU56 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_56),
	.C2V_2 (C2V_91_56),
	.C2V_3 (C2V_106_56),
	.C2V_4 (C2V_123_56),
	.C2V_5 (C2V_248_56),
	.C2V_6 (C2V_287_56),
	.L (L_56),
	.V2C_1 (V2C_56_18),
	.V2C_2 (V2C_56_91),
	.V2C_3 (V2C_56_106),
	.V2C_4 (V2C_56_123),
	.V2C_5 (V2C_56_248),
	.V2C_6 (V2C_56_287),
	.V (V_56)
);

VNU_6 #(quan_width) VNU57 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_57),
	.C2V_2 (C2V_24_57),
	.C2V_3 (C2V_97_57),
	.C2V_4 (C2V_112_57),
	.C2V_5 (C2V_129_57),
	.C2V_6 (C2V_254_57),
	.L (L_57),
	.V2C_1 (V2C_57_5),
	.V2C_2 (V2C_57_24),
	.V2C_3 (V2C_57_97),
	.V2C_4 (V2C_57_112),
	.V2C_5 (V2C_57_129),
	.V2C_6 (V2C_57_254),
	.V (V_57)
);

VNU_6 #(quan_width) VNU58 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_58),
	.C2V_2 (C2V_30_58),
	.C2V_3 (C2V_103_58),
	.C2V_4 (C2V_118_58),
	.C2V_5 (C2V_135_58),
	.C2V_6 (C2V_260_58),
	.L (L_58),
	.V2C_1 (V2C_58_11),
	.V2C_2 (V2C_58_30),
	.V2C_3 (V2C_58_103),
	.V2C_4 (V2C_58_118),
	.V2C_5 (V2C_58_135),
	.V2C_6 (V2C_58_260),
	.V (V_58)
);

VNU_6 #(quan_width) VNU59 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_59),
	.C2V_2 (C2V_36_59),
	.C2V_3 (C2V_109_59),
	.C2V_4 (C2V_124_59),
	.C2V_5 (C2V_141_59),
	.C2V_6 (C2V_266_59),
	.L (L_59),
	.V2C_1 (V2C_59_17),
	.V2C_2 (V2C_59_36),
	.V2C_3 (V2C_59_109),
	.V2C_4 (V2C_59_124),
	.V2C_5 (V2C_59_141),
	.V2C_6 (V2C_59_266),
	.V (V_59)
);

VNU_6 #(quan_width) VNU60 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_60),
	.C2V_2 (C2V_42_60),
	.C2V_3 (C2V_115_60),
	.C2V_4 (C2V_130_60),
	.C2V_5 (C2V_147_60),
	.C2V_6 (C2V_272_60),
	.L (L_60),
	.V2C_1 (V2C_60_23),
	.V2C_2 (V2C_60_42),
	.V2C_3 (V2C_60_115),
	.V2C_4 (V2C_60_130),
	.V2C_5 (V2C_60_147),
	.V2C_6 (V2C_60_272),
	.V (V_60)
);

VNU_6 #(quan_width) VNU61 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_61),
	.C2V_2 (C2V_48_61),
	.C2V_3 (C2V_121_61),
	.C2V_4 (C2V_136_61),
	.C2V_5 (C2V_153_61),
	.C2V_6 (C2V_278_61),
	.L (L_61),
	.V2C_1 (V2C_61_29),
	.V2C_2 (V2C_61_48),
	.V2C_3 (V2C_61_121),
	.V2C_4 (V2C_61_136),
	.V2C_5 (V2C_61_153),
	.V2C_6 (V2C_61_278),
	.V (V_61)
);

VNU_6 #(quan_width) VNU62 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_62),
	.C2V_2 (C2V_54_62),
	.C2V_3 (C2V_127_62),
	.C2V_4 (C2V_142_62),
	.C2V_5 (C2V_159_62),
	.C2V_6 (C2V_284_62),
	.L (L_62),
	.V2C_1 (V2C_62_35),
	.V2C_2 (V2C_62_54),
	.V2C_3 (V2C_62_127),
	.V2C_4 (V2C_62_142),
	.V2C_5 (V2C_62_159),
	.V2C_6 (V2C_62_284),
	.V (V_62)
);

VNU_6 #(quan_width) VNU63 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_63),
	.C2V_2 (C2V_41_63),
	.C2V_3 (C2V_60_63),
	.C2V_4 (C2V_133_63),
	.C2V_5 (C2V_148_63),
	.C2V_6 (C2V_165_63),
	.L (L_63),
	.V2C_1 (V2C_63_2),
	.V2C_2 (V2C_63_41),
	.V2C_3 (V2C_63_60),
	.V2C_4 (V2C_63_133),
	.V2C_5 (V2C_63_148),
	.V2C_6 (V2C_63_165),
	.V (V_63)
);

VNU_6 #(quan_width) VNU64 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_64),
	.C2V_2 (C2V_47_64),
	.C2V_3 (C2V_66_64),
	.C2V_4 (C2V_139_64),
	.C2V_5 (C2V_154_64),
	.C2V_6 (C2V_171_64),
	.L (L_64),
	.V2C_1 (V2C_64_8),
	.V2C_2 (V2C_64_47),
	.V2C_3 (V2C_64_66),
	.V2C_4 (V2C_64_139),
	.V2C_5 (V2C_64_154),
	.V2C_6 (V2C_64_171),
	.V (V_64)
);

VNU_6 #(quan_width) VNU65 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_65),
	.C2V_2 (C2V_53_65),
	.C2V_3 (C2V_72_65),
	.C2V_4 (C2V_145_65),
	.C2V_5 (C2V_160_65),
	.C2V_6 (C2V_177_65),
	.L (L_65),
	.V2C_1 (V2C_65_14),
	.V2C_2 (V2C_65_53),
	.V2C_3 (V2C_65_72),
	.V2C_4 (V2C_65_145),
	.V2C_5 (V2C_65_160),
	.V2C_6 (V2C_65_177),
	.V (V_65)
);

VNU_6 #(quan_width) VNU66 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_66),
	.C2V_2 (C2V_59_66),
	.C2V_3 (C2V_78_66),
	.C2V_4 (C2V_151_66),
	.C2V_5 (C2V_166_66),
	.C2V_6 (C2V_183_66),
	.L (L_66),
	.V2C_1 (V2C_66_20),
	.V2C_2 (V2C_66_59),
	.V2C_3 (V2C_66_78),
	.V2C_4 (V2C_66_151),
	.V2C_5 (V2C_66_166),
	.V2C_6 (V2C_66_183),
	.V (V_66)
);

VNU_6 #(quan_width) VNU67 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_67),
	.C2V_2 (C2V_65_67),
	.C2V_3 (C2V_84_67),
	.C2V_4 (C2V_157_67),
	.C2V_5 (C2V_172_67),
	.C2V_6 (C2V_189_67),
	.L (L_67),
	.V2C_1 (V2C_67_26),
	.V2C_2 (V2C_67_65),
	.V2C_3 (V2C_67_84),
	.V2C_4 (V2C_67_157),
	.V2C_5 (V2C_67_172),
	.V2C_6 (V2C_67_189),
	.V (V_67)
);

VNU_6 #(quan_width) VNU68 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_68),
	.C2V_2 (C2V_71_68),
	.C2V_3 (C2V_90_68),
	.C2V_4 (C2V_163_68),
	.C2V_5 (C2V_178_68),
	.C2V_6 (C2V_195_68),
	.L (L_68),
	.V2C_1 (V2C_68_32),
	.V2C_2 (V2C_68_71),
	.V2C_3 (V2C_68_90),
	.V2C_4 (V2C_68_163),
	.V2C_5 (V2C_68_178),
	.V2C_6 (V2C_68_195),
	.V (V_68)
);

VNU_6 #(quan_width) VNU69 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_69),
	.C2V_2 (C2V_77_69),
	.C2V_3 (C2V_96_69),
	.C2V_4 (C2V_169_69),
	.C2V_5 (C2V_184_69),
	.C2V_6 (C2V_201_69),
	.L (L_69),
	.V2C_1 (V2C_69_38),
	.V2C_2 (V2C_69_77),
	.V2C_3 (V2C_69_96),
	.V2C_4 (V2C_69_169),
	.V2C_5 (V2C_69_184),
	.V2C_6 (V2C_69_201),
	.V (V_69)
);

VNU_6 #(quan_width) VNU70 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_70),
	.C2V_2 (C2V_83_70),
	.C2V_3 (C2V_102_70),
	.C2V_4 (C2V_175_70),
	.C2V_5 (C2V_190_70),
	.C2V_6 (C2V_207_70),
	.L (L_70),
	.V2C_1 (V2C_70_44),
	.V2C_2 (V2C_70_83),
	.V2C_3 (V2C_70_102),
	.V2C_4 (V2C_70_175),
	.V2C_5 (V2C_70_190),
	.V2C_6 (V2C_70_207),
	.V (V_70)
);

VNU_6 #(quan_width) VNU71 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_71),
	.C2V_2 (C2V_89_71),
	.C2V_3 (C2V_108_71),
	.C2V_4 (C2V_181_71),
	.C2V_5 (C2V_196_71),
	.C2V_6 (C2V_213_71),
	.L (L_71),
	.V2C_1 (V2C_71_50),
	.V2C_2 (V2C_71_89),
	.V2C_3 (V2C_71_108),
	.V2C_4 (V2C_71_181),
	.V2C_5 (V2C_71_196),
	.V2C_6 (V2C_71_213),
	.V (V_71)
);

VNU_6 #(quan_width) VNU72 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_72),
	.C2V_2 (C2V_95_72),
	.C2V_3 (C2V_114_72),
	.C2V_4 (C2V_187_72),
	.C2V_5 (C2V_202_72),
	.C2V_6 (C2V_219_72),
	.L (L_72),
	.V2C_1 (V2C_72_56),
	.V2C_2 (V2C_72_95),
	.V2C_3 (V2C_72_114),
	.V2C_4 (V2C_72_187),
	.V2C_5 (V2C_72_202),
	.V2C_6 (V2C_72_219),
	.V (V_72)
);

VNU_6 #(quan_width) VNU73 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_73),
	.C2V_2 (C2V_101_73),
	.C2V_3 (C2V_120_73),
	.C2V_4 (C2V_193_73),
	.C2V_5 (C2V_208_73),
	.C2V_6 (C2V_225_73),
	.L (L_73),
	.V2C_1 (V2C_73_62),
	.V2C_2 (V2C_73_101),
	.V2C_3 (V2C_73_120),
	.V2C_4 (V2C_73_193),
	.V2C_5 (V2C_73_208),
	.V2C_6 (V2C_73_225),
	.V (V_73)
);

VNU_6 #(quan_width) VNU74 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_74),
	.C2V_2 (C2V_107_74),
	.C2V_3 (C2V_126_74),
	.C2V_4 (C2V_199_74),
	.C2V_5 (C2V_214_74),
	.C2V_6 (C2V_231_74),
	.L (L_74),
	.V2C_1 (V2C_74_68),
	.V2C_2 (V2C_74_107),
	.V2C_3 (V2C_74_126),
	.V2C_4 (V2C_74_199),
	.V2C_5 (V2C_74_214),
	.V2C_6 (V2C_74_231),
	.V (V_74)
);

VNU_6 #(quan_width) VNU75 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_75),
	.C2V_2 (C2V_113_75),
	.C2V_3 (C2V_132_75),
	.C2V_4 (C2V_205_75),
	.C2V_5 (C2V_220_75),
	.C2V_6 (C2V_237_75),
	.L (L_75),
	.V2C_1 (V2C_75_74),
	.V2C_2 (V2C_75_113),
	.V2C_3 (V2C_75_132),
	.V2C_4 (V2C_75_205),
	.V2C_5 (V2C_75_220),
	.V2C_6 (V2C_75_237),
	.V (V_75)
);

VNU_6 #(quan_width) VNU76 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_80_76),
	.C2V_2 (C2V_119_76),
	.C2V_3 (C2V_138_76),
	.C2V_4 (C2V_211_76),
	.C2V_5 (C2V_226_76),
	.C2V_6 (C2V_243_76),
	.L (L_76),
	.V2C_1 (V2C_76_80),
	.V2C_2 (V2C_76_119),
	.V2C_3 (V2C_76_138),
	.V2C_4 (V2C_76_211),
	.V2C_5 (V2C_76_226),
	.V2C_6 (V2C_76_243),
	.V (V_76)
);

VNU_6 #(quan_width) VNU77 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_86_77),
	.C2V_2 (C2V_125_77),
	.C2V_3 (C2V_144_77),
	.C2V_4 (C2V_217_77),
	.C2V_5 (C2V_232_77),
	.C2V_6 (C2V_249_77),
	.L (L_77),
	.V2C_1 (V2C_77_86),
	.V2C_2 (V2C_77_125),
	.V2C_3 (V2C_77_144),
	.V2C_4 (V2C_77_217),
	.V2C_5 (V2C_77_232),
	.V2C_6 (V2C_77_249),
	.V (V_77)
);

VNU_6 #(quan_width) VNU78 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_92_78),
	.C2V_2 (C2V_131_78),
	.C2V_3 (C2V_150_78),
	.C2V_4 (C2V_223_78),
	.C2V_5 (C2V_238_78),
	.C2V_6 (C2V_255_78),
	.L (L_78),
	.V2C_1 (V2C_78_92),
	.V2C_2 (V2C_78_131),
	.V2C_3 (V2C_78_150),
	.V2C_4 (V2C_78_223),
	.V2C_5 (V2C_78_238),
	.V2C_6 (V2C_78_255),
	.V (V_78)
);

VNU_6 #(quan_width) VNU79 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_98_79),
	.C2V_2 (C2V_137_79),
	.C2V_3 (C2V_156_79),
	.C2V_4 (C2V_229_79),
	.C2V_5 (C2V_244_79),
	.C2V_6 (C2V_261_79),
	.L (L_79),
	.V2C_1 (V2C_79_98),
	.V2C_2 (V2C_79_137),
	.V2C_3 (V2C_79_156),
	.V2C_4 (V2C_79_229),
	.V2C_5 (V2C_79_244),
	.V2C_6 (V2C_79_261),
	.V (V_79)
);

VNU_6 #(quan_width) VNU80 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_104_80),
	.C2V_2 (C2V_143_80),
	.C2V_3 (C2V_162_80),
	.C2V_4 (C2V_235_80),
	.C2V_5 (C2V_250_80),
	.C2V_6 (C2V_267_80),
	.L (L_80),
	.V2C_1 (V2C_80_104),
	.V2C_2 (V2C_80_143),
	.V2C_3 (V2C_80_162),
	.V2C_4 (V2C_80_235),
	.V2C_5 (V2C_80_250),
	.V2C_6 (V2C_80_267),
	.V (V_80)
);

VNU_6 #(quan_width) VNU81 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_110_81),
	.C2V_2 (C2V_149_81),
	.C2V_3 (C2V_168_81),
	.C2V_4 (C2V_241_81),
	.C2V_5 (C2V_256_81),
	.C2V_6 (C2V_273_81),
	.L (L_81),
	.V2C_1 (V2C_81_110),
	.V2C_2 (V2C_81_149),
	.V2C_3 (V2C_81_168),
	.V2C_4 (V2C_81_241),
	.V2C_5 (V2C_81_256),
	.V2C_6 (V2C_81_273),
	.V (V_81)
);

VNU_6 #(quan_width) VNU82 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_116_82),
	.C2V_2 (C2V_155_82),
	.C2V_3 (C2V_174_82),
	.C2V_4 (C2V_247_82),
	.C2V_5 (C2V_262_82),
	.C2V_6 (C2V_279_82),
	.L (L_82),
	.V2C_1 (V2C_82_116),
	.V2C_2 (V2C_82_155),
	.V2C_3 (V2C_82_174),
	.V2C_4 (V2C_82_247),
	.V2C_5 (V2C_82_262),
	.V2C_6 (V2C_82_279),
	.V (V_82)
);

VNU_6 #(quan_width) VNU83 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_122_83),
	.C2V_2 (C2V_161_83),
	.C2V_3 (C2V_180_83),
	.C2V_4 (C2V_253_83),
	.C2V_5 (C2V_268_83),
	.C2V_6 (C2V_285_83),
	.L (L_83),
	.V2C_1 (V2C_83_122),
	.V2C_2 (V2C_83_161),
	.V2C_3 (V2C_83_180),
	.V2C_4 (V2C_83_253),
	.V2C_5 (V2C_83_268),
	.V2C_6 (V2C_83_285),
	.V (V_83)
);

VNU_6 #(quan_width) VNU84 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_84),
	.C2V_2 (C2V_128_84),
	.C2V_3 (C2V_167_84),
	.C2V_4 (C2V_186_84),
	.C2V_5 (C2V_259_84),
	.C2V_6 (C2V_274_84),
	.L (L_84),
	.V2C_1 (V2C_84_3),
	.V2C_2 (V2C_84_128),
	.V2C_3 (V2C_84_167),
	.V2C_4 (V2C_84_186),
	.V2C_5 (V2C_84_259),
	.V2C_6 (V2C_84_274),
	.V (V_84)
);

VNU_6 #(quan_width) VNU85 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_85),
	.C2V_2 (C2V_134_85),
	.C2V_3 (C2V_173_85),
	.C2V_4 (C2V_192_85),
	.C2V_5 (C2V_265_85),
	.C2V_6 (C2V_280_85),
	.L (L_85),
	.V2C_1 (V2C_85_9),
	.V2C_2 (V2C_85_134),
	.V2C_3 (V2C_85_173),
	.V2C_4 (V2C_85_192),
	.V2C_5 (V2C_85_265),
	.V2C_6 (V2C_85_280),
	.V (V_85)
);

VNU_6 #(quan_width) VNU86 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_86),
	.C2V_2 (C2V_140_86),
	.C2V_3 (C2V_179_86),
	.C2V_4 (C2V_198_86),
	.C2V_5 (C2V_271_86),
	.C2V_6 (C2V_286_86),
	.L (L_86),
	.V2C_1 (V2C_86_15),
	.V2C_2 (V2C_86_140),
	.V2C_3 (V2C_86_179),
	.V2C_4 (V2C_86_198),
	.V2C_5 (V2C_86_271),
	.V2C_6 (V2C_86_286),
	.V (V_86)
);

VNU_6 #(quan_width) VNU87 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_87),
	.C2V_2 (C2V_21_87),
	.C2V_3 (C2V_146_87),
	.C2V_4 (C2V_185_87),
	.C2V_5 (C2V_204_87),
	.C2V_6 (C2V_277_87),
	.L (L_87),
	.V2C_1 (V2C_87_4),
	.V2C_2 (V2C_87_21),
	.V2C_3 (V2C_87_146),
	.V2C_4 (V2C_87_185),
	.V2C_5 (V2C_87_204),
	.V2C_6 (V2C_87_277),
	.V (V_87)
);

VNU_6 #(quan_width) VNU88 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_88),
	.C2V_2 (C2V_27_88),
	.C2V_3 (C2V_152_88),
	.C2V_4 (C2V_191_88),
	.C2V_5 (C2V_210_88),
	.C2V_6 (C2V_283_88),
	.L (L_88),
	.V2C_1 (V2C_88_10),
	.V2C_2 (V2C_88_27),
	.V2C_3 (V2C_88_152),
	.V2C_4 (V2C_88_191),
	.V2C_5 (V2C_88_210),
	.V2C_6 (V2C_88_283),
	.V (V_88)
);

VNU_6 #(quan_width) VNU89 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_89),
	.C2V_2 (C2V_16_89),
	.C2V_3 (C2V_33_89),
	.C2V_4 (C2V_158_89),
	.C2V_5 (C2V_197_89),
	.C2V_6 (C2V_216_89),
	.L (L_89),
	.V2C_1 (V2C_89_1),
	.V2C_2 (V2C_89_16),
	.V2C_3 (V2C_89_33),
	.V2C_4 (V2C_89_158),
	.V2C_5 (V2C_89_197),
	.V2C_6 (V2C_89_216),
	.V (V_89)
);

VNU_6 #(quan_width) VNU90 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_90),
	.C2V_2 (C2V_22_90),
	.C2V_3 (C2V_39_90),
	.C2V_4 (C2V_164_90),
	.C2V_5 (C2V_203_90),
	.C2V_6 (C2V_222_90),
	.L (L_90),
	.V2C_1 (V2C_90_7),
	.V2C_2 (V2C_90_22),
	.V2C_3 (V2C_90_39),
	.V2C_4 (V2C_90_164),
	.V2C_5 (V2C_90_203),
	.V2C_6 (V2C_90_222),
	.V (V_90)
);

VNU_6 #(quan_width) VNU91 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_91),
	.C2V_2 (C2V_28_91),
	.C2V_3 (C2V_45_91),
	.C2V_4 (C2V_170_91),
	.C2V_5 (C2V_209_91),
	.C2V_6 (C2V_228_91),
	.L (L_91),
	.V2C_1 (V2C_91_13),
	.V2C_2 (V2C_91_28),
	.V2C_3 (V2C_91_45),
	.V2C_4 (V2C_91_170),
	.V2C_5 (V2C_91_209),
	.V2C_6 (V2C_91_228),
	.V (V_91)
);

VNU_6 #(quan_width) VNU92 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_92),
	.C2V_2 (C2V_34_92),
	.C2V_3 (C2V_51_92),
	.C2V_4 (C2V_176_92),
	.C2V_5 (C2V_215_92),
	.C2V_6 (C2V_234_92),
	.L (L_92),
	.V2C_1 (V2C_92_19),
	.V2C_2 (V2C_92_34),
	.V2C_3 (V2C_92_51),
	.V2C_4 (V2C_92_176),
	.V2C_5 (V2C_92_215),
	.V2C_6 (V2C_92_234),
	.V (V_92)
);

VNU_6 #(quan_width) VNU93 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_93),
	.C2V_2 (C2V_40_93),
	.C2V_3 (C2V_57_93),
	.C2V_4 (C2V_182_93),
	.C2V_5 (C2V_221_93),
	.C2V_6 (C2V_240_93),
	.L (L_93),
	.V2C_1 (V2C_93_25),
	.V2C_2 (V2C_93_40),
	.V2C_3 (V2C_93_57),
	.V2C_4 (V2C_93_182),
	.V2C_5 (V2C_93_221),
	.V2C_6 (V2C_93_240),
	.V (V_93)
);

VNU_6 #(quan_width) VNU94 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_94),
	.C2V_2 (C2V_46_94),
	.C2V_3 (C2V_63_94),
	.C2V_4 (C2V_188_94),
	.C2V_5 (C2V_227_94),
	.C2V_6 (C2V_246_94),
	.L (L_94),
	.V2C_1 (V2C_94_31),
	.V2C_2 (V2C_94_46),
	.V2C_3 (V2C_94_63),
	.V2C_4 (V2C_94_188),
	.V2C_5 (V2C_94_227),
	.V2C_6 (V2C_94_246),
	.V (V_94)
);

VNU_6 #(quan_width) VNU95 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_95),
	.C2V_2 (C2V_52_95),
	.C2V_3 (C2V_69_95),
	.C2V_4 (C2V_194_95),
	.C2V_5 (C2V_233_95),
	.C2V_6 (C2V_252_95),
	.L (L_95),
	.V2C_1 (V2C_95_37),
	.V2C_2 (V2C_95_52),
	.V2C_3 (V2C_95_69),
	.V2C_4 (V2C_95_194),
	.V2C_5 (V2C_95_233),
	.V2C_6 (V2C_95_252),
	.V (V_95)
);

VNU_6 #(quan_width) VNU96 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_96),
	.C2V_2 (C2V_58_96),
	.C2V_3 (C2V_75_96),
	.C2V_4 (C2V_200_96),
	.C2V_5 (C2V_239_96),
	.C2V_6 (C2V_258_96),
	.L (L_96),
	.V2C_1 (V2C_96_43),
	.V2C_2 (V2C_96_58),
	.V2C_3 (V2C_96_75),
	.V2C_4 (V2C_96_200),
	.V2C_5 (V2C_96_239),
	.V2C_6 (V2C_96_258),
	.V (V_96)
);

VNU_6 #(quan_width) VNU97 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_97),
	.C2V_2 (C2V_35_97),
	.C2V_3 (C2V_118_97),
	.C2V_4 (C2V_158_97),
	.C2V_5 (C2V_217_97),
	.C2V_6 (C2V_267_97),
	.L (L_97),
	.V2C_1 (V2C_97_24),
	.V2C_2 (V2C_97_35),
	.V2C_3 (V2C_97_118),
	.V2C_4 (V2C_97_158),
	.V2C_5 (V2C_97_217),
	.V2C_6 (V2C_97_267),
	.V (V_97)
);

VNU_6 #(quan_width) VNU98 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_98),
	.C2V_2 (C2V_41_98),
	.C2V_3 (C2V_124_98),
	.C2V_4 (C2V_164_98),
	.C2V_5 (C2V_223_98),
	.C2V_6 (C2V_273_98),
	.L (L_98),
	.V2C_1 (V2C_98_30),
	.V2C_2 (V2C_98_41),
	.V2C_3 (V2C_98_124),
	.V2C_4 (V2C_98_164),
	.V2C_5 (V2C_98_223),
	.V2C_6 (V2C_98_273),
	.V (V_98)
);

VNU_6 #(quan_width) VNU99 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_99),
	.C2V_2 (C2V_47_99),
	.C2V_3 (C2V_130_99),
	.C2V_4 (C2V_170_99),
	.C2V_5 (C2V_229_99),
	.C2V_6 (C2V_279_99),
	.L (L_99),
	.V2C_1 (V2C_99_36),
	.V2C_2 (V2C_99_47),
	.V2C_3 (V2C_99_130),
	.V2C_4 (V2C_99_170),
	.V2C_5 (V2C_99_229),
	.V2C_6 (V2C_99_279),
	.V (V_99)
);

VNU_6 #(quan_width) VNU100 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_100),
	.C2V_2 (C2V_53_100),
	.C2V_3 (C2V_136_100),
	.C2V_4 (C2V_176_100),
	.C2V_5 (C2V_235_100),
	.C2V_6 (C2V_285_100),
	.L (L_100),
	.V2C_1 (V2C_100_42),
	.V2C_2 (V2C_100_53),
	.V2C_3 (V2C_100_136),
	.V2C_4 (V2C_100_176),
	.V2C_5 (V2C_100_235),
	.V2C_6 (V2C_100_285),
	.V (V_100)
);

VNU_6 #(quan_width) VNU101 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_101),
	.C2V_2 (C2V_48_101),
	.C2V_3 (C2V_59_101),
	.C2V_4 (C2V_142_101),
	.C2V_5 (C2V_182_101),
	.C2V_6 (C2V_241_101),
	.L (L_101),
	.V2C_1 (V2C_101_3),
	.V2C_2 (V2C_101_48),
	.V2C_3 (V2C_101_59),
	.V2C_4 (V2C_101_142),
	.V2C_5 (V2C_101_182),
	.V2C_6 (V2C_101_241),
	.V (V_101)
);

VNU_6 #(quan_width) VNU102 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_102),
	.C2V_2 (C2V_54_102),
	.C2V_3 (C2V_65_102),
	.C2V_4 (C2V_148_102),
	.C2V_5 (C2V_188_102),
	.C2V_6 (C2V_247_102),
	.L (L_102),
	.V2C_1 (V2C_102_9),
	.V2C_2 (V2C_102_54),
	.V2C_3 (V2C_102_65),
	.V2C_4 (V2C_102_148),
	.V2C_5 (V2C_102_188),
	.V2C_6 (V2C_102_247),
	.V (V_102)
);

VNU_6 #(quan_width) VNU103 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_103),
	.C2V_2 (C2V_60_103),
	.C2V_3 (C2V_71_103),
	.C2V_4 (C2V_154_103),
	.C2V_5 (C2V_194_103),
	.C2V_6 (C2V_253_103),
	.L (L_103),
	.V2C_1 (V2C_103_15),
	.V2C_2 (V2C_103_60),
	.V2C_3 (V2C_103_71),
	.V2C_4 (V2C_103_154),
	.V2C_5 (V2C_103_194),
	.V2C_6 (V2C_103_253),
	.V (V_103)
);

VNU_6 #(quan_width) VNU104 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_104),
	.C2V_2 (C2V_66_104),
	.C2V_3 (C2V_77_104),
	.C2V_4 (C2V_160_104),
	.C2V_5 (C2V_200_104),
	.C2V_6 (C2V_259_104),
	.L (L_104),
	.V2C_1 (V2C_104_21),
	.V2C_2 (V2C_104_66),
	.V2C_3 (V2C_104_77),
	.V2C_4 (V2C_104_160),
	.V2C_5 (V2C_104_200),
	.V2C_6 (V2C_104_259),
	.V (V_104)
);

VNU_6 #(quan_width) VNU105 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_105),
	.C2V_2 (C2V_72_105),
	.C2V_3 (C2V_83_105),
	.C2V_4 (C2V_166_105),
	.C2V_5 (C2V_206_105),
	.C2V_6 (C2V_265_105),
	.L (L_105),
	.V2C_1 (V2C_105_27),
	.V2C_2 (V2C_105_72),
	.V2C_3 (V2C_105_83),
	.V2C_4 (V2C_105_166),
	.V2C_5 (V2C_105_206),
	.V2C_6 (V2C_105_265),
	.V (V_105)
);

VNU_6 #(quan_width) VNU106 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_106),
	.C2V_2 (C2V_78_106),
	.C2V_3 (C2V_89_106),
	.C2V_4 (C2V_172_106),
	.C2V_5 (C2V_212_106),
	.C2V_6 (C2V_271_106),
	.L (L_106),
	.V2C_1 (V2C_106_33),
	.V2C_2 (V2C_106_78),
	.V2C_3 (V2C_106_89),
	.V2C_4 (V2C_106_172),
	.V2C_5 (V2C_106_212),
	.V2C_6 (V2C_106_271),
	.V (V_106)
);

VNU_6 #(quan_width) VNU107 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_107),
	.C2V_2 (C2V_84_107),
	.C2V_3 (C2V_95_107),
	.C2V_4 (C2V_178_107),
	.C2V_5 (C2V_218_107),
	.C2V_6 (C2V_277_107),
	.L (L_107),
	.V2C_1 (V2C_107_39),
	.V2C_2 (V2C_107_84),
	.V2C_3 (V2C_107_95),
	.V2C_4 (V2C_107_178),
	.V2C_5 (V2C_107_218),
	.V2C_6 (V2C_107_277),
	.V (V_107)
);

VNU_6 #(quan_width) VNU108 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_108),
	.C2V_2 (C2V_90_108),
	.C2V_3 (C2V_101_108),
	.C2V_4 (C2V_184_108),
	.C2V_5 (C2V_224_108),
	.C2V_6 (C2V_283_108),
	.L (L_108),
	.V2C_1 (V2C_108_45),
	.V2C_2 (V2C_108_90),
	.V2C_3 (V2C_108_101),
	.V2C_4 (V2C_108_184),
	.V2C_5 (V2C_108_224),
	.V2C_6 (V2C_108_283),
	.V (V_108)
);

VNU_6 #(quan_width) VNU109 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_109),
	.C2V_2 (C2V_51_109),
	.C2V_3 (C2V_96_109),
	.C2V_4 (C2V_107_109),
	.C2V_5 (C2V_190_109),
	.C2V_6 (C2V_230_109),
	.L (L_109),
	.V2C_1 (V2C_109_1),
	.V2C_2 (V2C_109_51),
	.V2C_3 (V2C_109_96),
	.V2C_4 (V2C_109_107),
	.V2C_5 (V2C_109_190),
	.V2C_6 (V2C_109_230),
	.V (V_109)
);

VNU_6 #(quan_width) VNU110 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_110),
	.C2V_2 (C2V_57_110),
	.C2V_3 (C2V_102_110),
	.C2V_4 (C2V_113_110),
	.C2V_5 (C2V_196_110),
	.C2V_6 (C2V_236_110),
	.L (L_110),
	.V2C_1 (V2C_110_7),
	.V2C_2 (V2C_110_57),
	.V2C_3 (V2C_110_102),
	.V2C_4 (V2C_110_113),
	.V2C_5 (V2C_110_196),
	.V2C_6 (V2C_110_236),
	.V (V_110)
);

VNU_6 #(quan_width) VNU111 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_111),
	.C2V_2 (C2V_63_111),
	.C2V_3 (C2V_108_111),
	.C2V_4 (C2V_119_111),
	.C2V_5 (C2V_202_111),
	.C2V_6 (C2V_242_111),
	.L (L_111),
	.V2C_1 (V2C_111_13),
	.V2C_2 (V2C_111_63),
	.V2C_3 (V2C_111_108),
	.V2C_4 (V2C_111_119),
	.V2C_5 (V2C_111_202),
	.V2C_6 (V2C_111_242),
	.V (V_111)
);

VNU_6 #(quan_width) VNU112 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_112),
	.C2V_2 (C2V_69_112),
	.C2V_3 (C2V_114_112),
	.C2V_4 (C2V_125_112),
	.C2V_5 (C2V_208_112),
	.C2V_6 (C2V_248_112),
	.L (L_112),
	.V2C_1 (V2C_112_19),
	.V2C_2 (V2C_112_69),
	.V2C_3 (V2C_112_114),
	.V2C_4 (V2C_112_125),
	.V2C_5 (V2C_112_208),
	.V2C_6 (V2C_112_248),
	.V (V_112)
);

VNU_6 #(quan_width) VNU113 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_113),
	.C2V_2 (C2V_75_113),
	.C2V_3 (C2V_120_113),
	.C2V_4 (C2V_131_113),
	.C2V_5 (C2V_214_113),
	.C2V_6 (C2V_254_113),
	.L (L_113),
	.V2C_1 (V2C_113_25),
	.V2C_2 (V2C_113_75),
	.V2C_3 (V2C_113_120),
	.V2C_4 (V2C_113_131),
	.V2C_5 (V2C_113_214),
	.V2C_6 (V2C_113_254),
	.V (V_113)
);

VNU_6 #(quan_width) VNU114 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_114),
	.C2V_2 (C2V_81_114),
	.C2V_3 (C2V_126_114),
	.C2V_4 (C2V_137_114),
	.C2V_5 (C2V_220_114),
	.C2V_6 (C2V_260_114),
	.L (L_114),
	.V2C_1 (V2C_114_31),
	.V2C_2 (V2C_114_81),
	.V2C_3 (V2C_114_126),
	.V2C_4 (V2C_114_137),
	.V2C_5 (V2C_114_220),
	.V2C_6 (V2C_114_260),
	.V (V_114)
);

VNU_6 #(quan_width) VNU115 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_115),
	.C2V_2 (C2V_87_115),
	.C2V_3 (C2V_132_115),
	.C2V_4 (C2V_143_115),
	.C2V_5 (C2V_226_115),
	.C2V_6 (C2V_266_115),
	.L (L_115),
	.V2C_1 (V2C_115_37),
	.V2C_2 (V2C_115_87),
	.V2C_3 (V2C_115_132),
	.V2C_4 (V2C_115_143),
	.V2C_5 (V2C_115_226),
	.V2C_6 (V2C_115_266),
	.V (V_115)
);

VNU_6 #(quan_width) VNU116 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_116),
	.C2V_2 (C2V_93_116),
	.C2V_3 (C2V_138_116),
	.C2V_4 (C2V_149_116),
	.C2V_5 (C2V_232_116),
	.C2V_6 (C2V_272_116),
	.L (L_116),
	.V2C_1 (V2C_116_43),
	.V2C_2 (V2C_116_93),
	.V2C_3 (V2C_116_138),
	.V2C_4 (V2C_116_149),
	.V2C_5 (V2C_116_232),
	.V2C_6 (V2C_116_272),
	.V (V_116)
);

VNU_6 #(quan_width) VNU117 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_117),
	.C2V_2 (C2V_99_117),
	.C2V_3 (C2V_144_117),
	.C2V_4 (C2V_155_117),
	.C2V_5 (C2V_238_117),
	.C2V_6 (C2V_278_117),
	.L (L_117),
	.V2C_1 (V2C_117_49),
	.V2C_2 (V2C_117_99),
	.V2C_3 (V2C_117_144),
	.V2C_4 (V2C_117_155),
	.V2C_5 (V2C_117_238),
	.V2C_6 (V2C_117_278),
	.V (V_117)
);

VNU_6 #(quan_width) VNU118 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_118),
	.C2V_2 (C2V_105_118),
	.C2V_3 (C2V_150_118),
	.C2V_4 (C2V_161_118),
	.C2V_5 (C2V_244_118),
	.C2V_6 (C2V_284_118),
	.L (L_118),
	.V2C_1 (V2C_118_55),
	.V2C_2 (V2C_118_105),
	.V2C_3 (V2C_118_150),
	.V2C_4 (V2C_118_161),
	.V2C_5 (V2C_118_244),
	.V2C_6 (V2C_118_284),
	.V (V_118)
);

VNU_6 #(quan_width) VNU119 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_119),
	.C2V_2 (C2V_61_119),
	.C2V_3 (C2V_111_119),
	.C2V_4 (C2V_156_119),
	.C2V_5 (C2V_167_119),
	.C2V_6 (C2V_250_119),
	.L (L_119),
	.V2C_1 (V2C_119_2),
	.V2C_2 (V2C_119_61),
	.V2C_3 (V2C_119_111),
	.V2C_4 (V2C_119_156),
	.V2C_5 (V2C_119_167),
	.V2C_6 (V2C_119_250),
	.V (V_119)
);

VNU_6 #(quan_width) VNU120 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_120),
	.C2V_2 (C2V_67_120),
	.C2V_3 (C2V_117_120),
	.C2V_4 (C2V_162_120),
	.C2V_5 (C2V_173_120),
	.C2V_6 (C2V_256_120),
	.L (L_120),
	.V2C_1 (V2C_120_8),
	.V2C_2 (V2C_120_67),
	.V2C_3 (V2C_120_117),
	.V2C_4 (V2C_120_162),
	.V2C_5 (V2C_120_173),
	.V2C_6 (V2C_120_256),
	.V (V_120)
);

VNU_6 #(quan_width) VNU121 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_121),
	.C2V_2 (C2V_73_121),
	.C2V_3 (C2V_123_121),
	.C2V_4 (C2V_168_121),
	.C2V_5 (C2V_179_121),
	.C2V_6 (C2V_262_121),
	.L (L_121),
	.V2C_1 (V2C_121_14),
	.V2C_2 (V2C_121_73),
	.V2C_3 (V2C_121_123),
	.V2C_4 (V2C_121_168),
	.V2C_5 (V2C_121_179),
	.V2C_6 (V2C_121_262),
	.V (V_121)
);

VNU_6 #(quan_width) VNU122 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_122),
	.C2V_2 (C2V_79_122),
	.C2V_3 (C2V_129_122),
	.C2V_4 (C2V_174_122),
	.C2V_5 (C2V_185_122),
	.C2V_6 (C2V_268_122),
	.L (L_122),
	.V2C_1 (V2C_122_20),
	.V2C_2 (V2C_122_79),
	.V2C_3 (V2C_122_129),
	.V2C_4 (V2C_122_174),
	.V2C_5 (V2C_122_185),
	.V2C_6 (V2C_122_268),
	.V (V_122)
);

VNU_6 #(quan_width) VNU123 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_123),
	.C2V_2 (C2V_85_123),
	.C2V_3 (C2V_135_123),
	.C2V_4 (C2V_180_123),
	.C2V_5 (C2V_191_123),
	.C2V_6 (C2V_274_123),
	.L (L_123),
	.V2C_1 (V2C_123_26),
	.V2C_2 (V2C_123_85),
	.V2C_3 (V2C_123_135),
	.V2C_4 (V2C_123_180),
	.V2C_5 (V2C_123_191),
	.V2C_6 (V2C_123_274),
	.V (V_123)
);

VNU_6 #(quan_width) VNU124 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_124),
	.C2V_2 (C2V_91_124),
	.C2V_3 (C2V_141_124),
	.C2V_4 (C2V_186_124),
	.C2V_5 (C2V_197_124),
	.C2V_6 (C2V_280_124),
	.L (L_124),
	.V2C_1 (V2C_124_32),
	.V2C_2 (V2C_124_91),
	.V2C_3 (V2C_124_141),
	.V2C_4 (V2C_124_186),
	.V2C_5 (V2C_124_197),
	.V2C_6 (V2C_124_280),
	.V (V_124)
);

VNU_6 #(quan_width) VNU125 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_125),
	.C2V_2 (C2V_97_125),
	.C2V_3 (C2V_147_125),
	.C2V_4 (C2V_192_125),
	.C2V_5 (C2V_203_125),
	.C2V_6 (C2V_286_125),
	.L (L_125),
	.V2C_1 (V2C_125_38),
	.V2C_2 (V2C_125_97),
	.V2C_3 (V2C_125_147),
	.V2C_4 (V2C_125_192),
	.V2C_5 (V2C_125_203),
	.V2C_6 (V2C_125_286),
	.V (V_125)
);

VNU_6 #(quan_width) VNU126 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_126),
	.C2V_2 (C2V_44_126),
	.C2V_3 (C2V_103_126),
	.C2V_4 (C2V_153_126),
	.C2V_5 (C2V_198_126),
	.C2V_6 (C2V_209_126),
	.L (L_126),
	.V2C_1 (V2C_126_4),
	.V2C_2 (V2C_126_44),
	.V2C_3 (V2C_126_103),
	.V2C_4 (V2C_126_153),
	.V2C_5 (V2C_126_198),
	.V2C_6 (V2C_126_209),
	.V (V_126)
);

VNU_6 #(quan_width) VNU127 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_127),
	.C2V_2 (C2V_50_127),
	.C2V_3 (C2V_109_127),
	.C2V_4 (C2V_159_127),
	.C2V_5 (C2V_204_127),
	.C2V_6 (C2V_215_127),
	.L (L_127),
	.V2C_1 (V2C_127_10),
	.V2C_2 (V2C_127_50),
	.V2C_3 (V2C_127_109),
	.V2C_4 (V2C_127_159),
	.V2C_5 (V2C_127_204),
	.V2C_6 (V2C_127_215),
	.V (V_127)
);

VNU_6 #(quan_width) VNU128 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_128),
	.C2V_2 (C2V_56_128),
	.C2V_3 (C2V_115_128),
	.C2V_4 (C2V_165_128),
	.C2V_5 (C2V_210_128),
	.C2V_6 (C2V_221_128),
	.L (L_128),
	.V2C_1 (V2C_128_16),
	.V2C_2 (V2C_128_56),
	.V2C_3 (V2C_128_115),
	.V2C_4 (V2C_128_165),
	.V2C_5 (V2C_128_210),
	.V2C_6 (V2C_128_221),
	.V (V_128)
);

VNU_6 #(quan_width) VNU129 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_129),
	.C2V_2 (C2V_62_129),
	.C2V_3 (C2V_121_129),
	.C2V_4 (C2V_171_129),
	.C2V_5 (C2V_216_129),
	.C2V_6 (C2V_227_129),
	.L (L_129),
	.V2C_1 (V2C_129_22),
	.V2C_2 (V2C_129_62),
	.V2C_3 (V2C_129_121),
	.V2C_4 (V2C_129_171),
	.V2C_5 (V2C_129_216),
	.V2C_6 (V2C_129_227),
	.V (V_129)
);

VNU_6 #(quan_width) VNU130 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_130),
	.C2V_2 (C2V_68_130),
	.C2V_3 (C2V_127_130),
	.C2V_4 (C2V_177_130),
	.C2V_5 (C2V_222_130),
	.C2V_6 (C2V_233_130),
	.L (L_130),
	.V2C_1 (V2C_130_28),
	.V2C_2 (V2C_130_68),
	.V2C_3 (V2C_130_127),
	.V2C_4 (V2C_130_177),
	.V2C_5 (V2C_130_222),
	.V2C_6 (V2C_130_233),
	.V (V_130)
);

VNU_6 #(quan_width) VNU131 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_131),
	.C2V_2 (C2V_74_131),
	.C2V_3 (C2V_133_131),
	.C2V_4 (C2V_183_131),
	.C2V_5 (C2V_228_131),
	.C2V_6 (C2V_239_131),
	.L (L_131),
	.V2C_1 (V2C_131_34),
	.V2C_2 (V2C_131_74),
	.V2C_3 (V2C_131_133),
	.V2C_4 (V2C_131_183),
	.V2C_5 (V2C_131_228),
	.V2C_6 (V2C_131_239),
	.V (V_131)
);

VNU_6 #(quan_width) VNU132 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_132),
	.C2V_2 (C2V_80_132),
	.C2V_3 (C2V_139_132),
	.C2V_4 (C2V_189_132),
	.C2V_5 (C2V_234_132),
	.C2V_6 (C2V_245_132),
	.L (L_132),
	.V2C_1 (V2C_132_40),
	.V2C_2 (V2C_132_80),
	.V2C_3 (V2C_132_139),
	.V2C_4 (V2C_132_189),
	.V2C_5 (V2C_132_234),
	.V2C_6 (V2C_132_245),
	.V (V_132)
);

VNU_6 #(quan_width) VNU133 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_133),
	.C2V_2 (C2V_86_133),
	.C2V_3 (C2V_145_133),
	.C2V_4 (C2V_195_133),
	.C2V_5 (C2V_240_133),
	.C2V_6 (C2V_251_133),
	.L (L_133),
	.V2C_1 (V2C_133_46),
	.V2C_2 (V2C_133_86),
	.V2C_3 (V2C_133_145),
	.V2C_4 (V2C_133_195),
	.V2C_5 (V2C_133_240),
	.V2C_6 (V2C_133_251),
	.V (V_133)
);

VNU_6 #(quan_width) VNU134 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_134),
	.C2V_2 (C2V_92_134),
	.C2V_3 (C2V_151_134),
	.C2V_4 (C2V_201_134),
	.C2V_5 (C2V_246_134),
	.C2V_6 (C2V_257_134),
	.L (L_134),
	.V2C_1 (V2C_134_52),
	.V2C_2 (V2C_134_92),
	.V2C_3 (V2C_134_151),
	.V2C_4 (V2C_134_201),
	.V2C_5 (V2C_134_246),
	.V2C_6 (V2C_134_257),
	.V (V_134)
);

VNU_6 #(quan_width) VNU135 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_135),
	.C2V_2 (C2V_98_135),
	.C2V_3 (C2V_157_135),
	.C2V_4 (C2V_207_135),
	.C2V_5 (C2V_252_135),
	.C2V_6 (C2V_263_135),
	.L (L_135),
	.V2C_1 (V2C_135_58),
	.V2C_2 (V2C_135_98),
	.V2C_3 (V2C_135_157),
	.V2C_4 (V2C_135_207),
	.V2C_5 (V2C_135_252),
	.V2C_6 (V2C_135_263),
	.V (V_135)
);

VNU_6 #(quan_width) VNU136 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_136),
	.C2V_2 (C2V_104_136),
	.C2V_3 (C2V_163_136),
	.C2V_4 (C2V_213_136),
	.C2V_5 (C2V_258_136),
	.C2V_6 (C2V_269_136),
	.L (L_136),
	.V2C_1 (V2C_136_64),
	.V2C_2 (V2C_136_104),
	.V2C_3 (V2C_136_163),
	.V2C_4 (V2C_136_213),
	.V2C_5 (V2C_136_258),
	.V2C_6 (V2C_136_269),
	.V (V_136)
);

VNU_6 #(quan_width) VNU137 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_137),
	.C2V_2 (C2V_110_137),
	.C2V_3 (C2V_169_137),
	.C2V_4 (C2V_219_137),
	.C2V_5 (C2V_264_137),
	.C2V_6 (C2V_275_137),
	.L (L_137),
	.V2C_1 (V2C_137_70),
	.V2C_2 (V2C_137_110),
	.V2C_3 (V2C_137_169),
	.V2C_4 (V2C_137_219),
	.V2C_5 (V2C_137_264),
	.V2C_6 (V2C_137_275),
	.V (V_137)
);

VNU_6 #(quan_width) VNU138 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_138),
	.C2V_2 (C2V_116_138),
	.C2V_3 (C2V_175_138),
	.C2V_4 (C2V_225_138),
	.C2V_5 (C2V_270_138),
	.C2V_6 (C2V_281_138),
	.L (L_138),
	.V2C_1 (V2C_138_76),
	.V2C_2 (V2C_138_116),
	.V2C_3 (V2C_138_175),
	.V2C_4 (V2C_138_225),
	.V2C_5 (V2C_138_270),
	.V2C_6 (V2C_138_281),
	.V (V_138)
);

VNU_6 #(quan_width) VNU139 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_139),
	.C2V_2 (C2V_122_139),
	.C2V_3 (C2V_181_139),
	.C2V_4 (C2V_231_139),
	.C2V_5 (C2V_276_139),
	.C2V_6 (C2V_287_139),
	.L (L_139),
	.V2C_1 (V2C_139_82),
	.V2C_2 (V2C_139_122),
	.V2C_3 (V2C_139_181),
	.V2C_4 (V2C_139_231),
	.V2C_5 (V2C_139_276),
	.V2C_6 (V2C_139_287),
	.V (V_139)
);

VNU_6 #(quan_width) VNU140 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_140),
	.C2V_2 (C2V_88_140),
	.C2V_3 (C2V_128_140),
	.C2V_4 (C2V_187_140),
	.C2V_5 (C2V_237_140),
	.C2V_6 (C2V_282_140),
	.L (L_140),
	.V2C_1 (V2C_140_5),
	.V2C_2 (V2C_140_88),
	.V2C_3 (V2C_140_128),
	.V2C_4 (V2C_140_187),
	.V2C_5 (V2C_140_237),
	.V2C_6 (V2C_140_282),
	.V (V_140)
);

VNU_6 #(quan_width) VNU141 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_141),
	.C2V_2 (C2V_94_141),
	.C2V_3 (C2V_134_141),
	.C2V_4 (C2V_193_141),
	.C2V_5 (C2V_243_141),
	.C2V_6 (C2V_288_141),
	.L (L_141),
	.V2C_1 (V2C_141_11),
	.V2C_2 (V2C_141_94),
	.V2C_3 (V2C_141_134),
	.V2C_4 (V2C_141_193),
	.V2C_5 (V2C_141_243),
	.V2C_6 (V2C_141_288),
	.V (V_141)
);

VNU_6 #(quan_width) VNU142 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_142),
	.C2V_2 (C2V_17_142),
	.C2V_3 (C2V_100_142),
	.C2V_4 (C2V_140_142),
	.C2V_5 (C2V_199_142),
	.C2V_6 (C2V_249_142),
	.L (L_142),
	.V2C_1 (V2C_142_6),
	.V2C_2 (V2C_142_17),
	.V2C_3 (V2C_142_100),
	.V2C_4 (V2C_142_140),
	.V2C_5 (V2C_142_199),
	.V2C_6 (V2C_142_249),
	.V (V_142)
);

VNU_6 #(quan_width) VNU143 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_143),
	.C2V_2 (C2V_23_143),
	.C2V_3 (C2V_106_143),
	.C2V_4 (C2V_146_143),
	.C2V_5 (C2V_205_143),
	.C2V_6 (C2V_255_143),
	.L (L_143),
	.V2C_1 (V2C_143_12),
	.V2C_2 (V2C_143_23),
	.V2C_3 (V2C_143_106),
	.V2C_4 (V2C_143_146),
	.V2C_5 (V2C_143_205),
	.V2C_6 (V2C_143_255),
	.V (V_143)
);

VNU_6 #(quan_width) VNU144 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_144),
	.C2V_2 (C2V_29_144),
	.C2V_3 (C2V_112_144),
	.C2V_4 (C2V_152_144),
	.C2V_5 (C2V_211_144),
	.C2V_6 (C2V_261_144),
	.L (L_144),
	.V2C_1 (V2C_144_18),
	.V2C_2 (V2C_144_29),
	.V2C_3 (V2C_144_112),
	.V2C_4 (V2C_144_152),
	.V2C_5 (V2C_144_211),
	.V2C_6 (V2C_144_261),
	.V (V_144)
);

VNU_6 #(quan_width) VNU145 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_145),
	.C2V_2 (C2V_70_145),
	.C2V_3 (C2V_139_145),
	.C2V_4 (C2V_158_145),
	.C2V_5 (C2V_185_145),
	.C2V_6 (C2V_192_145),
	.L (L_145),
	.V2C_1 (V2C_145_63),
	.V2C_2 (V2C_145_70),
	.V2C_3 (V2C_145_139),
	.V2C_4 (V2C_145_158),
	.V2C_5 (V2C_145_185),
	.V2C_6 (V2C_145_192),
	.V (V_145)
);

VNU_6 #(quan_width) VNU146 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_146),
	.C2V_2 (C2V_76_146),
	.C2V_3 (C2V_145_146),
	.C2V_4 (C2V_164_146),
	.C2V_5 (C2V_191_146),
	.C2V_6 (C2V_198_146),
	.L (L_146),
	.V2C_1 (V2C_146_69),
	.V2C_2 (V2C_146_76),
	.V2C_3 (V2C_146_145),
	.V2C_4 (V2C_146_164),
	.V2C_5 (V2C_146_191),
	.V2C_6 (V2C_146_198),
	.V (V_146)
);

VNU_6 #(quan_width) VNU147 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_147),
	.C2V_2 (C2V_82_147),
	.C2V_3 (C2V_151_147),
	.C2V_4 (C2V_170_147),
	.C2V_5 (C2V_197_147),
	.C2V_6 (C2V_204_147),
	.L (L_147),
	.V2C_1 (V2C_147_75),
	.V2C_2 (V2C_147_82),
	.V2C_3 (V2C_147_151),
	.V2C_4 (V2C_147_170),
	.V2C_5 (V2C_147_197),
	.V2C_6 (V2C_147_204),
	.V (V_147)
);

VNU_6 #(quan_width) VNU148 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_148),
	.C2V_2 (C2V_88_148),
	.C2V_3 (C2V_157_148),
	.C2V_4 (C2V_176_148),
	.C2V_5 (C2V_203_148),
	.C2V_6 (C2V_210_148),
	.L (L_148),
	.V2C_1 (V2C_148_81),
	.V2C_2 (V2C_148_88),
	.V2C_3 (V2C_148_157),
	.V2C_4 (V2C_148_176),
	.V2C_5 (V2C_148_203),
	.V2C_6 (V2C_148_210),
	.V (V_148)
);

VNU_6 #(quan_width) VNU149 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_149),
	.C2V_2 (C2V_94_149),
	.C2V_3 (C2V_163_149),
	.C2V_4 (C2V_182_149),
	.C2V_5 (C2V_209_149),
	.C2V_6 (C2V_216_149),
	.L (L_149),
	.V2C_1 (V2C_149_87),
	.V2C_2 (V2C_149_94),
	.V2C_3 (V2C_149_163),
	.V2C_4 (V2C_149_182),
	.V2C_5 (V2C_149_209),
	.V2C_6 (V2C_149_216),
	.V (V_149)
);

VNU_6 #(quan_width) VNU150 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_93_150),
	.C2V_2 (C2V_100_150),
	.C2V_3 (C2V_169_150),
	.C2V_4 (C2V_188_150),
	.C2V_5 (C2V_215_150),
	.C2V_6 (C2V_222_150),
	.L (L_150),
	.V2C_1 (V2C_150_93),
	.V2C_2 (V2C_150_100),
	.V2C_3 (V2C_150_169),
	.V2C_4 (V2C_150_188),
	.V2C_5 (V2C_150_215),
	.V2C_6 (V2C_150_222),
	.V (V_150)
);

VNU_6 #(quan_width) VNU151 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_99_151),
	.C2V_2 (C2V_106_151),
	.C2V_3 (C2V_175_151),
	.C2V_4 (C2V_194_151),
	.C2V_5 (C2V_221_151),
	.C2V_6 (C2V_228_151),
	.L (L_151),
	.V2C_1 (V2C_151_99),
	.V2C_2 (V2C_151_106),
	.V2C_3 (V2C_151_175),
	.V2C_4 (V2C_151_194),
	.V2C_5 (V2C_151_221),
	.V2C_6 (V2C_151_228),
	.V (V_151)
);

VNU_6 #(quan_width) VNU152 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_105_152),
	.C2V_2 (C2V_112_152),
	.C2V_3 (C2V_181_152),
	.C2V_4 (C2V_200_152),
	.C2V_5 (C2V_227_152),
	.C2V_6 (C2V_234_152),
	.L (L_152),
	.V2C_1 (V2C_152_105),
	.V2C_2 (V2C_152_112),
	.V2C_3 (V2C_152_181),
	.V2C_4 (V2C_152_200),
	.V2C_5 (V2C_152_227),
	.V2C_6 (V2C_152_234),
	.V (V_152)
);

VNU_6 #(quan_width) VNU153 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_111_153),
	.C2V_2 (C2V_118_153),
	.C2V_3 (C2V_187_153),
	.C2V_4 (C2V_206_153),
	.C2V_5 (C2V_233_153),
	.C2V_6 (C2V_240_153),
	.L (L_153),
	.V2C_1 (V2C_153_111),
	.V2C_2 (V2C_153_118),
	.V2C_3 (V2C_153_187),
	.V2C_4 (V2C_153_206),
	.V2C_5 (V2C_153_233),
	.V2C_6 (V2C_153_240),
	.V (V_153)
);

VNU_6 #(quan_width) VNU154 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_117_154),
	.C2V_2 (C2V_124_154),
	.C2V_3 (C2V_193_154),
	.C2V_4 (C2V_212_154),
	.C2V_5 (C2V_239_154),
	.C2V_6 (C2V_246_154),
	.L (L_154),
	.V2C_1 (V2C_154_117),
	.V2C_2 (V2C_154_124),
	.V2C_3 (V2C_154_193),
	.V2C_4 (V2C_154_212),
	.V2C_5 (V2C_154_239),
	.V2C_6 (V2C_154_246),
	.V (V_154)
);

VNU_6 #(quan_width) VNU155 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_123_155),
	.C2V_2 (C2V_130_155),
	.C2V_3 (C2V_199_155),
	.C2V_4 (C2V_218_155),
	.C2V_5 (C2V_245_155),
	.C2V_6 (C2V_252_155),
	.L (L_155),
	.V2C_1 (V2C_155_123),
	.V2C_2 (V2C_155_130),
	.V2C_3 (V2C_155_199),
	.V2C_4 (V2C_155_218),
	.V2C_5 (V2C_155_245),
	.V2C_6 (V2C_155_252),
	.V (V_155)
);

VNU_6 #(quan_width) VNU156 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_129_156),
	.C2V_2 (C2V_136_156),
	.C2V_3 (C2V_205_156),
	.C2V_4 (C2V_224_156),
	.C2V_5 (C2V_251_156),
	.C2V_6 (C2V_258_156),
	.L (L_156),
	.V2C_1 (V2C_156_129),
	.V2C_2 (V2C_156_136),
	.V2C_3 (V2C_156_205),
	.V2C_4 (V2C_156_224),
	.V2C_5 (V2C_156_251),
	.V2C_6 (V2C_156_258),
	.V (V_156)
);

VNU_6 #(quan_width) VNU157 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_135_157),
	.C2V_2 (C2V_142_157),
	.C2V_3 (C2V_211_157),
	.C2V_4 (C2V_230_157),
	.C2V_5 (C2V_257_157),
	.C2V_6 (C2V_264_157),
	.L (L_157),
	.V2C_1 (V2C_157_135),
	.V2C_2 (V2C_157_142),
	.V2C_3 (V2C_157_211),
	.V2C_4 (V2C_157_230),
	.V2C_5 (V2C_157_257),
	.V2C_6 (V2C_157_264),
	.V (V_157)
);

VNU_6 #(quan_width) VNU158 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_141_158),
	.C2V_2 (C2V_148_158),
	.C2V_3 (C2V_217_158),
	.C2V_4 (C2V_236_158),
	.C2V_5 (C2V_263_158),
	.C2V_6 (C2V_270_158),
	.L (L_158),
	.V2C_1 (V2C_158_141),
	.V2C_2 (V2C_158_148),
	.V2C_3 (V2C_158_217),
	.V2C_4 (V2C_158_236),
	.V2C_5 (V2C_158_263),
	.V2C_6 (V2C_158_270),
	.V (V_158)
);

VNU_6 #(quan_width) VNU159 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_147_159),
	.C2V_2 (C2V_154_159),
	.C2V_3 (C2V_223_159),
	.C2V_4 (C2V_242_159),
	.C2V_5 (C2V_269_159),
	.C2V_6 (C2V_276_159),
	.L (L_159),
	.V2C_1 (V2C_159_147),
	.V2C_2 (V2C_159_154),
	.V2C_3 (V2C_159_223),
	.V2C_4 (V2C_159_242),
	.V2C_5 (V2C_159_269),
	.V2C_6 (V2C_159_276),
	.V (V_159)
);

VNU_6 #(quan_width) VNU160 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_153_160),
	.C2V_2 (C2V_160_160),
	.C2V_3 (C2V_229_160),
	.C2V_4 (C2V_248_160),
	.C2V_5 (C2V_275_160),
	.C2V_6 (C2V_282_160),
	.L (L_160),
	.V2C_1 (V2C_160_153),
	.V2C_2 (V2C_160_160),
	.V2C_3 (V2C_160_229),
	.V2C_4 (V2C_160_248),
	.V2C_5 (V2C_160_275),
	.V2C_6 (V2C_160_282),
	.V (V_160)
);

VNU_6 #(quan_width) VNU161 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_159_161),
	.C2V_2 (C2V_166_161),
	.C2V_3 (C2V_235_161),
	.C2V_4 (C2V_254_161),
	.C2V_5 (C2V_281_161),
	.C2V_6 (C2V_288_161),
	.L (L_161),
	.V2C_1 (V2C_161_159),
	.V2C_2 (V2C_161_166),
	.V2C_3 (V2C_161_235),
	.V2C_4 (V2C_161_254),
	.V2C_5 (V2C_161_281),
	.V2C_6 (V2C_161_288),
	.V (V_161)
);

VNU_6 #(quan_width) VNU162 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_162),
	.C2V_2 (C2V_165_162),
	.C2V_3 (C2V_172_162),
	.C2V_4 (C2V_241_162),
	.C2V_5 (C2V_260_162),
	.C2V_6 (C2V_287_162),
	.L (L_162),
	.V2C_1 (V2C_162_6),
	.V2C_2 (V2C_162_165),
	.V2C_3 (V2C_162_172),
	.V2C_4 (V2C_162_241),
	.V2C_5 (V2C_162_260),
	.V2C_6 (V2C_162_287),
	.V (V_162)
);

VNU_6 #(quan_width) VNU163 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_163),
	.C2V_2 (C2V_12_163),
	.C2V_3 (C2V_171_163),
	.C2V_4 (C2V_178_163),
	.C2V_5 (C2V_247_163),
	.C2V_6 (C2V_266_163),
	.L (L_163),
	.V2C_1 (V2C_163_5),
	.V2C_2 (V2C_163_12),
	.V2C_3 (V2C_163_171),
	.V2C_4 (V2C_163_178),
	.V2C_5 (V2C_163_247),
	.V2C_6 (V2C_163_266),
	.V (V_163)
);

VNU_6 #(quan_width) VNU164 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_164),
	.C2V_2 (C2V_18_164),
	.C2V_3 (C2V_177_164),
	.C2V_4 (C2V_184_164),
	.C2V_5 (C2V_253_164),
	.C2V_6 (C2V_272_164),
	.L (L_164),
	.V2C_1 (V2C_164_11),
	.V2C_2 (V2C_164_18),
	.V2C_3 (V2C_164_177),
	.V2C_4 (V2C_164_184),
	.V2C_5 (V2C_164_253),
	.V2C_6 (V2C_164_272),
	.V (V_164)
);

VNU_6 #(quan_width) VNU165 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_165),
	.C2V_2 (C2V_24_165),
	.C2V_3 (C2V_183_165),
	.C2V_4 (C2V_190_165),
	.C2V_5 (C2V_259_165),
	.C2V_6 (C2V_278_165),
	.L (L_165),
	.V2C_1 (V2C_165_17),
	.V2C_2 (V2C_165_24),
	.V2C_3 (V2C_165_183),
	.V2C_4 (V2C_165_190),
	.V2C_5 (V2C_165_259),
	.V2C_6 (V2C_165_278),
	.V (V_165)
);

VNU_6 #(quan_width) VNU166 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_166),
	.C2V_2 (C2V_30_166),
	.C2V_3 (C2V_189_166),
	.C2V_4 (C2V_196_166),
	.C2V_5 (C2V_265_166),
	.C2V_6 (C2V_284_166),
	.L (L_166),
	.V2C_1 (V2C_166_23),
	.V2C_2 (V2C_166_30),
	.V2C_3 (V2C_166_189),
	.V2C_4 (V2C_166_196),
	.V2C_5 (V2C_166_265),
	.V2C_6 (V2C_166_284),
	.V (V_166)
);

VNU_6 #(quan_width) VNU167 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_167),
	.C2V_2 (C2V_29_167),
	.C2V_3 (C2V_36_167),
	.C2V_4 (C2V_195_167),
	.C2V_5 (C2V_202_167),
	.C2V_6 (C2V_271_167),
	.L (L_167),
	.V2C_1 (V2C_167_2),
	.V2C_2 (V2C_167_29),
	.V2C_3 (V2C_167_36),
	.V2C_4 (V2C_167_195),
	.V2C_5 (V2C_167_202),
	.V2C_6 (V2C_167_271),
	.V (V_167)
);

VNU_6 #(quan_width) VNU168 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_168),
	.C2V_2 (C2V_35_168),
	.C2V_3 (C2V_42_168),
	.C2V_4 (C2V_201_168),
	.C2V_5 (C2V_208_168),
	.C2V_6 (C2V_277_168),
	.L (L_168),
	.V2C_1 (V2C_168_8),
	.V2C_2 (V2C_168_35),
	.V2C_3 (V2C_168_42),
	.V2C_4 (V2C_168_201),
	.V2C_5 (V2C_168_208),
	.V2C_6 (V2C_168_277),
	.V (V_168)
);

VNU_6 #(quan_width) VNU169 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_169),
	.C2V_2 (C2V_41_169),
	.C2V_3 (C2V_48_169),
	.C2V_4 (C2V_207_169),
	.C2V_5 (C2V_214_169),
	.C2V_6 (C2V_283_169),
	.L (L_169),
	.V2C_1 (V2C_169_14),
	.V2C_2 (V2C_169_41),
	.V2C_3 (V2C_169_48),
	.V2C_4 (V2C_169_207),
	.V2C_5 (V2C_169_214),
	.V2C_6 (V2C_169_283),
	.V (V_169)
);

VNU_6 #(quan_width) VNU170 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_170),
	.C2V_2 (C2V_20_170),
	.C2V_3 (C2V_47_170),
	.C2V_4 (C2V_54_170),
	.C2V_5 (C2V_213_170),
	.C2V_6 (C2V_220_170),
	.L (L_170),
	.V2C_1 (V2C_170_1),
	.V2C_2 (V2C_170_20),
	.V2C_3 (V2C_170_47),
	.V2C_4 (V2C_170_54),
	.V2C_5 (V2C_170_213),
	.V2C_6 (V2C_170_220),
	.V (V_170)
);

VNU_6 #(quan_width) VNU171 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_171),
	.C2V_2 (C2V_26_171),
	.C2V_3 (C2V_53_171),
	.C2V_4 (C2V_60_171),
	.C2V_5 (C2V_219_171),
	.C2V_6 (C2V_226_171),
	.L (L_171),
	.V2C_1 (V2C_171_7),
	.V2C_2 (V2C_171_26),
	.V2C_3 (V2C_171_53),
	.V2C_4 (V2C_171_60),
	.V2C_5 (V2C_171_219),
	.V2C_6 (V2C_171_226),
	.V (V_171)
);

VNU_6 #(quan_width) VNU172 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_172),
	.C2V_2 (C2V_32_172),
	.C2V_3 (C2V_59_172),
	.C2V_4 (C2V_66_172),
	.C2V_5 (C2V_225_172),
	.C2V_6 (C2V_232_172),
	.L (L_172),
	.V2C_1 (V2C_172_13),
	.V2C_2 (V2C_172_32),
	.V2C_3 (V2C_172_59),
	.V2C_4 (V2C_172_66),
	.V2C_5 (V2C_172_225),
	.V2C_6 (V2C_172_232),
	.V (V_172)
);

VNU_6 #(quan_width) VNU173 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_173),
	.C2V_2 (C2V_38_173),
	.C2V_3 (C2V_65_173),
	.C2V_4 (C2V_72_173),
	.C2V_5 (C2V_231_173),
	.C2V_6 (C2V_238_173),
	.L (L_173),
	.V2C_1 (V2C_173_19),
	.V2C_2 (V2C_173_38),
	.V2C_3 (V2C_173_65),
	.V2C_4 (V2C_173_72),
	.V2C_5 (V2C_173_231),
	.V2C_6 (V2C_173_238),
	.V (V_173)
);

VNU_6 #(quan_width) VNU174 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_174),
	.C2V_2 (C2V_44_174),
	.C2V_3 (C2V_71_174),
	.C2V_4 (C2V_78_174),
	.C2V_5 (C2V_237_174),
	.C2V_6 (C2V_244_174),
	.L (L_174),
	.V2C_1 (V2C_174_25),
	.V2C_2 (V2C_174_44),
	.V2C_3 (V2C_174_71),
	.V2C_4 (V2C_174_78),
	.V2C_5 (V2C_174_237),
	.V2C_6 (V2C_174_244),
	.V (V_174)
);

VNU_6 #(quan_width) VNU175 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_175),
	.C2V_2 (C2V_50_175),
	.C2V_3 (C2V_77_175),
	.C2V_4 (C2V_84_175),
	.C2V_5 (C2V_243_175),
	.C2V_6 (C2V_250_175),
	.L (L_175),
	.V2C_1 (V2C_175_31),
	.V2C_2 (V2C_175_50),
	.V2C_3 (V2C_175_77),
	.V2C_4 (V2C_175_84),
	.V2C_5 (V2C_175_243),
	.V2C_6 (V2C_175_250),
	.V (V_175)
);

VNU_6 #(quan_width) VNU176 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_176),
	.C2V_2 (C2V_56_176),
	.C2V_3 (C2V_83_176),
	.C2V_4 (C2V_90_176),
	.C2V_5 (C2V_249_176),
	.C2V_6 (C2V_256_176),
	.L (L_176),
	.V2C_1 (V2C_176_37),
	.V2C_2 (V2C_176_56),
	.V2C_3 (V2C_176_83),
	.V2C_4 (V2C_176_90),
	.V2C_5 (V2C_176_249),
	.V2C_6 (V2C_176_256),
	.V (V_176)
);

VNU_6 #(quan_width) VNU177 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_177),
	.C2V_2 (C2V_62_177),
	.C2V_3 (C2V_89_177),
	.C2V_4 (C2V_96_177),
	.C2V_5 (C2V_255_177),
	.C2V_6 (C2V_262_177),
	.L (L_177),
	.V2C_1 (V2C_177_43),
	.V2C_2 (V2C_177_62),
	.V2C_3 (V2C_177_89),
	.V2C_4 (V2C_177_96),
	.V2C_5 (V2C_177_255),
	.V2C_6 (V2C_177_262),
	.V (V_177)
);

VNU_6 #(quan_width) VNU178 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_178),
	.C2V_2 (C2V_68_178),
	.C2V_3 (C2V_95_178),
	.C2V_4 (C2V_102_178),
	.C2V_5 (C2V_261_178),
	.C2V_6 (C2V_268_178),
	.L (L_178),
	.V2C_1 (V2C_178_49),
	.V2C_2 (V2C_178_68),
	.V2C_3 (V2C_178_95),
	.V2C_4 (V2C_178_102),
	.V2C_5 (V2C_178_261),
	.V2C_6 (V2C_178_268),
	.V (V_178)
);

VNU_6 #(quan_width) VNU179 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_179),
	.C2V_2 (C2V_74_179),
	.C2V_3 (C2V_101_179),
	.C2V_4 (C2V_108_179),
	.C2V_5 (C2V_267_179),
	.C2V_6 (C2V_274_179),
	.L (L_179),
	.V2C_1 (V2C_179_55),
	.V2C_2 (V2C_179_74),
	.V2C_3 (V2C_179_101),
	.V2C_4 (V2C_179_108),
	.V2C_5 (V2C_179_267),
	.V2C_6 (V2C_179_274),
	.V (V_179)
);

VNU_6 #(quan_width) VNU180 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_180),
	.C2V_2 (C2V_80_180),
	.C2V_3 (C2V_107_180),
	.C2V_4 (C2V_114_180),
	.C2V_5 (C2V_273_180),
	.C2V_6 (C2V_280_180),
	.L (L_180),
	.V2C_1 (V2C_180_61),
	.V2C_2 (V2C_180_80),
	.V2C_3 (V2C_180_107),
	.V2C_4 (V2C_180_114),
	.V2C_5 (V2C_180_273),
	.V2C_6 (V2C_180_280),
	.V (V_180)
);

VNU_6 #(quan_width) VNU181 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_181),
	.C2V_2 (C2V_86_181),
	.C2V_3 (C2V_113_181),
	.C2V_4 (C2V_120_181),
	.C2V_5 (C2V_279_181),
	.C2V_6 (C2V_286_181),
	.L (L_181),
	.V2C_1 (V2C_181_67),
	.V2C_2 (V2C_181_86),
	.V2C_3 (V2C_181_113),
	.V2C_4 (V2C_181_120),
	.V2C_5 (V2C_181_279),
	.V2C_6 (V2C_181_286),
	.V (V_181)
);

VNU_6 #(quan_width) VNU182 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_182),
	.C2V_2 (C2V_73_182),
	.C2V_3 (C2V_92_182),
	.C2V_4 (C2V_119_182),
	.C2V_5 (C2V_126_182),
	.C2V_6 (C2V_285_182),
	.L (L_182),
	.V2C_1 (V2C_182_4),
	.V2C_2 (V2C_182_73),
	.V2C_3 (V2C_182_92),
	.V2C_4 (V2C_182_119),
	.V2C_5 (V2C_182_126),
	.V2C_6 (V2C_182_285),
	.V (V_182)
);

VNU_6 #(quan_width) VNU183 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_183),
	.C2V_2 (C2V_10_183),
	.C2V_3 (C2V_79_183),
	.C2V_4 (C2V_98_183),
	.C2V_5 (C2V_125_183),
	.C2V_6 (C2V_132_183),
	.L (L_183),
	.V2C_1 (V2C_183_3),
	.V2C_2 (V2C_183_10),
	.V2C_3 (V2C_183_79),
	.V2C_4 (V2C_183_98),
	.V2C_5 (V2C_183_125),
	.V2C_6 (V2C_183_132),
	.V (V_183)
);

VNU_6 #(quan_width) VNU184 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_184),
	.C2V_2 (C2V_16_184),
	.C2V_3 (C2V_85_184),
	.C2V_4 (C2V_104_184),
	.C2V_5 (C2V_131_184),
	.C2V_6 (C2V_138_184),
	.L (L_184),
	.V2C_1 (V2C_184_9),
	.V2C_2 (V2C_184_16),
	.V2C_3 (V2C_184_85),
	.V2C_4 (V2C_184_104),
	.V2C_5 (V2C_184_131),
	.V2C_6 (V2C_184_138),
	.V (V_184)
);

VNU_6 #(quan_width) VNU185 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_185),
	.C2V_2 (C2V_22_185),
	.C2V_3 (C2V_91_185),
	.C2V_4 (C2V_110_185),
	.C2V_5 (C2V_137_185),
	.C2V_6 (C2V_144_185),
	.L (L_185),
	.V2C_1 (V2C_185_15),
	.V2C_2 (V2C_185_22),
	.V2C_3 (V2C_185_91),
	.V2C_4 (V2C_185_110),
	.V2C_5 (V2C_185_137),
	.V2C_6 (V2C_185_144),
	.V (V_185)
);

VNU_6 #(quan_width) VNU186 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_186),
	.C2V_2 (C2V_28_186),
	.C2V_3 (C2V_97_186),
	.C2V_4 (C2V_116_186),
	.C2V_5 (C2V_143_186),
	.C2V_6 (C2V_150_186),
	.L (L_186),
	.V2C_1 (V2C_186_21),
	.V2C_2 (V2C_186_28),
	.V2C_3 (V2C_186_97),
	.V2C_4 (V2C_186_116),
	.V2C_5 (V2C_186_143),
	.V2C_6 (V2C_186_150),
	.V (V_186)
);

VNU_6 #(quan_width) VNU187 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_187),
	.C2V_2 (C2V_34_187),
	.C2V_3 (C2V_103_187),
	.C2V_4 (C2V_122_187),
	.C2V_5 (C2V_149_187),
	.C2V_6 (C2V_156_187),
	.L (L_187),
	.V2C_1 (V2C_187_27),
	.V2C_2 (V2C_187_34),
	.V2C_3 (V2C_187_103),
	.V2C_4 (V2C_187_122),
	.V2C_5 (V2C_187_149),
	.V2C_6 (V2C_187_156),
	.V (V_187)
);

VNU_6 #(quan_width) VNU188 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_188),
	.C2V_2 (C2V_40_188),
	.C2V_3 (C2V_109_188),
	.C2V_4 (C2V_128_188),
	.C2V_5 (C2V_155_188),
	.C2V_6 (C2V_162_188),
	.L (L_188),
	.V2C_1 (V2C_188_33),
	.V2C_2 (V2C_188_40),
	.V2C_3 (V2C_188_109),
	.V2C_4 (V2C_188_128),
	.V2C_5 (V2C_188_155),
	.V2C_6 (V2C_188_162),
	.V (V_188)
);

VNU_6 #(quan_width) VNU189 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_189),
	.C2V_2 (C2V_46_189),
	.C2V_3 (C2V_115_189),
	.C2V_4 (C2V_134_189),
	.C2V_5 (C2V_161_189),
	.C2V_6 (C2V_168_189),
	.L (L_189),
	.V2C_1 (V2C_189_39),
	.V2C_2 (V2C_189_46),
	.V2C_3 (V2C_189_115),
	.V2C_4 (V2C_189_134),
	.V2C_5 (V2C_189_161),
	.V2C_6 (V2C_189_168),
	.V (V_189)
);

VNU_6 #(quan_width) VNU190 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_190),
	.C2V_2 (C2V_52_190),
	.C2V_3 (C2V_121_190),
	.C2V_4 (C2V_140_190),
	.C2V_5 (C2V_167_190),
	.C2V_6 (C2V_174_190),
	.L (L_190),
	.V2C_1 (V2C_190_45),
	.V2C_2 (V2C_190_52),
	.V2C_3 (V2C_190_121),
	.V2C_4 (V2C_190_140),
	.V2C_5 (V2C_190_167),
	.V2C_6 (V2C_190_174),
	.V (V_190)
);

VNU_6 #(quan_width) VNU191 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_191),
	.C2V_2 (C2V_58_191),
	.C2V_3 (C2V_127_191),
	.C2V_4 (C2V_146_191),
	.C2V_5 (C2V_173_191),
	.C2V_6 (C2V_180_191),
	.L (L_191),
	.V2C_1 (V2C_191_51),
	.V2C_2 (V2C_191_58),
	.V2C_3 (V2C_191_127),
	.V2C_4 (V2C_191_146),
	.V2C_5 (V2C_191_173),
	.V2C_6 (V2C_191_180),
	.V (V_191)
);

VNU_6 #(quan_width) VNU192 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_192),
	.C2V_2 (C2V_64_192),
	.C2V_3 (C2V_133_192),
	.C2V_4 (C2V_152_192),
	.C2V_5 (C2V_179_192),
	.C2V_6 (C2V_186_192),
	.L (L_192),
	.V2C_1 (V2C_192_57),
	.V2C_2 (V2C_192_64),
	.V2C_3 (V2C_192_133),
	.V2C_4 (V2C_192_152),
	.V2C_5 (V2C_192_179),
	.V2C_6 (V2C_192_186),
	.V (V_192)
);

VNU_6 #(quan_width) VNU193 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_193),
	.C2V_2 (C2V_89_193),
	.C2V_3 (C2V_243_193),
	.C2V_4 (C2V_256_193),
	.C2V_5 (C2V_272_193),
	.C2V_6 (C2V_276_193),
	.L (L_193),
	.V2C_1 (V2C_193_55),
	.V2C_2 (V2C_193_89),
	.V2C_3 (V2C_193_243),
	.V2C_4 (V2C_193_256),
	.V2C_5 (V2C_193_272),
	.V2C_6 (V2C_193_276),
	.V (V_193)
);

VNU_6 #(quan_width) VNU194 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_194),
	.C2V_2 (C2V_95_194),
	.C2V_3 (C2V_249_194),
	.C2V_4 (C2V_262_194),
	.C2V_5 (C2V_278_194),
	.C2V_6 (C2V_282_194),
	.L (L_194),
	.V2C_1 (V2C_194_61),
	.V2C_2 (V2C_194_95),
	.V2C_3 (V2C_194_249),
	.V2C_4 (V2C_194_262),
	.V2C_5 (V2C_194_278),
	.V2C_6 (V2C_194_282),
	.V (V_194)
);

VNU_6 #(quan_width) VNU195 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_195),
	.C2V_2 (C2V_101_195),
	.C2V_3 (C2V_255_195),
	.C2V_4 (C2V_268_195),
	.C2V_5 (C2V_284_195),
	.C2V_6 (C2V_288_195),
	.L (L_195),
	.V2C_1 (V2C_195_67),
	.V2C_2 (V2C_195_101),
	.V2C_3 (V2C_195_255),
	.V2C_4 (V2C_195_268),
	.V2C_5 (V2C_195_284),
	.V2C_6 (V2C_195_288),
	.V (V_195)
);

VNU_6 #(quan_width) VNU196 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_196),
	.C2V_2 (C2V_6_196),
	.C2V_3 (C2V_73_196),
	.C2V_4 (C2V_107_196),
	.C2V_5 (C2V_261_196),
	.C2V_6 (C2V_274_196),
	.L (L_196),
	.V2C_1 (V2C_196_2),
	.V2C_2 (V2C_196_6),
	.V2C_3 (V2C_196_73),
	.V2C_4 (V2C_196_107),
	.V2C_5 (V2C_196_261),
	.V2C_6 (V2C_196_274),
	.V (V_196)
);

VNU_6 #(quan_width) VNU197 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_197),
	.C2V_2 (C2V_12_197),
	.C2V_3 (C2V_79_197),
	.C2V_4 (C2V_113_197),
	.C2V_5 (C2V_267_197),
	.C2V_6 (C2V_280_197),
	.L (L_197),
	.V2C_1 (V2C_197_8),
	.V2C_2 (V2C_197_12),
	.V2C_3 (V2C_197_79),
	.V2C_4 (V2C_197_113),
	.V2C_5 (V2C_197_267),
	.V2C_6 (V2C_197_280),
	.V (V_197)
);

VNU_6 #(quan_width) VNU198 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_198),
	.C2V_2 (C2V_18_198),
	.C2V_3 (C2V_85_198),
	.C2V_4 (C2V_119_198),
	.C2V_5 (C2V_273_198),
	.C2V_6 (C2V_286_198),
	.L (L_198),
	.V2C_1 (V2C_198_14),
	.V2C_2 (V2C_198_18),
	.V2C_3 (V2C_198_85),
	.V2C_4 (V2C_198_119),
	.V2C_5 (V2C_198_273),
	.V2C_6 (V2C_198_286),
	.V (V_198)
);

VNU_6 #(quan_width) VNU199 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_199),
	.C2V_2 (C2V_20_199),
	.C2V_3 (C2V_24_199),
	.C2V_4 (C2V_91_199),
	.C2V_5 (C2V_125_199),
	.C2V_6 (C2V_279_199),
	.L (L_199),
	.V2C_1 (V2C_199_4),
	.V2C_2 (V2C_199_20),
	.V2C_3 (V2C_199_24),
	.V2C_4 (V2C_199_91),
	.V2C_5 (V2C_199_125),
	.V2C_6 (V2C_199_279),
	.V (V_199)
);

VNU_6 #(quan_width) VNU200 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_200),
	.C2V_2 (C2V_26_200),
	.C2V_3 (C2V_30_200),
	.C2V_4 (C2V_97_200),
	.C2V_5 (C2V_131_200),
	.C2V_6 (C2V_285_200),
	.L (L_200),
	.V2C_1 (V2C_200_10),
	.V2C_2 (V2C_200_26),
	.V2C_3 (V2C_200_30),
	.V2C_4 (V2C_200_97),
	.V2C_5 (V2C_200_131),
	.V2C_6 (V2C_200_285),
	.V (V_200)
);

VNU_6 #(quan_width) VNU201 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_201),
	.C2V_2 (C2V_16_201),
	.C2V_3 (C2V_32_201),
	.C2V_4 (C2V_36_201),
	.C2V_5 (C2V_103_201),
	.C2V_6 (C2V_137_201),
	.L (L_201),
	.V2C_1 (V2C_201_3),
	.V2C_2 (V2C_201_16),
	.V2C_3 (V2C_201_32),
	.V2C_4 (V2C_201_36),
	.V2C_5 (V2C_201_103),
	.V2C_6 (V2C_201_137),
	.V (V_201)
);

VNU_6 #(quan_width) VNU202 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_202),
	.C2V_2 (C2V_22_202),
	.C2V_3 (C2V_38_202),
	.C2V_4 (C2V_42_202),
	.C2V_5 (C2V_109_202),
	.C2V_6 (C2V_143_202),
	.L (L_202),
	.V2C_1 (V2C_202_9),
	.V2C_2 (V2C_202_22),
	.V2C_3 (V2C_202_38),
	.V2C_4 (V2C_202_42),
	.V2C_5 (V2C_202_109),
	.V2C_6 (V2C_202_143),
	.V (V_202)
);

VNU_6 #(quan_width) VNU203 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_203),
	.C2V_2 (C2V_28_203),
	.C2V_3 (C2V_44_203),
	.C2V_4 (C2V_48_203),
	.C2V_5 (C2V_115_203),
	.C2V_6 (C2V_149_203),
	.L (L_203),
	.V2C_1 (V2C_203_15),
	.V2C_2 (V2C_203_28),
	.V2C_3 (V2C_203_44),
	.V2C_4 (V2C_203_48),
	.V2C_5 (V2C_203_115),
	.V2C_6 (V2C_203_149),
	.V (V_203)
);

VNU_6 #(quan_width) VNU204 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_204),
	.C2V_2 (C2V_34_204),
	.C2V_3 (C2V_50_204),
	.C2V_4 (C2V_54_204),
	.C2V_5 (C2V_121_204),
	.C2V_6 (C2V_155_204),
	.L (L_204),
	.V2C_1 (V2C_204_21),
	.V2C_2 (V2C_204_34),
	.V2C_3 (V2C_204_50),
	.V2C_4 (V2C_204_54),
	.V2C_5 (V2C_204_121),
	.V2C_6 (V2C_204_155),
	.V (V_204)
);

VNU_6 #(quan_width) VNU205 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_205),
	.C2V_2 (C2V_40_205),
	.C2V_3 (C2V_56_205),
	.C2V_4 (C2V_60_205),
	.C2V_5 (C2V_127_205),
	.C2V_6 (C2V_161_205),
	.L (L_205),
	.V2C_1 (V2C_205_27),
	.V2C_2 (V2C_205_40),
	.V2C_3 (V2C_205_56),
	.V2C_4 (V2C_205_60),
	.V2C_5 (V2C_205_127),
	.V2C_6 (V2C_205_161),
	.V (V_205)
);

VNU_6 #(quan_width) VNU206 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_206),
	.C2V_2 (C2V_46_206),
	.C2V_3 (C2V_62_206),
	.C2V_4 (C2V_66_206),
	.C2V_5 (C2V_133_206),
	.C2V_6 (C2V_167_206),
	.L (L_206),
	.V2C_1 (V2C_206_33),
	.V2C_2 (V2C_206_46),
	.V2C_3 (V2C_206_62),
	.V2C_4 (V2C_206_66),
	.V2C_5 (V2C_206_133),
	.V2C_6 (V2C_206_167),
	.V (V_206)
);

VNU_6 #(quan_width) VNU207 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_207),
	.C2V_2 (C2V_52_207),
	.C2V_3 (C2V_68_207),
	.C2V_4 (C2V_72_207),
	.C2V_5 (C2V_139_207),
	.C2V_6 (C2V_173_207),
	.L (L_207),
	.V2C_1 (V2C_207_39),
	.V2C_2 (V2C_207_52),
	.V2C_3 (V2C_207_68),
	.V2C_4 (V2C_207_72),
	.V2C_5 (V2C_207_139),
	.V2C_6 (V2C_207_173),
	.V (V_207)
);

VNU_6 #(quan_width) VNU208 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_208),
	.C2V_2 (C2V_58_208),
	.C2V_3 (C2V_74_208),
	.C2V_4 (C2V_78_208),
	.C2V_5 (C2V_145_208),
	.C2V_6 (C2V_179_208),
	.L (L_208),
	.V2C_1 (V2C_208_45),
	.V2C_2 (V2C_208_58),
	.V2C_3 (V2C_208_74),
	.V2C_4 (V2C_208_78),
	.V2C_5 (V2C_208_145),
	.V2C_6 (V2C_208_179),
	.V (V_208)
);

VNU_6 #(quan_width) VNU209 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_209),
	.C2V_2 (C2V_64_209),
	.C2V_3 (C2V_80_209),
	.C2V_4 (C2V_84_209),
	.C2V_5 (C2V_151_209),
	.C2V_6 (C2V_185_209),
	.L (L_209),
	.V2C_1 (V2C_209_51),
	.V2C_2 (V2C_209_64),
	.V2C_3 (V2C_209_80),
	.V2C_4 (V2C_209_84),
	.V2C_5 (V2C_209_151),
	.V2C_6 (V2C_209_185),
	.V (V_209)
);

VNU_6 #(quan_width) VNU210 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_210),
	.C2V_2 (C2V_70_210),
	.C2V_3 (C2V_86_210),
	.C2V_4 (C2V_90_210),
	.C2V_5 (C2V_157_210),
	.C2V_6 (C2V_191_210),
	.L (L_210),
	.V2C_1 (V2C_210_57),
	.V2C_2 (V2C_210_70),
	.V2C_3 (V2C_210_86),
	.V2C_4 (V2C_210_90),
	.V2C_5 (V2C_210_157),
	.V2C_6 (V2C_210_191),
	.V (V_210)
);

VNU_6 #(quan_width) VNU211 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_211),
	.C2V_2 (C2V_76_211),
	.C2V_3 (C2V_92_211),
	.C2V_4 (C2V_96_211),
	.C2V_5 (C2V_163_211),
	.C2V_6 (C2V_197_211),
	.L (L_211),
	.V2C_1 (V2C_211_63),
	.V2C_2 (V2C_211_76),
	.V2C_3 (V2C_211_92),
	.V2C_4 (V2C_211_96),
	.V2C_5 (V2C_211_163),
	.V2C_6 (V2C_211_197),
	.V (V_211)
);

VNU_6 #(quan_width) VNU212 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_212),
	.C2V_2 (C2V_82_212),
	.C2V_3 (C2V_98_212),
	.C2V_4 (C2V_102_212),
	.C2V_5 (C2V_169_212),
	.C2V_6 (C2V_203_212),
	.L (L_212),
	.V2C_1 (V2C_212_69),
	.V2C_2 (V2C_212_82),
	.V2C_3 (V2C_212_98),
	.V2C_4 (V2C_212_102),
	.V2C_5 (V2C_212_169),
	.V2C_6 (V2C_212_203),
	.V (V_212)
);

VNU_6 #(quan_width) VNU213 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_213),
	.C2V_2 (C2V_88_213),
	.C2V_3 (C2V_104_213),
	.C2V_4 (C2V_108_213),
	.C2V_5 (C2V_175_213),
	.C2V_6 (C2V_209_213),
	.L (L_213),
	.V2C_1 (V2C_213_75),
	.V2C_2 (V2C_213_88),
	.V2C_3 (V2C_213_104),
	.V2C_4 (V2C_213_108),
	.V2C_5 (V2C_213_175),
	.V2C_6 (V2C_213_209),
	.V (V_213)
);

VNU_6 #(quan_width) VNU214 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_214),
	.C2V_2 (C2V_94_214),
	.C2V_3 (C2V_110_214),
	.C2V_4 (C2V_114_214),
	.C2V_5 (C2V_181_214),
	.C2V_6 (C2V_215_214),
	.L (L_214),
	.V2C_1 (V2C_214_81),
	.V2C_2 (V2C_214_94),
	.V2C_3 (V2C_214_110),
	.V2C_4 (V2C_214_114),
	.V2C_5 (V2C_214_181),
	.V2C_6 (V2C_214_215),
	.V (V_214)
);

VNU_6 #(quan_width) VNU215 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_215),
	.C2V_2 (C2V_100_215),
	.C2V_3 (C2V_116_215),
	.C2V_4 (C2V_120_215),
	.C2V_5 (C2V_187_215),
	.C2V_6 (C2V_221_215),
	.L (L_215),
	.V2C_1 (V2C_215_87),
	.V2C_2 (V2C_215_100),
	.V2C_3 (V2C_215_116),
	.V2C_4 (V2C_215_120),
	.V2C_5 (V2C_215_187),
	.V2C_6 (V2C_215_221),
	.V (V_215)
);

VNU_6 #(quan_width) VNU216 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_93_216),
	.C2V_2 (C2V_106_216),
	.C2V_3 (C2V_122_216),
	.C2V_4 (C2V_126_216),
	.C2V_5 (C2V_193_216),
	.C2V_6 (C2V_227_216),
	.L (L_216),
	.V2C_1 (V2C_216_93),
	.V2C_2 (V2C_216_106),
	.V2C_3 (V2C_216_122),
	.V2C_4 (V2C_216_126),
	.V2C_5 (V2C_216_193),
	.V2C_6 (V2C_216_227),
	.V (V_216)
);

VNU_6 #(quan_width) VNU217 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_99_217),
	.C2V_2 (C2V_112_217),
	.C2V_3 (C2V_128_217),
	.C2V_4 (C2V_132_217),
	.C2V_5 (C2V_199_217),
	.C2V_6 (C2V_233_217),
	.L (L_217),
	.V2C_1 (V2C_217_99),
	.V2C_2 (V2C_217_112),
	.V2C_3 (V2C_217_128),
	.V2C_4 (V2C_217_132),
	.V2C_5 (V2C_217_199),
	.V2C_6 (V2C_217_233),
	.V (V_217)
);

VNU_6 #(quan_width) VNU218 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_105_218),
	.C2V_2 (C2V_118_218),
	.C2V_3 (C2V_134_218),
	.C2V_4 (C2V_138_218),
	.C2V_5 (C2V_205_218),
	.C2V_6 (C2V_239_218),
	.L (L_218),
	.V2C_1 (V2C_218_105),
	.V2C_2 (V2C_218_118),
	.V2C_3 (V2C_218_134),
	.V2C_4 (V2C_218_138),
	.V2C_5 (V2C_218_205),
	.V2C_6 (V2C_218_239),
	.V (V_218)
);

VNU_6 #(quan_width) VNU219 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_111_219),
	.C2V_2 (C2V_124_219),
	.C2V_3 (C2V_140_219),
	.C2V_4 (C2V_144_219),
	.C2V_5 (C2V_211_219),
	.C2V_6 (C2V_245_219),
	.L (L_219),
	.V2C_1 (V2C_219_111),
	.V2C_2 (V2C_219_124),
	.V2C_3 (V2C_219_140),
	.V2C_4 (V2C_219_144),
	.V2C_5 (V2C_219_211),
	.V2C_6 (V2C_219_245),
	.V (V_219)
);

VNU_6 #(quan_width) VNU220 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_117_220),
	.C2V_2 (C2V_130_220),
	.C2V_3 (C2V_146_220),
	.C2V_4 (C2V_150_220),
	.C2V_5 (C2V_217_220),
	.C2V_6 (C2V_251_220),
	.L (L_220),
	.V2C_1 (V2C_220_117),
	.V2C_2 (V2C_220_130),
	.V2C_3 (V2C_220_146),
	.V2C_4 (V2C_220_150),
	.V2C_5 (V2C_220_217),
	.V2C_6 (V2C_220_251),
	.V (V_220)
);

VNU_6 #(quan_width) VNU221 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_123_221),
	.C2V_2 (C2V_136_221),
	.C2V_3 (C2V_152_221),
	.C2V_4 (C2V_156_221),
	.C2V_5 (C2V_223_221),
	.C2V_6 (C2V_257_221),
	.L (L_221),
	.V2C_1 (V2C_221_123),
	.V2C_2 (V2C_221_136),
	.V2C_3 (V2C_221_152),
	.V2C_4 (V2C_221_156),
	.V2C_5 (V2C_221_223),
	.V2C_6 (V2C_221_257),
	.V (V_221)
);

VNU_6 #(quan_width) VNU222 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_129_222),
	.C2V_2 (C2V_142_222),
	.C2V_3 (C2V_158_222),
	.C2V_4 (C2V_162_222),
	.C2V_5 (C2V_229_222),
	.C2V_6 (C2V_263_222),
	.L (L_222),
	.V2C_1 (V2C_222_129),
	.V2C_2 (V2C_222_142),
	.V2C_3 (V2C_222_158),
	.V2C_4 (V2C_222_162),
	.V2C_5 (V2C_222_229),
	.V2C_6 (V2C_222_263),
	.V (V_222)
);

VNU_6 #(quan_width) VNU223 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_135_223),
	.C2V_2 (C2V_148_223),
	.C2V_3 (C2V_164_223),
	.C2V_4 (C2V_168_223),
	.C2V_5 (C2V_235_223),
	.C2V_6 (C2V_269_223),
	.L (L_223),
	.V2C_1 (V2C_223_135),
	.V2C_2 (V2C_223_148),
	.V2C_3 (V2C_223_164),
	.V2C_4 (V2C_223_168),
	.V2C_5 (V2C_223_235),
	.V2C_6 (V2C_223_269),
	.V (V_223)
);

VNU_6 #(quan_width) VNU224 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_141_224),
	.C2V_2 (C2V_154_224),
	.C2V_3 (C2V_170_224),
	.C2V_4 (C2V_174_224),
	.C2V_5 (C2V_241_224),
	.C2V_6 (C2V_275_224),
	.L (L_224),
	.V2C_1 (V2C_224_141),
	.V2C_2 (V2C_224_154),
	.V2C_3 (V2C_224_170),
	.V2C_4 (V2C_224_174),
	.V2C_5 (V2C_224_241),
	.V2C_6 (V2C_224_275),
	.V (V_224)
);

VNU_6 #(quan_width) VNU225 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_147_225),
	.C2V_2 (C2V_160_225),
	.C2V_3 (C2V_176_225),
	.C2V_4 (C2V_180_225),
	.C2V_5 (C2V_247_225),
	.C2V_6 (C2V_281_225),
	.L (L_225),
	.V2C_1 (V2C_225_147),
	.V2C_2 (V2C_225_160),
	.V2C_3 (V2C_225_176),
	.V2C_4 (V2C_225_180),
	.V2C_5 (V2C_225_247),
	.V2C_6 (V2C_225_281),
	.V (V_225)
);

VNU_6 #(quan_width) VNU226 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_153_226),
	.C2V_2 (C2V_166_226),
	.C2V_3 (C2V_182_226),
	.C2V_4 (C2V_186_226),
	.C2V_5 (C2V_253_226),
	.C2V_6 (C2V_287_226),
	.L (L_226),
	.V2C_1 (V2C_226_153),
	.V2C_2 (V2C_226_166),
	.V2C_3 (V2C_226_182),
	.V2C_4 (V2C_226_186),
	.V2C_5 (V2C_226_253),
	.V2C_6 (V2C_226_287),
	.V (V_226)
);

VNU_6 #(quan_width) VNU227 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_227),
	.C2V_2 (C2V_159_227),
	.C2V_3 (C2V_172_227),
	.C2V_4 (C2V_188_227),
	.C2V_5 (C2V_192_227),
	.C2V_6 (C2V_259_227),
	.L (L_227),
	.V2C_1 (V2C_227_5),
	.V2C_2 (V2C_227_159),
	.V2C_3 (V2C_227_172),
	.V2C_4 (V2C_227_188),
	.V2C_5 (V2C_227_192),
	.V2C_6 (V2C_227_259),
	.V (V_227)
);

VNU_6 #(quan_width) VNU228 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_228),
	.C2V_2 (C2V_165_228),
	.C2V_3 (C2V_178_228),
	.C2V_4 (C2V_194_228),
	.C2V_5 (C2V_198_228),
	.C2V_6 (C2V_265_228),
	.L (L_228),
	.V2C_1 (V2C_228_11),
	.V2C_2 (V2C_228_165),
	.V2C_3 (V2C_228_178),
	.V2C_4 (V2C_228_194),
	.V2C_5 (V2C_228_198),
	.V2C_6 (V2C_228_265),
	.V (V_228)
);

VNU_6 #(quan_width) VNU229 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_229),
	.C2V_2 (C2V_171_229),
	.C2V_3 (C2V_184_229),
	.C2V_4 (C2V_200_229),
	.C2V_5 (C2V_204_229),
	.C2V_6 (C2V_271_229),
	.L (L_229),
	.V2C_1 (V2C_229_17),
	.V2C_2 (V2C_229_171),
	.V2C_3 (V2C_229_184),
	.V2C_4 (V2C_229_200),
	.V2C_5 (V2C_229_204),
	.V2C_6 (V2C_229_271),
	.V (V_229)
);

VNU_6 #(quan_width) VNU230 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_230),
	.C2V_2 (C2V_177_230),
	.C2V_3 (C2V_190_230),
	.C2V_4 (C2V_206_230),
	.C2V_5 (C2V_210_230),
	.C2V_6 (C2V_277_230),
	.L (L_230),
	.V2C_1 (V2C_230_23),
	.V2C_2 (V2C_230_177),
	.V2C_3 (V2C_230_190),
	.V2C_4 (V2C_230_206),
	.V2C_5 (V2C_230_210),
	.V2C_6 (V2C_230_277),
	.V (V_230)
);

VNU_6 #(quan_width) VNU231 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_231),
	.C2V_2 (C2V_183_231),
	.C2V_3 (C2V_196_231),
	.C2V_4 (C2V_212_231),
	.C2V_5 (C2V_216_231),
	.C2V_6 (C2V_283_231),
	.L (L_231),
	.V2C_1 (V2C_231_29),
	.V2C_2 (V2C_231_183),
	.V2C_3 (V2C_231_196),
	.V2C_4 (V2C_231_212),
	.V2C_5 (V2C_231_216),
	.V2C_6 (V2C_231_283),
	.V (V_231)
);

VNU_6 #(quan_width) VNU232 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_232),
	.C2V_2 (C2V_35_232),
	.C2V_3 (C2V_189_232),
	.C2V_4 (C2V_202_232),
	.C2V_5 (C2V_218_232),
	.C2V_6 (C2V_222_232),
	.L (L_232),
	.V2C_1 (V2C_232_1),
	.V2C_2 (V2C_232_35),
	.V2C_3 (V2C_232_189),
	.V2C_4 (V2C_232_202),
	.V2C_5 (V2C_232_218),
	.V2C_6 (V2C_232_222),
	.V (V_232)
);

VNU_6 #(quan_width) VNU233 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_233),
	.C2V_2 (C2V_41_233),
	.C2V_3 (C2V_195_233),
	.C2V_4 (C2V_208_233),
	.C2V_5 (C2V_224_233),
	.C2V_6 (C2V_228_233),
	.L (L_233),
	.V2C_1 (V2C_233_7),
	.V2C_2 (V2C_233_41),
	.V2C_3 (V2C_233_195),
	.V2C_4 (V2C_233_208),
	.V2C_5 (V2C_233_224),
	.V2C_6 (V2C_233_228),
	.V (V_233)
);

VNU_6 #(quan_width) VNU234 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_234),
	.C2V_2 (C2V_47_234),
	.C2V_3 (C2V_201_234),
	.C2V_4 (C2V_214_234),
	.C2V_5 (C2V_230_234),
	.C2V_6 (C2V_234_234),
	.L (L_234),
	.V2C_1 (V2C_234_13),
	.V2C_2 (V2C_234_47),
	.V2C_3 (V2C_234_201),
	.V2C_4 (V2C_234_214),
	.V2C_5 (V2C_234_230),
	.V2C_6 (V2C_234_234),
	.V (V_234)
);

VNU_6 #(quan_width) VNU235 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_235),
	.C2V_2 (C2V_53_235),
	.C2V_3 (C2V_207_235),
	.C2V_4 (C2V_220_235),
	.C2V_5 (C2V_236_235),
	.C2V_6 (C2V_240_235),
	.L (L_235),
	.V2C_1 (V2C_235_19),
	.V2C_2 (V2C_235_53),
	.V2C_3 (V2C_235_207),
	.V2C_4 (V2C_235_220),
	.V2C_5 (V2C_235_236),
	.V2C_6 (V2C_235_240),
	.V (V_235)
);

VNU_6 #(quan_width) VNU236 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_236),
	.C2V_2 (C2V_59_236),
	.C2V_3 (C2V_213_236),
	.C2V_4 (C2V_226_236),
	.C2V_5 (C2V_242_236),
	.C2V_6 (C2V_246_236),
	.L (L_236),
	.V2C_1 (V2C_236_25),
	.V2C_2 (V2C_236_59),
	.V2C_3 (V2C_236_213),
	.V2C_4 (V2C_236_226),
	.V2C_5 (V2C_236_242),
	.V2C_6 (V2C_236_246),
	.V (V_236)
);

VNU_6 #(quan_width) VNU237 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_237),
	.C2V_2 (C2V_65_237),
	.C2V_3 (C2V_219_237),
	.C2V_4 (C2V_232_237),
	.C2V_5 (C2V_248_237),
	.C2V_6 (C2V_252_237),
	.L (L_237),
	.V2C_1 (V2C_237_31),
	.V2C_2 (V2C_237_65),
	.V2C_3 (V2C_237_219),
	.V2C_4 (V2C_237_232),
	.V2C_5 (V2C_237_248),
	.V2C_6 (V2C_237_252),
	.V (V_237)
);

VNU_6 #(quan_width) VNU238 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_238),
	.C2V_2 (C2V_71_238),
	.C2V_3 (C2V_225_238),
	.C2V_4 (C2V_238_238),
	.C2V_5 (C2V_254_238),
	.C2V_6 (C2V_258_238),
	.L (L_238),
	.V2C_1 (V2C_238_37),
	.V2C_2 (V2C_238_71),
	.V2C_3 (V2C_238_225),
	.V2C_4 (V2C_238_238),
	.V2C_5 (V2C_238_254),
	.V2C_6 (V2C_238_258),
	.V (V_238)
);

VNU_6 #(quan_width) VNU239 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_239),
	.C2V_2 (C2V_77_239),
	.C2V_3 (C2V_231_239),
	.C2V_4 (C2V_244_239),
	.C2V_5 (C2V_260_239),
	.C2V_6 (C2V_264_239),
	.L (L_239),
	.V2C_1 (V2C_239_43),
	.V2C_2 (V2C_239_77),
	.V2C_3 (V2C_239_231),
	.V2C_4 (V2C_239_244),
	.V2C_5 (V2C_239_260),
	.V2C_6 (V2C_239_264),
	.V (V_239)
);

VNU_6 #(quan_width) VNU240 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_240),
	.C2V_2 (C2V_83_240),
	.C2V_3 (C2V_237_240),
	.C2V_4 (C2V_250_240),
	.C2V_5 (C2V_266_240),
	.C2V_6 (C2V_270_240),
	.L (L_240),
	.V2C_1 (V2C_240_49),
	.V2C_2 (V2C_240_83),
	.V2C_3 (V2C_240_237),
	.V2C_4 (V2C_240_250),
	.V2C_5 (V2C_240_266),
	.V2C_6 (V2C_240_270),
	.V (V_240)
);

VNU_6 #(quan_width) VNU241 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_241),
	.C2V_2 (C2V_90_241),
	.C2V_3 (C2V_129_241),
	.C2V_4 (C2V_146_241),
	.C2V_5 (C2V_220_241),
	.C2V_6 (C2V_269_241),
	.L (L_241),
	.V2C_1 (V2C_241_85),
	.V2C_2 (V2C_241_90),
	.V2C_3 (V2C_241_129),
	.V2C_4 (V2C_241_146),
	.V2C_5 (V2C_241_220),
	.V2C_6 (V2C_241_269),
	.V (V_241)
);

VNU_6 #(quan_width) VNU242 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_91_242),
	.C2V_2 (C2V_96_242),
	.C2V_3 (C2V_135_242),
	.C2V_4 (C2V_152_242),
	.C2V_5 (C2V_226_242),
	.C2V_6 (C2V_275_242),
	.L (L_242),
	.V2C_1 (V2C_242_91),
	.V2C_2 (V2C_242_96),
	.V2C_3 (V2C_242_135),
	.V2C_4 (V2C_242_152),
	.V2C_5 (V2C_242_226),
	.V2C_6 (V2C_242_275),
	.V (V_242)
);

VNU_6 #(quan_width) VNU243 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_97_243),
	.C2V_2 (C2V_102_243),
	.C2V_3 (C2V_141_243),
	.C2V_4 (C2V_158_243),
	.C2V_5 (C2V_232_243),
	.C2V_6 (C2V_281_243),
	.L (L_243),
	.V2C_1 (V2C_243_97),
	.V2C_2 (V2C_243_102),
	.V2C_3 (V2C_243_141),
	.V2C_4 (V2C_243_158),
	.V2C_5 (V2C_243_232),
	.V2C_6 (V2C_243_281),
	.V (V_243)
);

VNU_6 #(quan_width) VNU244 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_103_244),
	.C2V_2 (C2V_108_244),
	.C2V_3 (C2V_147_244),
	.C2V_4 (C2V_164_244),
	.C2V_5 (C2V_238_244),
	.C2V_6 (C2V_287_244),
	.L (L_244),
	.V2C_1 (V2C_244_103),
	.V2C_2 (V2C_244_108),
	.V2C_3 (V2C_244_147),
	.V2C_4 (V2C_244_164),
	.V2C_5 (V2C_244_238),
	.V2C_6 (V2C_244_287),
	.V (V_244)
);

VNU_6 #(quan_width) VNU245 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_245),
	.C2V_2 (C2V_109_245),
	.C2V_3 (C2V_114_245),
	.C2V_4 (C2V_153_245),
	.C2V_5 (C2V_170_245),
	.C2V_6 (C2V_244_245),
	.L (L_245),
	.V2C_1 (V2C_245_5),
	.V2C_2 (V2C_245_109),
	.V2C_3 (V2C_245_114),
	.V2C_4 (V2C_245_153),
	.V2C_5 (V2C_245_170),
	.V2C_6 (V2C_245_244),
	.V (V_245)
);

VNU_6 #(quan_width) VNU246 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_246),
	.C2V_2 (C2V_115_246),
	.C2V_3 (C2V_120_246),
	.C2V_4 (C2V_159_246),
	.C2V_5 (C2V_176_246),
	.C2V_6 (C2V_250_246),
	.L (L_246),
	.V2C_1 (V2C_246_11),
	.V2C_2 (V2C_246_115),
	.V2C_3 (V2C_246_120),
	.V2C_4 (V2C_246_159),
	.V2C_5 (V2C_246_176),
	.V2C_6 (V2C_246_250),
	.V (V_246)
);

VNU_6 #(quan_width) VNU247 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_247),
	.C2V_2 (C2V_121_247),
	.C2V_3 (C2V_126_247),
	.C2V_4 (C2V_165_247),
	.C2V_5 (C2V_182_247),
	.C2V_6 (C2V_256_247),
	.L (L_247),
	.V2C_1 (V2C_247_17),
	.V2C_2 (V2C_247_121),
	.V2C_3 (V2C_247_126),
	.V2C_4 (V2C_247_165),
	.V2C_5 (V2C_247_182),
	.V2C_6 (V2C_247_256),
	.V (V_247)
);

VNU_6 #(quan_width) VNU248 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_248),
	.C2V_2 (C2V_127_248),
	.C2V_3 (C2V_132_248),
	.C2V_4 (C2V_171_248),
	.C2V_5 (C2V_188_248),
	.C2V_6 (C2V_262_248),
	.L (L_248),
	.V2C_1 (V2C_248_23),
	.V2C_2 (V2C_248_127),
	.V2C_3 (V2C_248_132),
	.V2C_4 (V2C_248_171),
	.V2C_5 (V2C_248_188),
	.V2C_6 (V2C_248_262),
	.V (V_248)
);

VNU_6 #(quan_width) VNU249 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_249),
	.C2V_2 (C2V_133_249),
	.C2V_3 (C2V_138_249),
	.C2V_4 (C2V_177_249),
	.C2V_5 (C2V_194_249),
	.C2V_6 (C2V_268_249),
	.L (L_249),
	.V2C_1 (V2C_249_29),
	.V2C_2 (V2C_249_133),
	.V2C_3 (V2C_249_138),
	.V2C_4 (V2C_249_177),
	.V2C_5 (V2C_249_194),
	.V2C_6 (V2C_249_268),
	.V (V_249)
);

VNU_6 #(quan_width) VNU250 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_250),
	.C2V_2 (C2V_139_250),
	.C2V_3 (C2V_144_250),
	.C2V_4 (C2V_183_250),
	.C2V_5 (C2V_200_250),
	.C2V_6 (C2V_274_250),
	.L (L_250),
	.V2C_1 (V2C_250_35),
	.V2C_2 (V2C_250_139),
	.V2C_3 (V2C_250_144),
	.V2C_4 (V2C_250_183),
	.V2C_5 (V2C_250_200),
	.V2C_6 (V2C_250_274),
	.V (V_250)
);

VNU_6 #(quan_width) VNU251 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_251),
	.C2V_2 (C2V_145_251),
	.C2V_3 (C2V_150_251),
	.C2V_4 (C2V_189_251),
	.C2V_5 (C2V_206_251),
	.C2V_6 (C2V_280_251),
	.L (L_251),
	.V2C_1 (V2C_251_41),
	.V2C_2 (V2C_251_145),
	.V2C_3 (V2C_251_150),
	.V2C_4 (V2C_251_189),
	.V2C_5 (V2C_251_206),
	.V2C_6 (V2C_251_280),
	.V (V_251)
);

VNU_6 #(quan_width) VNU252 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_252),
	.C2V_2 (C2V_151_252),
	.C2V_3 (C2V_156_252),
	.C2V_4 (C2V_195_252),
	.C2V_5 (C2V_212_252),
	.C2V_6 (C2V_286_252),
	.L (L_252),
	.V2C_1 (V2C_252_47),
	.V2C_2 (V2C_252_151),
	.V2C_3 (V2C_252_156),
	.V2C_4 (V2C_252_195),
	.V2C_5 (V2C_252_212),
	.V2C_6 (V2C_252_286),
	.V (V_252)
);

VNU_6 #(quan_width) VNU253 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_253),
	.C2V_2 (C2V_53_253),
	.C2V_3 (C2V_157_253),
	.C2V_4 (C2V_162_253),
	.C2V_5 (C2V_201_253),
	.C2V_6 (C2V_218_253),
	.L (L_253),
	.V2C_1 (V2C_253_4),
	.V2C_2 (V2C_253_53),
	.V2C_3 (V2C_253_157),
	.V2C_4 (V2C_253_162),
	.V2C_5 (V2C_253_201),
	.V2C_6 (V2C_253_218),
	.V (V_253)
);

VNU_6 #(quan_width) VNU254 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_254),
	.C2V_2 (C2V_59_254),
	.C2V_3 (C2V_163_254),
	.C2V_4 (C2V_168_254),
	.C2V_5 (C2V_207_254),
	.C2V_6 (C2V_224_254),
	.L (L_254),
	.V2C_1 (V2C_254_10),
	.V2C_2 (V2C_254_59),
	.V2C_3 (V2C_254_163),
	.V2C_4 (V2C_254_168),
	.V2C_5 (V2C_254_207),
	.V2C_6 (V2C_254_224),
	.V (V_254)
);

VNU_6 #(quan_width) VNU255 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_255),
	.C2V_2 (C2V_65_255),
	.C2V_3 (C2V_169_255),
	.C2V_4 (C2V_174_255),
	.C2V_5 (C2V_213_255),
	.C2V_6 (C2V_230_255),
	.L (L_255),
	.V2C_1 (V2C_255_16),
	.V2C_2 (V2C_255_65),
	.V2C_3 (V2C_255_169),
	.V2C_4 (V2C_255_174),
	.V2C_5 (V2C_255_213),
	.V2C_6 (V2C_255_230),
	.V (V_255)
);

VNU_6 #(quan_width) VNU256 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_256),
	.C2V_2 (C2V_71_256),
	.C2V_3 (C2V_175_256),
	.C2V_4 (C2V_180_256),
	.C2V_5 (C2V_219_256),
	.C2V_6 (C2V_236_256),
	.L (L_256),
	.V2C_1 (V2C_256_22),
	.V2C_2 (V2C_256_71),
	.V2C_3 (V2C_256_175),
	.V2C_4 (V2C_256_180),
	.V2C_5 (V2C_256_219),
	.V2C_6 (V2C_256_236),
	.V (V_256)
);

VNU_6 #(quan_width) VNU257 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_257),
	.C2V_2 (C2V_77_257),
	.C2V_3 (C2V_181_257),
	.C2V_4 (C2V_186_257),
	.C2V_5 (C2V_225_257),
	.C2V_6 (C2V_242_257),
	.L (L_257),
	.V2C_1 (V2C_257_28),
	.V2C_2 (V2C_257_77),
	.V2C_3 (V2C_257_181),
	.V2C_4 (V2C_257_186),
	.V2C_5 (V2C_257_225),
	.V2C_6 (V2C_257_242),
	.V (V_257)
);

VNU_6 #(quan_width) VNU258 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_258),
	.C2V_2 (C2V_83_258),
	.C2V_3 (C2V_187_258),
	.C2V_4 (C2V_192_258),
	.C2V_5 (C2V_231_258),
	.C2V_6 (C2V_248_258),
	.L (L_258),
	.V2C_1 (V2C_258_34),
	.V2C_2 (V2C_258_83),
	.V2C_3 (V2C_258_187),
	.V2C_4 (V2C_258_192),
	.V2C_5 (V2C_258_231),
	.V2C_6 (V2C_258_248),
	.V (V_258)
);

VNU_6 #(quan_width) VNU259 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_259),
	.C2V_2 (C2V_89_259),
	.C2V_3 (C2V_193_259),
	.C2V_4 (C2V_198_259),
	.C2V_5 (C2V_237_259),
	.C2V_6 (C2V_254_259),
	.L (L_259),
	.V2C_1 (V2C_259_40),
	.V2C_2 (V2C_259_89),
	.V2C_3 (V2C_259_193),
	.V2C_4 (V2C_259_198),
	.V2C_5 (V2C_259_237),
	.V2C_6 (V2C_259_254),
	.V (V_259)
);

VNU_6 #(quan_width) VNU260 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_260),
	.C2V_2 (C2V_95_260),
	.C2V_3 (C2V_199_260),
	.C2V_4 (C2V_204_260),
	.C2V_5 (C2V_243_260),
	.C2V_6 (C2V_260_260),
	.L (L_260),
	.V2C_1 (V2C_260_46),
	.V2C_2 (V2C_260_95),
	.V2C_3 (V2C_260_199),
	.V2C_4 (V2C_260_204),
	.V2C_5 (V2C_260_243),
	.V2C_6 (V2C_260_260),
	.V (V_260)
);

VNU_6 #(quan_width) VNU261 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_261),
	.C2V_2 (C2V_101_261),
	.C2V_3 (C2V_205_261),
	.C2V_4 (C2V_210_261),
	.C2V_5 (C2V_249_261),
	.C2V_6 (C2V_266_261),
	.L (L_261),
	.V2C_1 (V2C_261_52),
	.V2C_2 (V2C_261_101),
	.V2C_3 (V2C_261_205),
	.V2C_4 (V2C_261_210),
	.V2C_5 (V2C_261_249),
	.V2C_6 (V2C_261_266),
	.V (V_261)
);

VNU_6 #(quan_width) VNU262 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_262),
	.C2V_2 (C2V_107_262),
	.C2V_3 (C2V_211_262),
	.C2V_4 (C2V_216_262),
	.C2V_5 (C2V_255_262),
	.C2V_6 (C2V_272_262),
	.L (L_262),
	.V2C_1 (V2C_262_58),
	.V2C_2 (V2C_262_107),
	.V2C_3 (V2C_262_211),
	.V2C_4 (V2C_262_216),
	.V2C_5 (V2C_262_255),
	.V2C_6 (V2C_262_272),
	.V (V_262)
);

VNU_6 #(quan_width) VNU263 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_263),
	.C2V_2 (C2V_113_263),
	.C2V_3 (C2V_217_263),
	.C2V_4 (C2V_222_263),
	.C2V_5 (C2V_261_263),
	.C2V_6 (C2V_278_263),
	.L (L_263),
	.V2C_1 (V2C_263_64),
	.V2C_2 (V2C_263_113),
	.V2C_3 (V2C_263_217),
	.V2C_4 (V2C_263_222),
	.V2C_5 (V2C_263_261),
	.V2C_6 (V2C_263_278),
	.V (V_263)
);

VNU_6 #(quan_width) VNU264 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_264),
	.C2V_2 (C2V_119_264),
	.C2V_3 (C2V_223_264),
	.C2V_4 (C2V_228_264),
	.C2V_5 (C2V_267_264),
	.C2V_6 (C2V_284_264),
	.L (L_264),
	.V2C_1 (V2C_264_70),
	.V2C_2 (V2C_264_119),
	.V2C_3 (V2C_264_223),
	.V2C_4 (V2C_264_228),
	.V2C_5 (V2C_264_267),
	.V2C_6 (V2C_264_284),
	.V (V_264)
);

VNU_6 #(quan_width) VNU265 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_265),
	.C2V_2 (C2V_76_265),
	.C2V_3 (C2V_125_265),
	.C2V_4 (C2V_229_265),
	.C2V_5 (C2V_234_265),
	.C2V_6 (C2V_273_265),
	.L (L_265),
	.V2C_1 (V2C_265_2),
	.V2C_2 (V2C_265_76),
	.V2C_3 (V2C_265_125),
	.V2C_4 (V2C_265_229),
	.V2C_5 (V2C_265_234),
	.V2C_6 (V2C_265_273),
	.V (V_265)
);

VNU_6 #(quan_width) VNU266 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_266),
	.C2V_2 (C2V_82_266),
	.C2V_3 (C2V_131_266),
	.C2V_4 (C2V_235_266),
	.C2V_5 (C2V_240_266),
	.C2V_6 (C2V_279_266),
	.L (L_266),
	.V2C_1 (V2C_266_8),
	.V2C_2 (V2C_266_82),
	.V2C_3 (V2C_266_131),
	.V2C_4 (V2C_266_235),
	.V2C_5 (V2C_266_240),
	.V2C_6 (V2C_266_279),
	.V (V_266)
);

VNU_6 #(quan_width) VNU267 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_267),
	.C2V_2 (C2V_88_267),
	.C2V_3 (C2V_137_267),
	.C2V_4 (C2V_241_267),
	.C2V_5 (C2V_246_267),
	.C2V_6 (C2V_285_267),
	.L (L_267),
	.V2C_1 (V2C_267_14),
	.V2C_2 (V2C_267_88),
	.V2C_3 (V2C_267_137),
	.V2C_4 (V2C_267_241),
	.V2C_5 (V2C_267_246),
	.V2C_6 (V2C_267_285),
	.V (V_267)
);

VNU_6 #(quan_width) VNU268 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_268),
	.C2V_2 (C2V_20_268),
	.C2V_3 (C2V_94_268),
	.C2V_4 (C2V_143_268),
	.C2V_5 (C2V_247_268),
	.C2V_6 (C2V_252_268),
	.L (L_268),
	.V2C_1 (V2C_268_3),
	.V2C_2 (V2C_268_20),
	.V2C_3 (V2C_268_94),
	.V2C_4 (V2C_268_143),
	.V2C_5 (V2C_268_247),
	.V2C_6 (V2C_268_252),
	.V (V_268)
);

VNU_6 #(quan_width) VNU269 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_269),
	.C2V_2 (C2V_26_269),
	.C2V_3 (C2V_100_269),
	.C2V_4 (C2V_149_269),
	.C2V_5 (C2V_253_269),
	.C2V_6 (C2V_258_269),
	.L (L_269),
	.V2C_1 (V2C_269_9),
	.V2C_2 (V2C_269_26),
	.V2C_3 (V2C_269_100),
	.V2C_4 (V2C_269_149),
	.V2C_5 (V2C_269_253),
	.V2C_6 (V2C_269_258),
	.V (V_269)
);

VNU_6 #(quan_width) VNU270 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_270),
	.C2V_2 (C2V_32_270),
	.C2V_3 (C2V_106_270),
	.C2V_4 (C2V_155_270),
	.C2V_5 (C2V_259_270),
	.C2V_6 (C2V_264_270),
	.L (L_270),
	.V2C_1 (V2C_270_15),
	.V2C_2 (V2C_270_32),
	.V2C_3 (V2C_270_106),
	.V2C_4 (V2C_270_155),
	.V2C_5 (V2C_270_259),
	.V2C_6 (V2C_270_264),
	.V (V_270)
);

VNU_6 #(quan_width) VNU271 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_271),
	.C2V_2 (C2V_38_271),
	.C2V_3 (C2V_112_271),
	.C2V_4 (C2V_161_271),
	.C2V_5 (C2V_265_271),
	.C2V_6 (C2V_270_271),
	.L (L_271),
	.V2C_1 (V2C_271_21),
	.V2C_2 (V2C_271_38),
	.V2C_3 (V2C_271_112),
	.V2C_4 (V2C_271_161),
	.V2C_5 (V2C_271_265),
	.V2C_6 (V2C_271_270),
	.V (V_271)
);

VNU_6 #(quan_width) VNU272 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_272),
	.C2V_2 (C2V_44_272),
	.C2V_3 (C2V_118_272),
	.C2V_4 (C2V_167_272),
	.C2V_5 (C2V_271_272),
	.C2V_6 (C2V_276_272),
	.L (L_272),
	.V2C_1 (V2C_272_27),
	.V2C_2 (V2C_272_44),
	.V2C_3 (V2C_272_118),
	.V2C_4 (V2C_272_167),
	.V2C_5 (V2C_272_271),
	.V2C_6 (V2C_272_276),
	.V (V_272)
);

VNU_6 #(quan_width) VNU273 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_273),
	.C2V_2 (C2V_50_273),
	.C2V_3 (C2V_124_273),
	.C2V_4 (C2V_173_273),
	.C2V_5 (C2V_277_273),
	.C2V_6 (C2V_282_273),
	.L (L_273),
	.V2C_1 (V2C_273_33),
	.V2C_2 (V2C_273_50),
	.V2C_3 (V2C_273_124),
	.V2C_4 (V2C_273_173),
	.V2C_5 (V2C_273_277),
	.V2C_6 (V2C_273_282),
	.V (V_273)
);

VNU_6 #(quan_width) VNU274 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_274),
	.C2V_2 (C2V_56_274),
	.C2V_3 (C2V_130_274),
	.C2V_4 (C2V_179_274),
	.C2V_5 (C2V_283_274),
	.C2V_6 (C2V_288_274),
	.L (L_274),
	.V2C_1 (V2C_274_39),
	.V2C_2 (V2C_274_56),
	.V2C_3 (V2C_274_130),
	.V2C_4 (V2C_274_179),
	.V2C_5 (V2C_274_283),
	.V2C_6 (V2C_274_288),
	.V (V_274)
);

VNU_6 #(quan_width) VNU275 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_275),
	.C2V_2 (C2V_6_275),
	.C2V_3 (C2V_45_275),
	.C2V_4 (C2V_62_275),
	.C2V_5 (C2V_136_275),
	.C2V_6 (C2V_185_275),
	.L (L_275),
	.V2C_1 (V2C_275_1),
	.V2C_2 (V2C_275_6),
	.V2C_3 (V2C_275_45),
	.V2C_4 (V2C_275_62),
	.V2C_5 (V2C_275_136),
	.V2C_6 (V2C_275_185),
	.V (V_275)
);

VNU_6 #(quan_width) VNU276 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_276),
	.C2V_2 (C2V_12_276),
	.C2V_3 (C2V_51_276),
	.C2V_4 (C2V_68_276),
	.C2V_5 (C2V_142_276),
	.C2V_6 (C2V_191_276),
	.L (L_276),
	.V2C_1 (V2C_276_7),
	.V2C_2 (V2C_276_12),
	.V2C_3 (V2C_276_51),
	.V2C_4 (V2C_276_68),
	.V2C_5 (V2C_276_142),
	.V2C_6 (V2C_276_191),
	.V (V_276)
);

VNU_6 #(quan_width) VNU277 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_277),
	.C2V_2 (C2V_18_277),
	.C2V_3 (C2V_57_277),
	.C2V_4 (C2V_74_277),
	.C2V_5 (C2V_148_277),
	.C2V_6 (C2V_197_277),
	.L (L_277),
	.V2C_1 (V2C_277_13),
	.V2C_2 (V2C_277_18),
	.V2C_3 (V2C_277_57),
	.V2C_4 (V2C_277_74),
	.V2C_5 (V2C_277_148),
	.V2C_6 (V2C_277_197),
	.V (V_277)
);

VNU_6 #(quan_width) VNU278 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_278),
	.C2V_2 (C2V_24_278),
	.C2V_3 (C2V_63_278),
	.C2V_4 (C2V_80_278),
	.C2V_5 (C2V_154_278),
	.C2V_6 (C2V_203_278),
	.L (L_278),
	.V2C_1 (V2C_278_19),
	.V2C_2 (V2C_278_24),
	.V2C_3 (V2C_278_63),
	.V2C_4 (V2C_278_80),
	.V2C_5 (V2C_278_154),
	.V2C_6 (V2C_278_203),
	.V (V_278)
);

VNU_6 #(quan_width) VNU279 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_279),
	.C2V_2 (C2V_30_279),
	.C2V_3 (C2V_69_279),
	.C2V_4 (C2V_86_279),
	.C2V_5 (C2V_160_279),
	.C2V_6 (C2V_209_279),
	.L (L_279),
	.V2C_1 (V2C_279_25),
	.V2C_2 (V2C_279_30),
	.V2C_3 (V2C_279_69),
	.V2C_4 (V2C_279_86),
	.V2C_5 (V2C_279_160),
	.V2C_6 (V2C_279_209),
	.V (V_279)
);

VNU_6 #(quan_width) VNU280 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_280),
	.C2V_2 (C2V_36_280),
	.C2V_3 (C2V_75_280),
	.C2V_4 (C2V_92_280),
	.C2V_5 (C2V_166_280),
	.C2V_6 (C2V_215_280),
	.L (L_280),
	.V2C_1 (V2C_280_31),
	.V2C_2 (V2C_280_36),
	.V2C_3 (V2C_280_75),
	.V2C_4 (V2C_280_92),
	.V2C_5 (V2C_280_166),
	.V2C_6 (V2C_280_215),
	.V (V_280)
);

VNU_6 #(quan_width) VNU281 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_281),
	.C2V_2 (C2V_42_281),
	.C2V_3 (C2V_81_281),
	.C2V_4 (C2V_98_281),
	.C2V_5 (C2V_172_281),
	.C2V_6 (C2V_221_281),
	.L (L_281),
	.V2C_1 (V2C_281_37),
	.V2C_2 (V2C_281_42),
	.V2C_3 (V2C_281_81),
	.V2C_4 (V2C_281_98),
	.V2C_5 (V2C_281_172),
	.V2C_6 (V2C_281_221),
	.V (V_281)
);

VNU_6 #(quan_width) VNU282 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_282),
	.C2V_2 (C2V_48_282),
	.C2V_3 (C2V_87_282),
	.C2V_4 (C2V_104_282),
	.C2V_5 (C2V_178_282),
	.C2V_6 (C2V_227_282),
	.L (L_282),
	.V2C_1 (V2C_282_43),
	.V2C_2 (V2C_282_48),
	.V2C_3 (V2C_282_87),
	.V2C_4 (V2C_282_104),
	.V2C_5 (V2C_282_178),
	.V2C_6 (V2C_282_227),
	.V (V_282)
);

VNU_6 #(quan_width) VNU283 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_283),
	.C2V_2 (C2V_54_283),
	.C2V_3 (C2V_93_283),
	.C2V_4 (C2V_110_283),
	.C2V_5 (C2V_184_283),
	.C2V_6 (C2V_233_283),
	.L (L_283),
	.V2C_1 (V2C_283_49),
	.V2C_2 (V2C_283_54),
	.V2C_3 (V2C_283_93),
	.V2C_4 (V2C_283_110),
	.V2C_5 (V2C_283_184),
	.V2C_6 (V2C_283_233),
	.V (V_283)
);

VNU_6 #(quan_width) VNU284 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_284),
	.C2V_2 (C2V_60_284),
	.C2V_3 (C2V_99_284),
	.C2V_4 (C2V_116_284),
	.C2V_5 (C2V_190_284),
	.C2V_6 (C2V_239_284),
	.L (L_284),
	.V2C_1 (V2C_284_55),
	.V2C_2 (V2C_284_60),
	.V2C_3 (V2C_284_99),
	.V2C_4 (V2C_284_116),
	.V2C_5 (V2C_284_190),
	.V2C_6 (V2C_284_239),
	.V (V_284)
);

VNU_6 #(quan_width) VNU285 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_285),
	.C2V_2 (C2V_66_285),
	.C2V_3 (C2V_105_285),
	.C2V_4 (C2V_122_285),
	.C2V_5 (C2V_196_285),
	.C2V_6 (C2V_245_285),
	.L (L_285),
	.V2C_1 (V2C_285_61),
	.V2C_2 (V2C_285_66),
	.V2C_3 (V2C_285_105),
	.V2C_4 (V2C_285_122),
	.V2C_5 (V2C_285_196),
	.V2C_6 (V2C_285_245),
	.V (V_285)
);

VNU_6 #(quan_width) VNU286 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_286),
	.C2V_2 (C2V_72_286),
	.C2V_3 (C2V_111_286),
	.C2V_4 (C2V_128_286),
	.C2V_5 (C2V_202_286),
	.C2V_6 (C2V_251_286),
	.L (L_286),
	.V2C_1 (V2C_286_67),
	.V2C_2 (V2C_286_72),
	.V2C_3 (V2C_286_111),
	.V2C_4 (V2C_286_128),
	.V2C_5 (V2C_286_202),
	.V2C_6 (V2C_286_251),
	.V (V_286)
);

VNU_6 #(quan_width) VNU287 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_287),
	.C2V_2 (C2V_78_287),
	.C2V_3 (C2V_117_287),
	.C2V_4 (C2V_134_287),
	.C2V_5 (C2V_208_287),
	.C2V_6 (C2V_257_287),
	.L (L_287),
	.V2C_1 (V2C_287_73),
	.V2C_2 (V2C_287_78),
	.V2C_3 (V2C_287_117),
	.V2C_4 (V2C_287_134),
	.V2C_5 (V2C_287_208),
	.V2C_6 (V2C_287_257),
	.V (V_287)
);

VNU_6 #(quan_width) VNU288 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_288),
	.C2V_2 (C2V_84_288),
	.C2V_3 (C2V_123_288),
	.C2V_4 (C2V_140_288),
	.C2V_5 (C2V_214_288),
	.C2V_6 (C2V_263_288),
	.L (L_288),
	.V2C_1 (V2C_288_79),
	.V2C_2 (V2C_288_84),
	.V2C_3 (V2C_288_123),
	.V2C_4 (V2C_288_140),
	.V2C_5 (V2C_288_214),
	.V2C_6 (V2C_288_263),
	.V (V_288)
);

VNU_3 #(quan_width) VNU289 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_60_289),
	.C2V_2 (C2V_128_289),
	.C2V_3 (C2V_263_289),
	.L (L_289),
	.V2C_1 (V2C_289_60),
	.V2C_2 (V2C_289_128),
	.V2C_3 (V2C_289_263),
	.V (V_289)
);

VNU_3 #(quan_width) VNU290 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_66_290),
	.C2V_2 (C2V_134_290),
	.C2V_3 (C2V_269_290),
	.L (L_290),
	.V2C_1 (V2C_290_66),
	.V2C_2 (V2C_290_134),
	.V2C_3 (V2C_290_269),
	.V (V_290)
);

VNU_3 #(quan_width) VNU291 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_72_291),
	.C2V_2 (C2V_140_291),
	.C2V_3 (C2V_275_291),
	.L (L_291),
	.V2C_1 (V2C_291_72),
	.V2C_2 (V2C_291_140),
	.V2C_3 (V2C_291_275),
	.V (V_291)
);

VNU_3 #(quan_width) VNU292 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_78_292),
	.C2V_2 (C2V_146_292),
	.C2V_3 (C2V_281_292),
	.L (L_292),
	.V2C_1 (V2C_292_78),
	.V2C_2 (V2C_292_146),
	.V2C_3 (V2C_292_281),
	.V (V_292)
);

VNU_3 #(quan_width) VNU293 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_84_293),
	.C2V_2 (C2V_152_293),
	.C2V_3 (C2V_287_293),
	.L (L_293),
	.V2C_1 (V2C_293_84),
	.V2C_2 (V2C_293_152),
	.V2C_3 (V2C_293_287),
	.V (V_293)
);

VNU_3 #(quan_width) VNU294 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_294),
	.C2V_2 (C2V_90_294),
	.C2V_3 (C2V_158_294),
	.L (L_294),
	.V2C_1 (V2C_294_5),
	.V2C_2 (V2C_294_90),
	.V2C_3 (V2C_294_158),
	.V (V_294)
);

VNU_3 #(quan_width) VNU295 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_295),
	.C2V_2 (C2V_96_295),
	.C2V_3 (C2V_164_295),
	.L (L_295),
	.V2C_1 (V2C_295_11),
	.V2C_2 (V2C_295_96),
	.V2C_3 (V2C_295_164),
	.V (V_295)
);

VNU_3 #(quan_width) VNU296 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_296),
	.C2V_2 (C2V_102_296),
	.C2V_3 (C2V_170_296),
	.L (L_296),
	.V2C_1 (V2C_296_17),
	.V2C_2 (V2C_296_102),
	.V2C_3 (V2C_296_170),
	.V (V_296)
);

VNU_3 #(quan_width) VNU297 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_297),
	.C2V_2 (C2V_108_297),
	.C2V_3 (C2V_176_297),
	.L (L_297),
	.V2C_1 (V2C_297_23),
	.V2C_2 (V2C_297_108),
	.V2C_3 (V2C_297_176),
	.V (V_297)
);

VNU_3 #(quan_width) VNU298 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_298),
	.C2V_2 (C2V_114_298),
	.C2V_3 (C2V_182_298),
	.L (L_298),
	.V2C_1 (V2C_298_29),
	.V2C_2 (V2C_298_114),
	.V2C_3 (V2C_298_182),
	.V (V_298)
);

VNU_3 #(quan_width) VNU299 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_299),
	.C2V_2 (C2V_120_299),
	.C2V_3 (C2V_188_299),
	.L (L_299),
	.V2C_1 (V2C_299_35),
	.V2C_2 (V2C_299_120),
	.V2C_3 (V2C_299_188),
	.V (V_299)
);

VNU_3 #(quan_width) VNU300 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_300),
	.C2V_2 (C2V_126_300),
	.C2V_3 (C2V_194_300),
	.L (L_300),
	.V2C_1 (V2C_300_41),
	.V2C_2 (V2C_300_126),
	.V2C_3 (V2C_300_194),
	.V (V_300)
);

VNU_3 #(quan_width) VNU301 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_301),
	.C2V_2 (C2V_132_301),
	.C2V_3 (C2V_200_301),
	.L (L_301),
	.V2C_1 (V2C_301_47),
	.V2C_2 (V2C_301_132),
	.V2C_3 (V2C_301_200),
	.V (V_301)
);

VNU_3 #(quan_width) VNU302 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_302),
	.C2V_2 (C2V_138_302),
	.C2V_3 (C2V_206_302),
	.L (L_302),
	.V2C_1 (V2C_302_53),
	.V2C_2 (V2C_302_138),
	.V2C_3 (V2C_302_206),
	.V (V_302)
);

VNU_3 #(quan_width) VNU303 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_59_303),
	.C2V_2 (C2V_144_303),
	.C2V_3 (C2V_212_303),
	.L (L_303),
	.V2C_1 (V2C_303_59),
	.V2C_2 (V2C_303_144),
	.V2C_3 (V2C_303_212),
	.V (V_303)
);

VNU_3 #(quan_width) VNU304 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_65_304),
	.C2V_2 (C2V_150_304),
	.C2V_3 (C2V_218_304),
	.L (L_304),
	.V2C_1 (V2C_304_65),
	.V2C_2 (V2C_304_150),
	.V2C_3 (V2C_304_218),
	.V (V_304)
);

VNU_3 #(quan_width) VNU305 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_71_305),
	.C2V_2 (C2V_156_305),
	.C2V_3 (C2V_224_305),
	.L (L_305),
	.V2C_1 (V2C_305_71),
	.V2C_2 (V2C_305_156),
	.V2C_3 (V2C_305_224),
	.V (V_305)
);

VNU_3 #(quan_width) VNU306 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_77_306),
	.C2V_2 (C2V_162_306),
	.C2V_3 (C2V_230_306),
	.L (L_306),
	.V2C_1 (V2C_306_77),
	.V2C_2 (V2C_306_162),
	.V2C_3 (V2C_306_230),
	.V (V_306)
);

VNU_3 #(quan_width) VNU307 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_83_307),
	.C2V_2 (C2V_168_307),
	.C2V_3 (C2V_236_307),
	.L (L_307),
	.V2C_1 (V2C_307_83),
	.V2C_2 (V2C_307_168),
	.V2C_3 (V2C_307_236),
	.V (V_307)
);

VNU_3 #(quan_width) VNU308 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_89_308),
	.C2V_2 (C2V_174_308),
	.C2V_3 (C2V_242_308),
	.L (L_308),
	.V2C_1 (V2C_308_89),
	.V2C_2 (V2C_308_174),
	.V2C_3 (V2C_308_242),
	.V (V_308)
);

VNU_3 #(quan_width) VNU309 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_95_309),
	.C2V_2 (C2V_180_309),
	.C2V_3 (C2V_248_309),
	.L (L_309),
	.V2C_1 (V2C_309_95),
	.V2C_2 (V2C_309_180),
	.V2C_3 (V2C_309_248),
	.V (V_309)
);

VNU_3 #(quan_width) VNU310 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_101_310),
	.C2V_2 (C2V_186_310),
	.C2V_3 (C2V_254_310),
	.L (L_310),
	.V2C_1 (V2C_310_101),
	.V2C_2 (V2C_310_186),
	.V2C_3 (V2C_310_254),
	.V (V_310)
);

VNU_3 #(quan_width) VNU311 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_107_311),
	.C2V_2 (C2V_192_311),
	.C2V_3 (C2V_260_311),
	.L (L_311),
	.V2C_1 (V2C_311_107),
	.V2C_2 (V2C_311_192),
	.V2C_3 (V2C_311_260),
	.V (V_311)
);

VNU_3 #(quan_width) VNU312 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_113_312),
	.C2V_2 (C2V_198_312),
	.C2V_3 (C2V_266_312),
	.L (L_312),
	.V2C_1 (V2C_312_113),
	.V2C_2 (V2C_312_198),
	.V2C_3 (V2C_312_266),
	.V (V_312)
);

VNU_3 #(quan_width) VNU313 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_119_313),
	.C2V_2 (C2V_204_313),
	.C2V_3 (C2V_272_313),
	.L (L_313),
	.V2C_1 (V2C_313_119),
	.V2C_2 (V2C_313_204),
	.V2C_3 (V2C_313_272),
	.V (V_313)
);

VNU_3 #(quan_width) VNU314 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_125_314),
	.C2V_2 (C2V_210_314),
	.C2V_3 (C2V_278_314),
	.L (L_314),
	.V2C_1 (V2C_314_125),
	.V2C_2 (V2C_314_210),
	.V2C_3 (V2C_314_278),
	.V (V_314)
);

VNU_3 #(quan_width) VNU315 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_131_315),
	.C2V_2 (C2V_216_315),
	.C2V_3 (C2V_284_315),
	.L (L_315),
	.V2C_1 (V2C_315_131),
	.V2C_2 (V2C_315_216),
	.V2C_3 (V2C_315_284),
	.V (V_315)
);

VNU_3 #(quan_width) VNU316 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_316),
	.C2V_2 (C2V_137_316),
	.C2V_3 (C2V_222_316),
	.L (L_316),
	.V2C_1 (V2C_316_2),
	.V2C_2 (V2C_316_137),
	.V2C_3 (V2C_316_222),
	.V (V_316)
);

VNU_3 #(quan_width) VNU317 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_317),
	.C2V_2 (C2V_143_317),
	.C2V_3 (C2V_228_317),
	.L (L_317),
	.V2C_1 (V2C_317_8),
	.V2C_2 (V2C_317_143),
	.V2C_3 (V2C_317_228),
	.V (V_317)
);

VNU_3 #(quan_width) VNU318 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_318),
	.C2V_2 (C2V_149_318),
	.C2V_3 (C2V_234_318),
	.L (L_318),
	.V2C_1 (V2C_318_14),
	.V2C_2 (V2C_318_149),
	.V2C_3 (V2C_318_234),
	.V (V_318)
);

VNU_3 #(quan_width) VNU319 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_319),
	.C2V_2 (C2V_155_319),
	.C2V_3 (C2V_240_319),
	.L (L_319),
	.V2C_1 (V2C_319_20),
	.V2C_2 (V2C_319_155),
	.V2C_3 (V2C_319_240),
	.V (V_319)
);

VNU_3 #(quan_width) VNU320 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_320),
	.C2V_2 (C2V_161_320),
	.C2V_3 (C2V_246_320),
	.L (L_320),
	.V2C_1 (V2C_320_26),
	.V2C_2 (V2C_320_161),
	.V2C_3 (V2C_320_246),
	.V (V_320)
);

VNU_3 #(quan_width) VNU321 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_321),
	.C2V_2 (C2V_167_321),
	.C2V_3 (C2V_252_321),
	.L (L_321),
	.V2C_1 (V2C_321_32),
	.V2C_2 (V2C_321_167),
	.V2C_3 (V2C_321_252),
	.V (V_321)
);

VNU_3 #(quan_width) VNU322 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_322),
	.C2V_2 (C2V_173_322),
	.C2V_3 (C2V_258_322),
	.L (L_322),
	.V2C_1 (V2C_322_38),
	.V2C_2 (V2C_322_173),
	.V2C_3 (V2C_322_258),
	.V (V_322)
);

VNU_3 #(quan_width) VNU323 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_323),
	.C2V_2 (C2V_179_323),
	.C2V_3 (C2V_264_323),
	.L (L_323),
	.V2C_1 (V2C_323_44),
	.V2C_2 (V2C_323_179),
	.V2C_3 (V2C_323_264),
	.V (V_323)
);

VNU_3 #(quan_width) VNU324 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_324),
	.C2V_2 (C2V_185_324),
	.C2V_3 (C2V_270_324),
	.L (L_324),
	.V2C_1 (V2C_324_50),
	.V2C_2 (V2C_324_185),
	.V2C_3 (V2C_324_270),
	.V (V_324)
);

VNU_3 #(quan_width) VNU325 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_325),
	.C2V_2 (C2V_191_325),
	.C2V_3 (C2V_276_325),
	.L (L_325),
	.V2C_1 (V2C_325_56),
	.V2C_2 (V2C_325_191),
	.V2C_3 (V2C_325_276),
	.V (V_325)
);

VNU_3 #(quan_width) VNU326 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_326),
	.C2V_2 (C2V_197_326),
	.C2V_3 (C2V_282_326),
	.L (L_326),
	.V2C_1 (V2C_326_62),
	.V2C_2 (V2C_326_197),
	.V2C_3 (V2C_326_282),
	.V (V_326)
);

VNU_3 #(quan_width) VNU327 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_327),
	.C2V_2 (C2V_203_327),
	.C2V_3 (C2V_288_327),
	.L (L_327),
	.V2C_1 (V2C_327_68),
	.V2C_2 (V2C_327_203),
	.V2C_3 (V2C_327_288),
	.V (V_327)
);

VNU_3 #(quan_width) VNU328 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_328),
	.C2V_2 (C2V_74_328),
	.C2V_3 (C2V_209_328),
	.L (L_328),
	.V2C_1 (V2C_328_6),
	.V2C_2 (V2C_328_74),
	.V2C_3 (V2C_328_209),
	.V (V_328)
);

VNU_3 #(quan_width) VNU329 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_329),
	.C2V_2 (C2V_80_329),
	.C2V_3 (C2V_215_329),
	.L (L_329),
	.V2C_1 (V2C_329_12),
	.V2C_2 (V2C_329_80),
	.V2C_3 (V2C_329_215),
	.V (V_329)
);

VNU_3 #(quan_width) VNU330 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_330),
	.C2V_2 (C2V_86_330),
	.C2V_3 (C2V_221_330),
	.L (L_330),
	.V2C_1 (V2C_330_18),
	.V2C_2 (V2C_330_86),
	.V2C_3 (V2C_330_221),
	.V (V_330)
);

VNU_3 #(quan_width) VNU331 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_331),
	.C2V_2 (C2V_92_331),
	.C2V_3 (C2V_227_331),
	.L (L_331),
	.V2C_1 (V2C_331_24),
	.V2C_2 (V2C_331_92),
	.V2C_3 (V2C_331_227),
	.V (V_331)
);

VNU_3 #(quan_width) VNU332 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_332),
	.C2V_2 (C2V_98_332),
	.C2V_3 (C2V_233_332),
	.L (L_332),
	.V2C_1 (V2C_332_30),
	.V2C_2 (V2C_332_98),
	.V2C_3 (V2C_332_233),
	.V (V_332)
);

VNU_3 #(quan_width) VNU333 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_333),
	.C2V_2 (C2V_104_333),
	.C2V_3 (C2V_239_333),
	.L (L_333),
	.V2C_1 (V2C_333_36),
	.V2C_2 (V2C_333_104),
	.V2C_3 (V2C_333_239),
	.V (V_333)
);

VNU_3 #(quan_width) VNU334 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_334),
	.C2V_2 (C2V_110_334),
	.C2V_3 (C2V_245_334),
	.L (L_334),
	.V2C_1 (V2C_334_42),
	.V2C_2 (V2C_334_110),
	.V2C_3 (V2C_334_245),
	.V (V_334)
);

VNU_3 #(quan_width) VNU335 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_335),
	.C2V_2 (C2V_116_335),
	.C2V_3 (C2V_251_335),
	.L (L_335),
	.V2C_1 (V2C_335_48),
	.V2C_2 (V2C_335_116),
	.V2C_3 (V2C_335_251),
	.V (V_335)
);

VNU_3 #(quan_width) VNU336 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_54_336),
	.C2V_2 (C2V_122_336),
	.C2V_3 (C2V_257_336),
	.L (L_336),
	.V2C_1 (V2C_336_54),
	.V2C_2 (V2C_336_122),
	.V2C_3 (V2C_336_257),
	.V (V_336)
);

VNU_3 #(quan_width) VNU337 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_337),
	.C2V_2 (C2V_123_337),
	.C2V_3 (C2V_149_337),
	.L (L_337),
	.V2C_1 (V2C_337_61),
	.V2C_2 (V2C_337_123),
	.V2C_3 (V2C_337_149),
	.V (V_337)
);

VNU_3 #(quan_width) VNU338 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_338),
	.C2V_2 (C2V_129_338),
	.C2V_3 (C2V_155_338),
	.L (L_338),
	.V2C_1 (V2C_338_67),
	.V2C_2 (V2C_338_129),
	.V2C_3 (V2C_338_155),
	.V (V_338)
);

VNU_3 #(quan_width) VNU339 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_339),
	.C2V_2 (C2V_135_339),
	.C2V_3 (C2V_161_339),
	.L (L_339),
	.V2C_1 (V2C_339_73),
	.V2C_2 (V2C_339_135),
	.V2C_3 (V2C_339_161),
	.V (V_339)
);

VNU_3 #(quan_width) VNU340 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_340),
	.C2V_2 (C2V_141_340),
	.C2V_3 (C2V_167_340),
	.L (L_340),
	.V2C_1 (V2C_340_79),
	.V2C_2 (V2C_340_141),
	.V2C_3 (V2C_340_167),
	.V (V_340)
);

VNU_3 #(quan_width) VNU341 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_341),
	.C2V_2 (C2V_147_341),
	.C2V_3 (C2V_173_341),
	.L (L_341),
	.V2C_1 (V2C_341_85),
	.V2C_2 (V2C_341_147),
	.V2C_3 (V2C_341_173),
	.V (V_341)
);

VNU_3 #(quan_width) VNU342 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_91_342),
	.C2V_2 (C2V_153_342),
	.C2V_3 (C2V_179_342),
	.L (L_342),
	.V2C_1 (V2C_342_91),
	.V2C_2 (V2C_342_153),
	.V2C_3 (V2C_342_179),
	.V (V_342)
);

VNU_3 #(quan_width) VNU343 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_97_343),
	.C2V_2 (C2V_159_343),
	.C2V_3 (C2V_185_343),
	.L (L_343),
	.V2C_1 (V2C_343_97),
	.V2C_2 (V2C_343_159),
	.V2C_3 (V2C_343_185),
	.V (V_343)
);

VNU_3 #(quan_width) VNU344 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_103_344),
	.C2V_2 (C2V_165_344),
	.C2V_3 (C2V_191_344),
	.L (L_344),
	.V2C_1 (V2C_344_103),
	.V2C_2 (V2C_344_165),
	.V2C_3 (V2C_344_191),
	.V (V_344)
);

VNU_3 #(quan_width) VNU345 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_109_345),
	.C2V_2 (C2V_171_345),
	.C2V_3 (C2V_197_345),
	.L (L_345),
	.V2C_1 (V2C_345_109),
	.V2C_2 (V2C_345_171),
	.V2C_3 (V2C_345_197),
	.V (V_345)
);

VNU_3 #(quan_width) VNU346 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_115_346),
	.C2V_2 (C2V_177_346),
	.C2V_3 (C2V_203_346),
	.L (L_346),
	.V2C_1 (V2C_346_115),
	.V2C_2 (V2C_346_177),
	.V2C_3 (V2C_346_203),
	.V (V_346)
);

VNU_3 #(quan_width) VNU347 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_121_347),
	.C2V_2 (C2V_183_347),
	.C2V_3 (C2V_209_347),
	.L (L_347),
	.V2C_1 (V2C_347_121),
	.V2C_2 (V2C_347_183),
	.V2C_3 (V2C_347_209),
	.V (V_347)
);

VNU_3 #(quan_width) VNU348 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_127_348),
	.C2V_2 (C2V_189_348),
	.C2V_3 (C2V_215_348),
	.L (L_348),
	.V2C_1 (V2C_348_127),
	.V2C_2 (V2C_348_189),
	.V2C_3 (V2C_348_215),
	.V (V_348)
);

VNU_3 #(quan_width) VNU349 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_133_349),
	.C2V_2 (C2V_195_349),
	.C2V_3 (C2V_221_349),
	.L (L_349),
	.V2C_1 (V2C_349_133),
	.V2C_2 (V2C_349_195),
	.V2C_3 (V2C_349_221),
	.V (V_349)
);

VNU_3 #(quan_width) VNU350 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_139_350),
	.C2V_2 (C2V_201_350),
	.C2V_3 (C2V_227_350),
	.L (L_350),
	.V2C_1 (V2C_350_139),
	.V2C_2 (V2C_350_201),
	.V2C_3 (V2C_350_227),
	.V (V_350)
);

VNU_3 #(quan_width) VNU351 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_145_351),
	.C2V_2 (C2V_207_351),
	.C2V_3 (C2V_233_351),
	.L (L_351),
	.V2C_1 (V2C_351_145),
	.V2C_2 (V2C_351_207),
	.V2C_3 (V2C_351_233),
	.V (V_351)
);

VNU_3 #(quan_width) VNU352 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_151_352),
	.C2V_2 (C2V_213_352),
	.C2V_3 (C2V_239_352),
	.L (L_352),
	.V2C_1 (V2C_352_151),
	.V2C_2 (V2C_352_213),
	.V2C_3 (V2C_352_239),
	.V (V_352)
);

VNU_3 #(quan_width) VNU353 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_157_353),
	.C2V_2 (C2V_219_353),
	.C2V_3 (C2V_245_353),
	.L (L_353),
	.V2C_1 (V2C_353_157),
	.V2C_2 (V2C_353_219),
	.V2C_3 (V2C_353_245),
	.V (V_353)
);

VNU_3 #(quan_width) VNU354 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_163_354),
	.C2V_2 (C2V_225_354),
	.C2V_3 (C2V_251_354),
	.L (L_354),
	.V2C_1 (V2C_354_163),
	.V2C_2 (V2C_354_225),
	.V2C_3 (V2C_354_251),
	.V (V_354)
);

VNU_3 #(quan_width) VNU355 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_169_355),
	.C2V_2 (C2V_231_355),
	.C2V_3 (C2V_257_355),
	.L (L_355),
	.V2C_1 (V2C_355_169),
	.V2C_2 (V2C_355_231),
	.V2C_3 (V2C_355_257),
	.V (V_355)
);

VNU_3 #(quan_width) VNU356 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_175_356),
	.C2V_2 (C2V_237_356),
	.C2V_3 (C2V_263_356),
	.L (L_356),
	.V2C_1 (V2C_356_175),
	.V2C_2 (V2C_356_237),
	.V2C_3 (V2C_356_263),
	.V (V_356)
);

VNU_3 #(quan_width) VNU357 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_181_357),
	.C2V_2 (C2V_243_357),
	.C2V_3 (C2V_269_357),
	.L (L_357),
	.V2C_1 (V2C_357_181),
	.V2C_2 (V2C_357_243),
	.V2C_3 (V2C_357_269),
	.V (V_357)
);

VNU_3 #(quan_width) VNU358 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_187_358),
	.C2V_2 (C2V_249_358),
	.C2V_3 (C2V_275_358),
	.L (L_358),
	.V2C_1 (V2C_358_187),
	.V2C_2 (V2C_358_249),
	.V2C_3 (V2C_358_275),
	.V (V_358)
);

VNU_3 #(quan_width) VNU359 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_193_359),
	.C2V_2 (C2V_255_359),
	.C2V_3 (C2V_281_359),
	.L (L_359),
	.V2C_1 (V2C_359_193),
	.V2C_2 (V2C_359_255),
	.V2C_3 (V2C_359_281),
	.V (V_359)
);

VNU_3 #(quan_width) VNU360 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_199_360),
	.C2V_2 (C2V_261_360),
	.C2V_3 (C2V_287_360),
	.L (L_360),
	.V2C_1 (V2C_360_199),
	.V2C_2 (V2C_360_261),
	.V2C_3 (V2C_360_287),
	.V (V_360)
);

VNU_3 #(quan_width) VNU361 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_361),
	.C2V_2 (C2V_205_361),
	.C2V_3 (C2V_267_361),
	.L (L_361),
	.V2C_1 (V2C_361_5),
	.V2C_2 (V2C_361_205),
	.V2C_3 (V2C_361_267),
	.V (V_361)
);

VNU_3 #(quan_width) VNU362 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_362),
	.C2V_2 (C2V_211_362),
	.C2V_3 (C2V_273_362),
	.L (L_362),
	.V2C_1 (V2C_362_11),
	.V2C_2 (V2C_362_211),
	.V2C_3 (V2C_362_273),
	.V (V_362)
);

VNU_3 #(quan_width) VNU363 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_363),
	.C2V_2 (C2V_217_363),
	.C2V_3 (C2V_279_363),
	.L (L_363),
	.V2C_1 (V2C_363_17),
	.V2C_2 (V2C_363_217),
	.V2C_3 (V2C_363_279),
	.V (V_363)
);

VNU_3 #(quan_width) VNU364 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_364),
	.C2V_2 (C2V_223_364),
	.C2V_3 (C2V_285_364),
	.L (L_364),
	.V2C_1 (V2C_364_23),
	.V2C_2 (V2C_364_223),
	.V2C_3 (V2C_364_285),
	.V (V_364)
);

VNU_3 #(quan_width) VNU365 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_365),
	.C2V_2 (C2V_29_365),
	.C2V_3 (C2V_229_365),
	.L (L_365),
	.V2C_1 (V2C_365_3),
	.V2C_2 (V2C_365_29),
	.V2C_3 (V2C_365_229),
	.V (V_365)
);

VNU_3 #(quan_width) VNU366 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_366),
	.C2V_2 (C2V_35_366),
	.C2V_3 (C2V_235_366),
	.L (L_366),
	.V2C_1 (V2C_366_9),
	.V2C_2 (V2C_366_35),
	.V2C_3 (V2C_366_235),
	.V (V_366)
);

VNU_3 #(quan_width) VNU367 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_367),
	.C2V_2 (C2V_41_367),
	.C2V_3 (C2V_241_367),
	.L (L_367),
	.V2C_1 (V2C_367_15),
	.V2C_2 (V2C_367_41),
	.V2C_3 (V2C_367_241),
	.V (V_367)
);

VNU_3 #(quan_width) VNU368 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_368),
	.C2V_2 (C2V_47_368),
	.C2V_3 (C2V_247_368),
	.L (L_368),
	.V2C_1 (V2C_368_21),
	.V2C_2 (V2C_368_47),
	.V2C_3 (V2C_368_247),
	.V (V_368)
);

VNU_3 #(quan_width) VNU369 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_369),
	.C2V_2 (C2V_53_369),
	.C2V_3 (C2V_253_369),
	.L (L_369),
	.V2C_1 (V2C_369_27),
	.V2C_2 (V2C_369_53),
	.V2C_3 (V2C_369_253),
	.V (V_369)
);

VNU_3 #(quan_width) VNU370 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_370),
	.C2V_2 (C2V_59_370),
	.C2V_3 (C2V_259_370),
	.L (L_370),
	.V2C_1 (V2C_370_33),
	.V2C_2 (V2C_370_59),
	.V2C_3 (V2C_370_259),
	.V (V_370)
);

VNU_3 #(quan_width) VNU371 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_371),
	.C2V_2 (C2V_65_371),
	.C2V_3 (C2V_265_371),
	.L (L_371),
	.V2C_1 (V2C_371_39),
	.V2C_2 (V2C_371_65),
	.V2C_3 (V2C_371_265),
	.V (V_371)
);

VNU_3 #(quan_width) VNU372 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_372),
	.C2V_2 (C2V_71_372),
	.C2V_3 (C2V_271_372),
	.L (L_372),
	.V2C_1 (V2C_372_45),
	.V2C_2 (V2C_372_71),
	.V2C_3 (V2C_372_271),
	.V (V_372)
);

VNU_3 #(quan_width) VNU373 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_373),
	.C2V_2 (C2V_77_373),
	.C2V_3 (C2V_277_373),
	.L (L_373),
	.V2C_1 (V2C_373_51),
	.V2C_2 (V2C_373_77),
	.V2C_3 (V2C_373_277),
	.V (V_373)
);

VNU_3 #(quan_width) VNU374 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_374),
	.C2V_2 (C2V_83_374),
	.C2V_3 (C2V_283_374),
	.L (L_374),
	.V2C_1 (V2C_374_57),
	.V2C_2 (V2C_374_83),
	.V2C_3 (V2C_374_283),
	.V (V_374)
);

VNU_3 #(quan_width) VNU375 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_375),
	.C2V_2 (C2V_63_375),
	.C2V_3 (C2V_89_375),
	.L (L_375),
	.V2C_1 (V2C_375_1),
	.V2C_2 (V2C_375_63),
	.V2C_3 (V2C_375_89),
	.V (V_375)
);

VNU_3 #(quan_width) VNU376 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_376),
	.C2V_2 (C2V_69_376),
	.C2V_3 (C2V_95_376),
	.L (L_376),
	.V2C_1 (V2C_376_7),
	.V2C_2 (V2C_376_69),
	.V2C_3 (V2C_376_95),
	.V (V_376)
);

VNU_3 #(quan_width) VNU377 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_377),
	.C2V_2 (C2V_75_377),
	.C2V_3 (C2V_101_377),
	.L (L_377),
	.V2C_1 (V2C_377_13),
	.V2C_2 (V2C_377_75),
	.V2C_3 (V2C_377_101),
	.V (V_377)
);

VNU_3 #(quan_width) VNU378 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_378),
	.C2V_2 (C2V_81_378),
	.C2V_3 (C2V_107_378),
	.L (L_378),
	.V2C_1 (V2C_378_19),
	.V2C_2 (V2C_378_81),
	.V2C_3 (V2C_378_107),
	.V (V_378)
);

VNU_3 #(quan_width) VNU379 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_379),
	.C2V_2 (C2V_87_379),
	.C2V_3 (C2V_113_379),
	.L (L_379),
	.V2C_1 (V2C_379_25),
	.V2C_2 (V2C_379_87),
	.V2C_3 (V2C_379_113),
	.V (V_379)
);

VNU_3 #(quan_width) VNU380 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_380),
	.C2V_2 (C2V_93_380),
	.C2V_3 (C2V_119_380),
	.L (L_380),
	.V2C_1 (V2C_380_31),
	.V2C_2 (V2C_380_93),
	.V2C_3 (V2C_380_119),
	.V (V_380)
);

VNU_3 #(quan_width) VNU381 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_381),
	.C2V_2 (C2V_99_381),
	.C2V_3 (C2V_125_381),
	.L (L_381),
	.V2C_1 (V2C_381_37),
	.V2C_2 (V2C_381_99),
	.V2C_3 (V2C_381_125),
	.V (V_381)
);

VNU_3 #(quan_width) VNU382 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_382),
	.C2V_2 (C2V_105_382),
	.C2V_3 (C2V_131_382),
	.L (L_382),
	.V2C_1 (V2C_382_43),
	.V2C_2 (V2C_382_105),
	.V2C_3 (V2C_382_131),
	.V (V_382)
);

VNU_3 #(quan_width) VNU383 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_383),
	.C2V_2 (C2V_111_383),
	.C2V_3 (C2V_137_383),
	.L (L_383),
	.V2C_1 (V2C_383_49),
	.V2C_2 (V2C_383_111),
	.V2C_3 (V2C_383_137),
	.V (V_383)
);

VNU_3 #(quan_width) VNU384 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_384),
	.C2V_2 (C2V_117_384),
	.C2V_3 (C2V_143_384),
	.L (L_384),
	.V2C_1 (V2C_384_55),
	.V2C_2 (V2C_384_117),
	.V2C_3 (V2C_384_143),
	.V (V_384)
);

VNU_3 #(quan_width) VNU385 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_385),
	.C2V_2 (C2V_62_385),
	.C2V_3 (C2V_81_385),
	.L (L_385),
	.V2C_1 (V2C_385_25),
	.V2C_2 (V2C_385_62),
	.V2C_3 (V2C_385_81),
	.V (V_385)
);

VNU_3 #(quan_width) VNU386 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_386),
	.C2V_2 (C2V_68_386),
	.C2V_3 (C2V_87_386),
	.L (L_386),
	.V2C_1 (V2C_386_31),
	.V2C_2 (V2C_386_68),
	.V2C_3 (V2C_386_87),
	.V (V_386)
);

VNU_3 #(quan_width) VNU387 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_387),
	.C2V_2 (C2V_74_387),
	.C2V_3 (C2V_93_387),
	.L (L_387),
	.V2C_1 (V2C_387_37),
	.V2C_2 (V2C_387_74),
	.V2C_3 (V2C_387_93),
	.V (V_387)
);

VNU_3 #(quan_width) VNU388 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_388),
	.C2V_2 (C2V_80_388),
	.C2V_3 (C2V_99_388),
	.L (L_388),
	.V2C_1 (V2C_388_43),
	.V2C_2 (V2C_388_80),
	.V2C_3 (V2C_388_99),
	.V (V_388)
);

VNU_3 #(quan_width) VNU389 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_389),
	.C2V_2 (C2V_86_389),
	.C2V_3 (C2V_105_389),
	.L (L_389),
	.V2C_1 (V2C_389_49),
	.V2C_2 (V2C_389_86),
	.V2C_3 (V2C_389_105),
	.V (V_389)
);

VNU_3 #(quan_width) VNU390 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_390),
	.C2V_2 (C2V_92_390),
	.C2V_3 (C2V_111_390),
	.L (L_390),
	.V2C_1 (V2C_390_55),
	.V2C_2 (V2C_390_92),
	.V2C_3 (V2C_390_111),
	.V (V_390)
);

VNU_3 #(quan_width) VNU391 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_391),
	.C2V_2 (C2V_98_391),
	.C2V_3 (C2V_117_391),
	.L (L_391),
	.V2C_1 (V2C_391_61),
	.V2C_2 (V2C_391_98),
	.V2C_3 (V2C_391_117),
	.V (V_391)
);

VNU_3 #(quan_width) VNU392 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_392),
	.C2V_2 (C2V_104_392),
	.C2V_3 (C2V_123_392),
	.L (L_392),
	.V2C_1 (V2C_392_67),
	.V2C_2 (V2C_392_104),
	.V2C_3 (V2C_392_123),
	.V (V_392)
);

VNU_3 #(quan_width) VNU393 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_393),
	.C2V_2 (C2V_110_393),
	.C2V_3 (C2V_129_393),
	.L (L_393),
	.V2C_1 (V2C_393_73),
	.V2C_2 (V2C_393_110),
	.V2C_3 (V2C_393_129),
	.V (V_393)
);

VNU_3 #(quan_width) VNU394 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_394),
	.C2V_2 (C2V_116_394),
	.C2V_3 (C2V_135_394),
	.L (L_394),
	.V2C_1 (V2C_394_79),
	.V2C_2 (V2C_394_116),
	.V2C_3 (V2C_394_135),
	.V (V_394)
);

VNU_3 #(quan_width) VNU395 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_395),
	.C2V_2 (C2V_122_395),
	.C2V_3 (C2V_141_395),
	.L (L_395),
	.V2C_1 (V2C_395_85),
	.V2C_2 (V2C_395_122),
	.V2C_3 (V2C_395_141),
	.V (V_395)
);

VNU_3 #(quan_width) VNU396 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_91_396),
	.C2V_2 (C2V_128_396),
	.C2V_3 (C2V_147_396),
	.L (L_396),
	.V2C_1 (V2C_396_91),
	.V2C_2 (V2C_396_128),
	.V2C_3 (V2C_396_147),
	.V (V_396)
);

VNU_3 #(quan_width) VNU397 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_97_397),
	.C2V_2 (C2V_134_397),
	.C2V_3 (C2V_153_397),
	.L (L_397),
	.V2C_1 (V2C_397_97),
	.V2C_2 (V2C_397_134),
	.V2C_3 (V2C_397_153),
	.V (V_397)
);

VNU_3 #(quan_width) VNU398 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_103_398),
	.C2V_2 (C2V_140_398),
	.C2V_3 (C2V_159_398),
	.L (L_398),
	.V2C_1 (V2C_398_103),
	.V2C_2 (V2C_398_140),
	.V2C_3 (V2C_398_159),
	.V (V_398)
);

VNU_3 #(quan_width) VNU399 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_109_399),
	.C2V_2 (C2V_146_399),
	.C2V_3 (C2V_165_399),
	.L (L_399),
	.V2C_1 (V2C_399_109),
	.V2C_2 (V2C_399_146),
	.V2C_3 (V2C_399_165),
	.V (V_399)
);

VNU_3 #(quan_width) VNU400 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_115_400),
	.C2V_2 (C2V_152_400),
	.C2V_3 (C2V_171_400),
	.L (L_400),
	.V2C_1 (V2C_400_115),
	.V2C_2 (V2C_400_152),
	.V2C_3 (V2C_400_171),
	.V (V_400)
);

VNU_3 #(quan_width) VNU401 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_121_401),
	.C2V_2 (C2V_158_401),
	.C2V_3 (C2V_177_401),
	.L (L_401),
	.V2C_1 (V2C_401_121),
	.V2C_2 (V2C_401_158),
	.V2C_3 (V2C_401_177),
	.V (V_401)
);

VNU_3 #(quan_width) VNU402 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_127_402),
	.C2V_2 (C2V_164_402),
	.C2V_3 (C2V_183_402),
	.L (L_402),
	.V2C_1 (V2C_402_127),
	.V2C_2 (V2C_402_164),
	.V2C_3 (V2C_402_183),
	.V (V_402)
);

VNU_3 #(quan_width) VNU403 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_133_403),
	.C2V_2 (C2V_170_403),
	.C2V_3 (C2V_189_403),
	.L (L_403),
	.V2C_1 (V2C_403_133),
	.V2C_2 (V2C_403_170),
	.V2C_3 (V2C_403_189),
	.V (V_403)
);

VNU_3 #(quan_width) VNU404 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_139_404),
	.C2V_2 (C2V_176_404),
	.C2V_3 (C2V_195_404),
	.L (L_404),
	.V2C_1 (V2C_404_139),
	.V2C_2 (V2C_404_176),
	.V2C_3 (V2C_404_195),
	.V (V_404)
);

VNU_3 #(quan_width) VNU405 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_145_405),
	.C2V_2 (C2V_182_405),
	.C2V_3 (C2V_201_405),
	.L (L_405),
	.V2C_1 (V2C_405_145),
	.V2C_2 (V2C_405_182),
	.V2C_3 (V2C_405_201),
	.V (V_405)
);

VNU_3 #(quan_width) VNU406 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_151_406),
	.C2V_2 (C2V_188_406),
	.C2V_3 (C2V_207_406),
	.L (L_406),
	.V2C_1 (V2C_406_151),
	.V2C_2 (V2C_406_188),
	.V2C_3 (V2C_406_207),
	.V (V_406)
);

VNU_3 #(quan_width) VNU407 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_157_407),
	.C2V_2 (C2V_194_407),
	.C2V_3 (C2V_213_407),
	.L (L_407),
	.V2C_1 (V2C_407_157),
	.V2C_2 (V2C_407_194),
	.V2C_3 (V2C_407_213),
	.V (V_407)
);

VNU_3 #(quan_width) VNU408 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_163_408),
	.C2V_2 (C2V_200_408),
	.C2V_3 (C2V_219_408),
	.L (L_408),
	.V2C_1 (V2C_408_163),
	.V2C_2 (V2C_408_200),
	.V2C_3 (V2C_408_219),
	.V (V_408)
);

VNU_3 #(quan_width) VNU409 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_169_409),
	.C2V_2 (C2V_206_409),
	.C2V_3 (C2V_225_409),
	.L (L_409),
	.V2C_1 (V2C_409_169),
	.V2C_2 (V2C_409_206),
	.V2C_3 (V2C_409_225),
	.V (V_409)
);

VNU_3 #(quan_width) VNU410 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_175_410),
	.C2V_2 (C2V_212_410),
	.C2V_3 (C2V_231_410),
	.L (L_410),
	.V2C_1 (V2C_410_175),
	.V2C_2 (V2C_410_212),
	.V2C_3 (V2C_410_231),
	.V (V_410)
);

VNU_3 #(quan_width) VNU411 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_181_411),
	.C2V_2 (C2V_218_411),
	.C2V_3 (C2V_237_411),
	.L (L_411),
	.V2C_1 (V2C_411_181),
	.V2C_2 (V2C_411_218),
	.V2C_3 (V2C_411_237),
	.V (V_411)
);

VNU_3 #(quan_width) VNU412 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_187_412),
	.C2V_2 (C2V_224_412),
	.C2V_3 (C2V_243_412),
	.L (L_412),
	.V2C_1 (V2C_412_187),
	.V2C_2 (V2C_412_224),
	.V2C_3 (V2C_412_243),
	.V (V_412)
);

VNU_3 #(quan_width) VNU413 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_193_413),
	.C2V_2 (C2V_230_413),
	.C2V_3 (C2V_249_413),
	.L (L_413),
	.V2C_1 (V2C_413_193),
	.V2C_2 (V2C_413_230),
	.V2C_3 (V2C_413_249),
	.V (V_413)
);

VNU_3 #(quan_width) VNU414 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_199_414),
	.C2V_2 (C2V_236_414),
	.C2V_3 (C2V_255_414),
	.L (L_414),
	.V2C_1 (V2C_414_199),
	.V2C_2 (V2C_414_236),
	.V2C_3 (V2C_414_255),
	.V (V_414)
);

VNU_3 #(quan_width) VNU415 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_205_415),
	.C2V_2 (C2V_242_415),
	.C2V_3 (C2V_261_415),
	.L (L_415),
	.V2C_1 (V2C_415_205),
	.V2C_2 (V2C_415_242),
	.V2C_3 (V2C_415_261),
	.V (V_415)
);

VNU_3 #(quan_width) VNU416 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_211_416),
	.C2V_2 (C2V_248_416),
	.C2V_3 (C2V_267_416),
	.L (L_416),
	.V2C_1 (V2C_416_211),
	.V2C_2 (V2C_416_248),
	.V2C_3 (V2C_416_267),
	.V (V_416)
);

VNU_3 #(quan_width) VNU417 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_217_417),
	.C2V_2 (C2V_254_417),
	.C2V_3 (C2V_273_417),
	.L (L_417),
	.V2C_1 (V2C_417_217),
	.V2C_2 (V2C_417_254),
	.V2C_3 (V2C_417_273),
	.V (V_417)
);

VNU_3 #(quan_width) VNU418 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_223_418),
	.C2V_2 (C2V_260_418),
	.C2V_3 (C2V_279_418),
	.L (L_418),
	.V2C_1 (V2C_418_223),
	.V2C_2 (V2C_418_260),
	.V2C_3 (V2C_418_279),
	.V (V_418)
);

VNU_3 #(quan_width) VNU419 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_229_419),
	.C2V_2 (C2V_266_419),
	.C2V_3 (C2V_285_419),
	.L (L_419),
	.V2C_1 (V2C_419_229),
	.V2C_2 (V2C_419_266),
	.V2C_3 (V2C_419_285),
	.V (V_419)
);

VNU_3 #(quan_width) VNU420 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_420),
	.C2V_2 (C2V_235_420),
	.C2V_3 (C2V_272_420),
	.L (L_420),
	.V2C_1 (V2C_420_3),
	.V2C_2 (V2C_420_235),
	.V2C_3 (V2C_420_272),
	.V (V_420)
);

VNU_3 #(quan_width) VNU421 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_421),
	.C2V_2 (C2V_241_421),
	.C2V_3 (C2V_278_421),
	.L (L_421),
	.V2C_1 (V2C_421_9),
	.V2C_2 (V2C_421_241),
	.V2C_3 (V2C_421_278),
	.V (V_421)
);

VNU_3 #(quan_width) VNU422 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_422),
	.C2V_2 (C2V_247_422),
	.C2V_3 (C2V_284_422),
	.L (L_422),
	.V2C_1 (V2C_422_15),
	.V2C_2 (V2C_422_247),
	.V2C_3 (V2C_422_284),
	.V (V_422)
);

VNU_3 #(quan_width) VNU423 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_423),
	.C2V_2 (C2V_21_423),
	.C2V_3 (C2V_253_423),
	.L (L_423),
	.V2C_1 (V2C_423_2),
	.V2C_2 (V2C_423_21),
	.V2C_3 (V2C_423_253),
	.V (V_423)
);

VNU_3 #(quan_width) VNU424 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_424),
	.C2V_2 (C2V_27_424),
	.C2V_3 (C2V_259_424),
	.L (L_424),
	.V2C_1 (V2C_424_8),
	.V2C_2 (V2C_424_27),
	.V2C_3 (V2C_424_259),
	.V (V_424)
);

VNU_3 #(quan_width) VNU425 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_425),
	.C2V_2 (C2V_33_425),
	.C2V_3 (C2V_265_425),
	.L (L_425),
	.V2C_1 (V2C_425_14),
	.V2C_2 (V2C_425_33),
	.V2C_3 (V2C_425_265),
	.V (V_425)
);

VNU_3 #(quan_width) VNU426 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_426),
	.C2V_2 (C2V_39_426),
	.C2V_3 (C2V_271_426),
	.L (L_426),
	.V2C_1 (V2C_426_20),
	.V2C_2 (V2C_426_39),
	.V2C_3 (V2C_426_271),
	.V (V_426)
);

VNU_3 #(quan_width) VNU427 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_427),
	.C2V_2 (C2V_45_427),
	.C2V_3 (C2V_277_427),
	.L (L_427),
	.V2C_1 (V2C_427_26),
	.V2C_2 (V2C_427_45),
	.V2C_3 (V2C_427_277),
	.V (V_427)
);

VNU_3 #(quan_width) VNU428 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_428),
	.C2V_2 (C2V_51_428),
	.C2V_3 (C2V_283_428),
	.L (L_428),
	.V2C_1 (V2C_428_32),
	.V2C_2 (V2C_428_51),
	.V2C_3 (V2C_428_283),
	.V (V_428)
);

VNU_3 #(quan_width) VNU429 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_429),
	.C2V_2 (C2V_38_429),
	.C2V_3 (C2V_57_429),
	.L (L_429),
	.V2C_1 (V2C_429_1),
	.V2C_2 (V2C_429_38),
	.V2C_3 (V2C_429_57),
	.V (V_429)
);

VNU_3 #(quan_width) VNU430 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_430),
	.C2V_2 (C2V_44_430),
	.C2V_3 (C2V_63_430),
	.L (L_430),
	.V2C_1 (V2C_430_7),
	.V2C_2 (V2C_430_44),
	.V2C_3 (V2C_430_63),
	.V (V_430)
);

VNU_3 #(quan_width) VNU431 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_431),
	.C2V_2 (C2V_50_431),
	.C2V_3 (C2V_69_431),
	.L (L_431),
	.V2C_1 (V2C_431_13),
	.V2C_2 (V2C_431_50),
	.V2C_3 (V2C_431_69),
	.V (V_431)
);

VNU_3 #(quan_width) VNU432 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_432),
	.C2V_2 (C2V_56_432),
	.C2V_3 (C2V_75_432),
	.L (L_432),
	.V2C_1 (V2C_432_19),
	.V2C_2 (V2C_432_56),
	.V2C_3 (V2C_432_75),
	.V (V_432)
);

VNU_3 #(quan_width) VNU433 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_433),
	.C2V_2 (C2V_28_433),
	.C2V_3 (C2V_251_433),
	.L (L_433),
	.V2C_1 (V2C_433_12),
	.V2C_2 (V2C_433_28),
	.V2C_3 (V2C_433_251),
	.V (V_433)
);

VNU_3 #(quan_width) VNU434 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_434),
	.C2V_2 (C2V_34_434),
	.C2V_3 (C2V_257_434),
	.L (L_434),
	.V2C_1 (V2C_434_18),
	.V2C_2 (V2C_434_34),
	.V2C_3 (V2C_434_257),
	.V (V_434)
);

VNU_3 #(quan_width) VNU435 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_435),
	.C2V_2 (C2V_40_435),
	.C2V_3 (C2V_263_435),
	.L (L_435),
	.V2C_1 (V2C_435_24),
	.V2C_2 (V2C_435_40),
	.V2C_3 (V2C_435_263),
	.V (V_435)
);

VNU_3 #(quan_width) VNU436 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_436),
	.C2V_2 (C2V_46_436),
	.C2V_3 (C2V_269_436),
	.L (L_436),
	.V2C_1 (V2C_436_30),
	.V2C_2 (V2C_436_46),
	.V2C_3 (V2C_436_269),
	.V (V_436)
);

VNU_3 #(quan_width) VNU437 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_437),
	.C2V_2 (C2V_52_437),
	.C2V_3 (C2V_275_437),
	.L (L_437),
	.V2C_1 (V2C_437_36),
	.V2C_2 (V2C_437_52),
	.V2C_3 (V2C_437_275),
	.V (V_437)
);

VNU_3 #(quan_width) VNU438 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_438),
	.C2V_2 (C2V_58_438),
	.C2V_3 (C2V_281_438),
	.L (L_438),
	.V2C_1 (V2C_438_42),
	.V2C_2 (V2C_438_58),
	.V2C_3 (V2C_438_281),
	.V (V_438)
);

VNU_3 #(quan_width) VNU439 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_439),
	.C2V_2 (C2V_64_439),
	.C2V_3 (C2V_287_439),
	.L (L_439),
	.V2C_1 (V2C_439_48),
	.V2C_2 (V2C_439_64),
	.V2C_3 (V2C_439_287),
	.V (V_439)
);

VNU_3 #(quan_width) VNU440 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_440),
	.C2V_2 (C2V_54_440),
	.C2V_3 (C2V_70_440),
	.L (L_440),
	.V2C_1 (V2C_440_5),
	.V2C_2 (V2C_440_54),
	.V2C_3 (V2C_440_70),
	.V (V_440)
);

VNU_3 #(quan_width) VNU441 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_441),
	.C2V_2 (C2V_60_441),
	.C2V_3 (C2V_76_441),
	.L (L_441),
	.V2C_1 (V2C_441_11),
	.V2C_2 (V2C_441_60),
	.V2C_3 (V2C_441_76),
	.V (V_441)
);

VNU_3 #(quan_width) VNU442 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_442),
	.C2V_2 (C2V_66_442),
	.C2V_3 (C2V_82_442),
	.L (L_442),
	.V2C_1 (V2C_442_17),
	.V2C_2 (V2C_442_66),
	.V2C_3 (V2C_442_82),
	.V (V_442)
);

VNU_3 #(quan_width) VNU443 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_443),
	.C2V_2 (C2V_72_443),
	.C2V_3 (C2V_88_443),
	.L (L_443),
	.V2C_1 (V2C_443_23),
	.V2C_2 (V2C_443_72),
	.V2C_3 (V2C_443_88),
	.V (V_443)
);

VNU_3 #(quan_width) VNU444 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_444),
	.C2V_2 (C2V_78_444),
	.C2V_3 (C2V_94_444),
	.L (L_444),
	.V2C_1 (V2C_444_29),
	.V2C_2 (V2C_444_78),
	.V2C_3 (V2C_444_94),
	.V (V_444)
);

VNU_3 #(quan_width) VNU445 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_445),
	.C2V_2 (C2V_84_445),
	.C2V_3 (C2V_100_445),
	.L (L_445),
	.V2C_1 (V2C_445_35),
	.V2C_2 (V2C_445_84),
	.V2C_3 (V2C_445_100),
	.V (V_445)
);

VNU_3 #(quan_width) VNU446 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_446),
	.C2V_2 (C2V_90_446),
	.C2V_3 (C2V_106_446),
	.L (L_446),
	.V2C_1 (V2C_446_41),
	.V2C_2 (V2C_446_90),
	.V2C_3 (V2C_446_106),
	.V (V_446)
);

VNU_3 #(quan_width) VNU447 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_447),
	.C2V_2 (C2V_96_447),
	.C2V_3 (C2V_112_447),
	.L (L_447),
	.V2C_1 (V2C_447_47),
	.V2C_2 (V2C_447_96),
	.V2C_3 (V2C_447_112),
	.V (V_447)
);

VNU_3 #(quan_width) VNU448 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_448),
	.C2V_2 (C2V_102_448),
	.C2V_3 (C2V_118_448),
	.L (L_448),
	.V2C_1 (V2C_448_53),
	.V2C_2 (V2C_448_102),
	.V2C_3 (V2C_448_118),
	.V (V_448)
);

VNU_3 #(quan_width) VNU449 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_59_449),
	.C2V_2 (C2V_108_449),
	.C2V_3 (C2V_124_449),
	.L (L_449),
	.V2C_1 (V2C_449_59),
	.V2C_2 (V2C_449_108),
	.V2C_3 (V2C_449_124),
	.V (V_449)
);

VNU_3 #(quan_width) VNU450 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_65_450),
	.C2V_2 (C2V_114_450),
	.C2V_3 (C2V_130_450),
	.L (L_450),
	.V2C_1 (V2C_450_65),
	.V2C_2 (V2C_450_114),
	.V2C_3 (V2C_450_130),
	.V (V_450)
);

VNU_3 #(quan_width) VNU451 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_71_451),
	.C2V_2 (C2V_120_451),
	.C2V_3 (C2V_136_451),
	.L (L_451),
	.V2C_1 (V2C_451_71),
	.V2C_2 (V2C_451_120),
	.V2C_3 (V2C_451_136),
	.V (V_451)
);

VNU_3 #(quan_width) VNU452 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_77_452),
	.C2V_2 (C2V_126_452),
	.C2V_3 (C2V_142_452),
	.L (L_452),
	.V2C_1 (V2C_452_77),
	.V2C_2 (V2C_452_126),
	.V2C_3 (V2C_452_142),
	.V (V_452)
);

VNU_3 #(quan_width) VNU453 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_83_453),
	.C2V_2 (C2V_132_453),
	.C2V_3 (C2V_148_453),
	.L (L_453),
	.V2C_1 (V2C_453_83),
	.V2C_2 (V2C_453_132),
	.V2C_3 (V2C_453_148),
	.V (V_453)
);

VNU_3 #(quan_width) VNU454 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_89_454),
	.C2V_2 (C2V_138_454),
	.C2V_3 (C2V_154_454),
	.L (L_454),
	.V2C_1 (V2C_454_89),
	.V2C_2 (V2C_454_138),
	.V2C_3 (V2C_454_154),
	.V (V_454)
);

VNU_3 #(quan_width) VNU455 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_95_455),
	.C2V_2 (C2V_144_455),
	.C2V_3 (C2V_160_455),
	.L (L_455),
	.V2C_1 (V2C_455_95),
	.V2C_2 (V2C_455_144),
	.V2C_3 (V2C_455_160),
	.V (V_455)
);

VNU_3 #(quan_width) VNU456 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_101_456),
	.C2V_2 (C2V_150_456),
	.C2V_3 (C2V_166_456),
	.L (L_456),
	.V2C_1 (V2C_456_101),
	.V2C_2 (V2C_456_150),
	.V2C_3 (V2C_456_166),
	.V (V_456)
);

VNU_3 #(quan_width) VNU457 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_107_457),
	.C2V_2 (C2V_156_457),
	.C2V_3 (C2V_172_457),
	.L (L_457),
	.V2C_1 (V2C_457_107),
	.V2C_2 (V2C_457_156),
	.V2C_3 (V2C_457_172),
	.V (V_457)
);

VNU_3 #(quan_width) VNU458 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_113_458),
	.C2V_2 (C2V_162_458),
	.C2V_3 (C2V_178_458),
	.L (L_458),
	.V2C_1 (V2C_458_113),
	.V2C_2 (V2C_458_162),
	.V2C_3 (V2C_458_178),
	.V (V_458)
);

VNU_3 #(quan_width) VNU459 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_119_459),
	.C2V_2 (C2V_168_459),
	.C2V_3 (C2V_184_459),
	.L (L_459),
	.V2C_1 (V2C_459_119),
	.V2C_2 (V2C_459_168),
	.V2C_3 (V2C_459_184),
	.V (V_459)
);

VNU_3 #(quan_width) VNU460 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_125_460),
	.C2V_2 (C2V_174_460),
	.C2V_3 (C2V_190_460),
	.L (L_460),
	.V2C_1 (V2C_460_125),
	.V2C_2 (V2C_460_174),
	.V2C_3 (V2C_460_190),
	.V (V_460)
);

VNU_3 #(quan_width) VNU461 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_131_461),
	.C2V_2 (C2V_180_461),
	.C2V_3 (C2V_196_461),
	.L (L_461),
	.V2C_1 (V2C_461_131),
	.V2C_2 (V2C_461_180),
	.V2C_3 (V2C_461_196),
	.V (V_461)
);

VNU_3 #(quan_width) VNU462 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_137_462),
	.C2V_2 (C2V_186_462),
	.C2V_3 (C2V_202_462),
	.L (L_462),
	.V2C_1 (V2C_462_137),
	.V2C_2 (V2C_462_186),
	.V2C_3 (V2C_462_202),
	.V (V_462)
);

VNU_3 #(quan_width) VNU463 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_143_463),
	.C2V_2 (C2V_192_463),
	.C2V_3 (C2V_208_463),
	.L (L_463),
	.V2C_1 (V2C_463_143),
	.V2C_2 (V2C_463_192),
	.V2C_3 (V2C_463_208),
	.V (V_463)
);

VNU_3 #(quan_width) VNU464 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_149_464),
	.C2V_2 (C2V_198_464),
	.C2V_3 (C2V_214_464),
	.L (L_464),
	.V2C_1 (V2C_464_149),
	.V2C_2 (V2C_464_198),
	.V2C_3 (V2C_464_214),
	.V (V_464)
);

VNU_3 #(quan_width) VNU465 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_155_465),
	.C2V_2 (C2V_204_465),
	.C2V_3 (C2V_220_465),
	.L (L_465),
	.V2C_1 (V2C_465_155),
	.V2C_2 (V2C_465_204),
	.V2C_3 (V2C_465_220),
	.V (V_465)
);

VNU_3 #(quan_width) VNU466 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_161_466),
	.C2V_2 (C2V_210_466),
	.C2V_3 (C2V_226_466),
	.L (L_466),
	.V2C_1 (V2C_466_161),
	.V2C_2 (V2C_466_210),
	.V2C_3 (V2C_466_226),
	.V (V_466)
);

VNU_3 #(quan_width) VNU467 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_167_467),
	.C2V_2 (C2V_216_467),
	.C2V_3 (C2V_232_467),
	.L (L_467),
	.V2C_1 (V2C_467_167),
	.V2C_2 (V2C_467_216),
	.V2C_3 (V2C_467_232),
	.V (V_467)
);

VNU_3 #(quan_width) VNU468 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_173_468),
	.C2V_2 (C2V_222_468),
	.C2V_3 (C2V_238_468),
	.L (L_468),
	.V2C_1 (V2C_468_173),
	.V2C_2 (V2C_468_222),
	.V2C_3 (V2C_468_238),
	.V (V_468)
);

VNU_3 #(quan_width) VNU469 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_179_469),
	.C2V_2 (C2V_228_469),
	.C2V_3 (C2V_244_469),
	.L (L_469),
	.V2C_1 (V2C_469_179),
	.V2C_2 (V2C_469_228),
	.V2C_3 (V2C_469_244),
	.V (V_469)
);

VNU_3 #(quan_width) VNU470 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_185_470),
	.C2V_2 (C2V_234_470),
	.C2V_3 (C2V_250_470),
	.L (L_470),
	.V2C_1 (V2C_470_185),
	.V2C_2 (V2C_470_234),
	.V2C_3 (V2C_470_250),
	.V (V_470)
);

VNU_3 #(quan_width) VNU471 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_191_471),
	.C2V_2 (C2V_240_471),
	.C2V_3 (C2V_256_471),
	.L (L_471),
	.V2C_1 (V2C_471_191),
	.V2C_2 (V2C_471_240),
	.V2C_3 (V2C_471_256),
	.V (V_471)
);

VNU_3 #(quan_width) VNU472 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_197_472),
	.C2V_2 (C2V_246_472),
	.C2V_3 (C2V_262_472),
	.L (L_472),
	.V2C_1 (V2C_472_197),
	.V2C_2 (V2C_472_246),
	.V2C_3 (V2C_472_262),
	.V (V_472)
);

VNU_3 #(quan_width) VNU473 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_203_473),
	.C2V_2 (C2V_252_473),
	.C2V_3 (C2V_268_473),
	.L (L_473),
	.V2C_1 (V2C_473_203),
	.V2C_2 (V2C_473_252),
	.V2C_3 (V2C_473_268),
	.V (V_473)
);

VNU_3 #(quan_width) VNU474 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_209_474),
	.C2V_2 (C2V_258_474),
	.C2V_3 (C2V_274_474),
	.L (L_474),
	.V2C_1 (V2C_474_209),
	.V2C_2 (V2C_474_258),
	.V2C_3 (V2C_474_274),
	.V (V_474)
);

VNU_3 #(quan_width) VNU475 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_215_475),
	.C2V_2 (C2V_264_475),
	.C2V_3 (C2V_280_475),
	.L (L_475),
	.V2C_1 (V2C_475_215),
	.V2C_2 (V2C_475_264),
	.V2C_3 (V2C_475_280),
	.V (V_475)
);

VNU_3 #(quan_width) VNU476 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_221_476),
	.C2V_2 (C2V_270_476),
	.C2V_3 (C2V_286_476),
	.L (L_476),
	.V2C_1 (V2C_476_221),
	.V2C_2 (V2C_476_270),
	.V2C_3 (V2C_476_286),
	.V (V_476)
);

VNU_3 #(quan_width) VNU477 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_477),
	.C2V_2 (C2V_227_477),
	.C2V_3 (C2V_276_477),
	.L (L_477),
	.V2C_1 (V2C_477_4),
	.V2C_2 (V2C_477_227),
	.V2C_3 (V2C_477_276),
	.V (V_477)
);

VNU_3 #(quan_width) VNU478 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_478),
	.C2V_2 (C2V_233_478),
	.C2V_3 (C2V_282_478),
	.L (L_478),
	.V2C_1 (V2C_478_10),
	.V2C_2 (V2C_478_233),
	.V2C_3 (V2C_478_282),
	.V (V_478)
);

VNU_3 #(quan_width) VNU479 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_479),
	.C2V_2 (C2V_239_479),
	.C2V_3 (C2V_288_479),
	.L (L_479),
	.V2C_1 (V2C_479_16),
	.V2C_2 (V2C_479_239),
	.V2C_3 (V2C_479_288),
	.V (V_479)
);

VNU_3 #(quan_width) VNU480 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_480),
	.C2V_2 (C2V_22_480),
	.C2V_3 (C2V_245_480),
	.L (L_480),
	.V2C_1 (V2C_480_6),
	.V2C_2 (V2C_480_22),
	.V2C_3 (V2C_480_245),
	.V (V_480)
);

VNU_3 #(quan_width) VNU481 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_481),
	.C2V_2 (C2V_76_481),
	.C2V_3 (C2V_104_481),
	.L (L_481),
	.V2C_1 (V2C_481_19),
	.V2C_2 (V2C_481_76),
	.V2C_3 (V2C_481_104),
	.V (V_481)
);

VNU_3 #(quan_width) VNU482 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_482),
	.C2V_2 (C2V_82_482),
	.C2V_3 (C2V_110_482),
	.L (L_482),
	.V2C_1 (V2C_482_25),
	.V2C_2 (V2C_482_82),
	.V2C_3 (V2C_482_110),
	.V (V_482)
);

VNU_3 #(quan_width) VNU483 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_483),
	.C2V_2 (C2V_88_483),
	.C2V_3 (C2V_116_483),
	.L (L_483),
	.V2C_1 (V2C_483_31),
	.V2C_2 (V2C_483_88),
	.V2C_3 (V2C_483_116),
	.V (V_483)
);

VNU_3 #(quan_width) VNU484 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_484),
	.C2V_2 (C2V_94_484),
	.C2V_3 (C2V_122_484),
	.L (L_484),
	.V2C_1 (V2C_484_37),
	.V2C_2 (V2C_484_94),
	.V2C_3 (V2C_484_122),
	.V (V_484)
);

VNU_3 #(quan_width) VNU485 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_485),
	.C2V_2 (C2V_100_485),
	.C2V_3 (C2V_128_485),
	.L (L_485),
	.V2C_1 (V2C_485_43),
	.V2C_2 (V2C_485_100),
	.V2C_3 (V2C_485_128),
	.V (V_485)
);

VNU_3 #(quan_width) VNU486 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_486),
	.C2V_2 (C2V_106_486),
	.C2V_3 (C2V_134_486),
	.L (L_486),
	.V2C_1 (V2C_486_49),
	.V2C_2 (V2C_486_106),
	.V2C_3 (V2C_486_134),
	.V (V_486)
);

VNU_3 #(quan_width) VNU487 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_487),
	.C2V_2 (C2V_112_487),
	.C2V_3 (C2V_140_487),
	.L (L_487),
	.V2C_1 (V2C_487_55),
	.V2C_2 (V2C_487_112),
	.V2C_3 (V2C_487_140),
	.V (V_487)
);

VNU_3 #(quan_width) VNU488 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_488),
	.C2V_2 (C2V_118_488),
	.C2V_3 (C2V_146_488),
	.L (L_488),
	.V2C_1 (V2C_488_61),
	.V2C_2 (V2C_488_118),
	.V2C_3 (V2C_488_146),
	.V (V_488)
);

VNU_3 #(quan_width) VNU489 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_489),
	.C2V_2 (C2V_124_489),
	.C2V_3 (C2V_152_489),
	.L (L_489),
	.V2C_1 (V2C_489_67),
	.V2C_2 (V2C_489_124),
	.V2C_3 (V2C_489_152),
	.V (V_489)
);

VNU_3 #(quan_width) VNU490 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_490),
	.C2V_2 (C2V_130_490),
	.C2V_3 (C2V_158_490),
	.L (L_490),
	.V2C_1 (V2C_490_73),
	.V2C_2 (V2C_490_130),
	.V2C_3 (V2C_490_158),
	.V (V_490)
);

VNU_3 #(quan_width) VNU491 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_491),
	.C2V_2 (C2V_136_491),
	.C2V_3 (C2V_164_491),
	.L (L_491),
	.V2C_1 (V2C_491_79),
	.V2C_2 (V2C_491_136),
	.V2C_3 (V2C_491_164),
	.V (V_491)
);

VNU_3 #(quan_width) VNU492 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_492),
	.C2V_2 (C2V_142_492),
	.C2V_3 (C2V_170_492),
	.L (L_492),
	.V2C_1 (V2C_492_85),
	.V2C_2 (V2C_492_142),
	.V2C_3 (V2C_492_170),
	.V (V_492)
);

VNU_3 #(quan_width) VNU493 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_91_493),
	.C2V_2 (C2V_148_493),
	.C2V_3 (C2V_176_493),
	.L (L_493),
	.V2C_1 (V2C_493_91),
	.V2C_2 (V2C_493_148),
	.V2C_3 (V2C_493_176),
	.V (V_493)
);

VNU_3 #(quan_width) VNU494 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_97_494),
	.C2V_2 (C2V_154_494),
	.C2V_3 (C2V_182_494),
	.L (L_494),
	.V2C_1 (V2C_494_97),
	.V2C_2 (V2C_494_154),
	.V2C_3 (V2C_494_182),
	.V (V_494)
);

VNU_3 #(quan_width) VNU495 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_103_495),
	.C2V_2 (C2V_160_495),
	.C2V_3 (C2V_188_495),
	.L (L_495),
	.V2C_1 (V2C_495_103),
	.V2C_2 (V2C_495_160),
	.V2C_3 (V2C_495_188),
	.V (V_495)
);

VNU_3 #(quan_width) VNU496 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_109_496),
	.C2V_2 (C2V_166_496),
	.C2V_3 (C2V_194_496),
	.L (L_496),
	.V2C_1 (V2C_496_109),
	.V2C_2 (V2C_496_166),
	.V2C_3 (V2C_496_194),
	.V (V_496)
);

VNU_3 #(quan_width) VNU497 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_115_497),
	.C2V_2 (C2V_172_497),
	.C2V_3 (C2V_200_497),
	.L (L_497),
	.V2C_1 (V2C_497_115),
	.V2C_2 (V2C_497_172),
	.V2C_3 (V2C_497_200),
	.V (V_497)
);

VNU_3 #(quan_width) VNU498 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_121_498),
	.C2V_2 (C2V_178_498),
	.C2V_3 (C2V_206_498),
	.L (L_498),
	.V2C_1 (V2C_498_121),
	.V2C_2 (V2C_498_178),
	.V2C_3 (V2C_498_206),
	.V (V_498)
);

VNU_3 #(quan_width) VNU499 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_127_499),
	.C2V_2 (C2V_184_499),
	.C2V_3 (C2V_212_499),
	.L (L_499),
	.V2C_1 (V2C_499_127),
	.V2C_2 (V2C_499_184),
	.V2C_3 (V2C_499_212),
	.V (V_499)
);

VNU_3 #(quan_width) VNU500 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_133_500),
	.C2V_2 (C2V_190_500),
	.C2V_3 (C2V_218_500),
	.L (L_500),
	.V2C_1 (V2C_500_133),
	.V2C_2 (V2C_500_190),
	.V2C_3 (V2C_500_218),
	.V (V_500)
);

VNU_3 #(quan_width) VNU501 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_139_501),
	.C2V_2 (C2V_196_501),
	.C2V_3 (C2V_224_501),
	.L (L_501),
	.V2C_1 (V2C_501_139),
	.V2C_2 (V2C_501_196),
	.V2C_3 (V2C_501_224),
	.V (V_501)
);

VNU_3 #(quan_width) VNU502 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_145_502),
	.C2V_2 (C2V_202_502),
	.C2V_3 (C2V_230_502),
	.L (L_502),
	.V2C_1 (V2C_502_145),
	.V2C_2 (V2C_502_202),
	.V2C_3 (V2C_502_230),
	.V (V_502)
);

VNU_3 #(quan_width) VNU503 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_151_503),
	.C2V_2 (C2V_208_503),
	.C2V_3 (C2V_236_503),
	.L (L_503),
	.V2C_1 (V2C_503_151),
	.V2C_2 (V2C_503_208),
	.V2C_3 (V2C_503_236),
	.V (V_503)
);

VNU_3 #(quan_width) VNU504 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_157_504),
	.C2V_2 (C2V_214_504),
	.C2V_3 (C2V_242_504),
	.L (L_504),
	.V2C_1 (V2C_504_157),
	.V2C_2 (V2C_504_214),
	.V2C_3 (V2C_504_242),
	.V (V_504)
);

VNU_3 #(quan_width) VNU505 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_163_505),
	.C2V_2 (C2V_220_505),
	.C2V_3 (C2V_248_505),
	.L (L_505),
	.V2C_1 (V2C_505_163),
	.V2C_2 (V2C_505_220),
	.V2C_3 (V2C_505_248),
	.V (V_505)
);

VNU_3 #(quan_width) VNU506 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_169_506),
	.C2V_2 (C2V_226_506),
	.C2V_3 (C2V_254_506),
	.L (L_506),
	.V2C_1 (V2C_506_169),
	.V2C_2 (V2C_506_226),
	.V2C_3 (V2C_506_254),
	.V (V_506)
);

VNU_3 #(quan_width) VNU507 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_175_507),
	.C2V_2 (C2V_232_507),
	.C2V_3 (C2V_260_507),
	.L (L_507),
	.V2C_1 (V2C_507_175),
	.V2C_2 (V2C_507_232),
	.V2C_3 (V2C_507_260),
	.V (V_507)
);

VNU_3 #(quan_width) VNU508 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_181_508),
	.C2V_2 (C2V_238_508),
	.C2V_3 (C2V_266_508),
	.L (L_508),
	.V2C_1 (V2C_508_181),
	.V2C_2 (V2C_508_238),
	.V2C_3 (V2C_508_266),
	.V (V_508)
);

VNU_3 #(quan_width) VNU509 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_187_509),
	.C2V_2 (C2V_244_509),
	.C2V_3 (C2V_272_509),
	.L (L_509),
	.V2C_1 (V2C_509_187),
	.V2C_2 (V2C_509_244),
	.V2C_3 (V2C_509_272),
	.V (V_509)
);

VNU_3 #(quan_width) VNU510 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_193_510),
	.C2V_2 (C2V_250_510),
	.C2V_3 (C2V_278_510),
	.L (L_510),
	.V2C_1 (V2C_510_193),
	.V2C_2 (V2C_510_250),
	.V2C_3 (V2C_510_278),
	.V (V_510)
);

VNU_3 #(quan_width) VNU511 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_199_511),
	.C2V_2 (C2V_256_511),
	.C2V_3 (C2V_284_511),
	.L (L_511),
	.V2C_1 (V2C_511_199),
	.V2C_2 (V2C_511_256),
	.V2C_3 (V2C_511_284),
	.V (V_511)
);

VNU_3 #(quan_width) VNU512 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_512),
	.C2V_2 (C2V_205_512),
	.C2V_3 (C2V_262_512),
	.L (L_512),
	.V2C_1 (V2C_512_2),
	.V2C_2 (V2C_512_205),
	.V2C_3 (V2C_512_262),
	.V (V_512)
);

VNU_3 #(quan_width) VNU513 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_513),
	.C2V_2 (C2V_211_513),
	.C2V_3 (C2V_268_513),
	.L (L_513),
	.V2C_1 (V2C_513_8),
	.V2C_2 (V2C_513_211),
	.V2C_3 (V2C_513_268),
	.V (V_513)
);

VNU_3 #(quan_width) VNU514 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_514),
	.C2V_2 (C2V_217_514),
	.C2V_3 (C2V_274_514),
	.L (L_514),
	.V2C_1 (V2C_514_14),
	.V2C_2 (V2C_514_217),
	.V2C_3 (V2C_514_274),
	.V (V_514)
);

VNU_3 #(quan_width) VNU515 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_515),
	.C2V_2 (C2V_223_515),
	.C2V_3 (C2V_280_515),
	.L (L_515),
	.V2C_1 (V2C_515_20),
	.V2C_2 (V2C_515_223),
	.V2C_3 (V2C_515_280),
	.V (V_515)
);

VNU_3 #(quan_width) VNU516 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_516),
	.C2V_2 (C2V_229_516),
	.C2V_3 (C2V_286_516),
	.L (L_516),
	.V2C_1 (V2C_516_26),
	.V2C_2 (V2C_516_229),
	.V2C_3 (V2C_516_286),
	.V (V_516)
);

VNU_3 #(quan_width) VNU517 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_517),
	.C2V_2 (C2V_32_517),
	.C2V_3 (C2V_235_517),
	.L (L_517),
	.V2C_1 (V2C_517_4),
	.V2C_2 (V2C_517_32),
	.V2C_3 (V2C_517_235),
	.V (V_517)
);

VNU_3 #(quan_width) VNU518 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_518),
	.C2V_2 (C2V_38_518),
	.C2V_3 (C2V_241_518),
	.L (L_518),
	.V2C_1 (V2C_518_10),
	.V2C_2 (V2C_518_38),
	.V2C_3 (V2C_518_241),
	.V (V_518)
);

VNU_3 #(quan_width) VNU519 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_519),
	.C2V_2 (C2V_44_519),
	.C2V_3 (C2V_247_519),
	.L (L_519),
	.V2C_1 (V2C_519_16),
	.V2C_2 (V2C_519_44),
	.V2C_3 (V2C_519_247),
	.V (V_519)
);

VNU_3 #(quan_width) VNU520 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_520),
	.C2V_2 (C2V_50_520),
	.C2V_3 (C2V_253_520),
	.L (L_520),
	.V2C_1 (V2C_520_22),
	.V2C_2 (V2C_520_50),
	.V2C_3 (V2C_520_253),
	.V (V_520)
);

VNU_3 #(quan_width) VNU521 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_521),
	.C2V_2 (C2V_56_521),
	.C2V_3 (C2V_259_521),
	.L (L_521),
	.V2C_1 (V2C_521_28),
	.V2C_2 (V2C_521_56),
	.V2C_3 (V2C_521_259),
	.V (V_521)
);

VNU_3 #(quan_width) VNU522 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_522),
	.C2V_2 (C2V_62_522),
	.C2V_3 (C2V_265_522),
	.L (L_522),
	.V2C_1 (V2C_522_34),
	.V2C_2 (V2C_522_62),
	.V2C_3 (V2C_522_265),
	.V (V_522)
);

VNU_3 #(quan_width) VNU523 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_523),
	.C2V_2 (C2V_68_523),
	.C2V_3 (C2V_271_523),
	.L (L_523),
	.V2C_1 (V2C_523_40),
	.V2C_2 (V2C_523_68),
	.V2C_3 (V2C_523_271),
	.V (V_523)
);

VNU_3 #(quan_width) VNU524 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_524),
	.C2V_2 (C2V_74_524),
	.C2V_3 (C2V_277_524),
	.L (L_524),
	.V2C_1 (V2C_524_46),
	.V2C_2 (V2C_524_74),
	.V2C_3 (V2C_524_277),
	.V (V_524)
);

VNU_3 #(quan_width) VNU525 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_525),
	.C2V_2 (C2V_80_525),
	.C2V_3 (C2V_283_525),
	.L (L_525),
	.V2C_1 (V2C_525_52),
	.V2C_2 (V2C_525_80),
	.V2C_3 (V2C_525_283),
	.V (V_525)
);

VNU_3 #(quan_width) VNU526 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_526),
	.C2V_2 (C2V_58_526),
	.C2V_3 (C2V_86_526),
	.L (L_526),
	.V2C_1 (V2C_526_1),
	.V2C_2 (V2C_526_58),
	.V2C_3 (V2C_526_86),
	.V (V_526)
);

VNU_3 #(quan_width) VNU527 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_527),
	.C2V_2 (C2V_64_527),
	.C2V_3 (C2V_92_527),
	.L (L_527),
	.V2C_1 (V2C_527_7),
	.V2C_2 (V2C_527_64),
	.V2C_3 (V2C_527_92),
	.V (V_527)
);

VNU_3 #(quan_width) VNU528 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_528),
	.C2V_2 (C2V_70_528),
	.C2V_3 (C2V_98_528),
	.L (L_528),
	.V2C_1 (V2C_528_13),
	.V2C_2 (V2C_528_70),
	.V2C_3 (V2C_528_98),
	.V (V_528)
);

VNU_3 #(quan_width) VNU529 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_529),
	.C2V_2 (C2V_148_529),
	.C2V_3 (C2V_279_529),
	.L (L_529),
	.V2C_1 (V2C_529_6),
	.V2C_2 (V2C_529_148),
	.V2C_3 (V2C_529_279),
	.V (V_529)
);

VNU_3 #(quan_width) VNU530 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_530),
	.C2V_2 (C2V_154_530),
	.C2V_3 (C2V_285_530),
	.L (L_530),
	.V2C_1 (V2C_530_12),
	.V2C_2 (V2C_530_154),
	.V2C_3 (V2C_530_285),
	.V (V_530)
);

VNU_3 #(quan_width) VNU531 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_531),
	.C2V_2 (C2V_18_531),
	.C2V_3 (C2V_160_531),
	.L (L_531),
	.V2C_1 (V2C_531_3),
	.V2C_2 (V2C_531_18),
	.V2C_3 (V2C_531_160),
	.V (V_531)
);

VNU_3 #(quan_width) VNU532 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_532),
	.C2V_2 (C2V_24_532),
	.C2V_3 (C2V_166_532),
	.L (L_532),
	.V2C_1 (V2C_532_9),
	.V2C_2 (V2C_532_24),
	.V2C_3 (V2C_532_166),
	.V (V_532)
);

VNU_3 #(quan_width) VNU533 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_533),
	.C2V_2 (C2V_30_533),
	.C2V_3 (C2V_172_533),
	.L (L_533),
	.V2C_1 (V2C_533_15),
	.V2C_2 (V2C_533_30),
	.V2C_3 (V2C_533_172),
	.V (V_533)
);

VNU_3 #(quan_width) VNU534 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_534),
	.C2V_2 (C2V_36_534),
	.C2V_3 (C2V_178_534),
	.L (L_534),
	.V2C_1 (V2C_534_21),
	.V2C_2 (V2C_534_36),
	.V2C_3 (V2C_534_178),
	.V (V_534)
);

VNU_3 #(quan_width) VNU535 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_535),
	.C2V_2 (C2V_42_535),
	.C2V_3 (C2V_184_535),
	.L (L_535),
	.V2C_1 (V2C_535_27),
	.V2C_2 (V2C_535_42),
	.V2C_3 (V2C_535_184),
	.V (V_535)
);

VNU_3 #(quan_width) VNU536 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_536),
	.C2V_2 (C2V_48_536),
	.C2V_3 (C2V_190_536),
	.L (L_536),
	.V2C_1 (V2C_536_33),
	.V2C_2 (V2C_536_48),
	.V2C_3 (V2C_536_190),
	.V (V_536)
);

VNU_3 #(quan_width) VNU537 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_537),
	.C2V_2 (C2V_54_537),
	.C2V_3 (C2V_196_537),
	.L (L_537),
	.V2C_1 (V2C_537_39),
	.V2C_2 (V2C_537_54),
	.V2C_3 (V2C_537_196),
	.V (V_537)
);

VNU_3 #(quan_width) VNU538 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_538),
	.C2V_2 (C2V_60_538),
	.C2V_3 (C2V_202_538),
	.L (L_538),
	.V2C_1 (V2C_538_45),
	.V2C_2 (V2C_538_60),
	.V2C_3 (V2C_538_202),
	.V (V_538)
);

VNU_3 #(quan_width) VNU539 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_539),
	.C2V_2 (C2V_66_539),
	.C2V_3 (C2V_208_539),
	.L (L_539),
	.V2C_1 (V2C_539_51),
	.V2C_2 (V2C_539_66),
	.V2C_3 (V2C_539_208),
	.V (V_539)
);

VNU_3 #(quan_width) VNU540 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_540),
	.C2V_2 (C2V_72_540),
	.C2V_3 (C2V_214_540),
	.L (L_540),
	.V2C_1 (V2C_540_57),
	.V2C_2 (V2C_540_72),
	.V2C_3 (V2C_540_214),
	.V (V_540)
);

VNU_3 #(quan_width) VNU541 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_541),
	.C2V_2 (C2V_78_541),
	.C2V_3 (C2V_220_541),
	.L (L_541),
	.V2C_1 (V2C_541_63),
	.V2C_2 (V2C_541_78),
	.V2C_3 (V2C_541_220),
	.V (V_541)
);

VNU_3 #(quan_width) VNU542 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_542),
	.C2V_2 (C2V_84_542),
	.C2V_3 (C2V_226_542),
	.L (L_542),
	.V2C_1 (V2C_542_69),
	.V2C_2 (V2C_542_84),
	.V2C_3 (V2C_542_226),
	.V (V_542)
);

VNU_3 #(quan_width) VNU543 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_543),
	.C2V_2 (C2V_90_543),
	.C2V_3 (C2V_232_543),
	.L (L_543),
	.V2C_1 (V2C_543_75),
	.V2C_2 (V2C_543_90),
	.V2C_3 (V2C_543_232),
	.V (V_543)
);

VNU_3 #(quan_width) VNU544 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_544),
	.C2V_2 (C2V_96_544),
	.C2V_3 (C2V_238_544),
	.L (L_544),
	.V2C_1 (V2C_544_81),
	.V2C_2 (V2C_544_96),
	.V2C_3 (V2C_544_238),
	.V (V_544)
);

VNU_3 #(quan_width) VNU545 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_545),
	.C2V_2 (C2V_102_545),
	.C2V_3 (C2V_244_545),
	.L (L_545),
	.V2C_1 (V2C_545_87),
	.V2C_2 (V2C_545_102),
	.V2C_3 (V2C_545_244),
	.V (V_545)
);

VNU_3 #(quan_width) VNU546 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_93_546),
	.C2V_2 (C2V_108_546),
	.C2V_3 (C2V_250_546),
	.L (L_546),
	.V2C_1 (V2C_546_93),
	.V2C_2 (V2C_546_108),
	.V2C_3 (V2C_546_250),
	.V (V_546)
);

VNU_3 #(quan_width) VNU547 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_99_547),
	.C2V_2 (C2V_114_547),
	.C2V_3 (C2V_256_547),
	.L (L_547),
	.V2C_1 (V2C_547_99),
	.V2C_2 (V2C_547_114),
	.V2C_3 (V2C_547_256),
	.V (V_547)
);

VNU_3 #(quan_width) VNU548 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_105_548),
	.C2V_2 (C2V_120_548),
	.C2V_3 (C2V_262_548),
	.L (L_548),
	.V2C_1 (V2C_548_105),
	.V2C_2 (V2C_548_120),
	.V2C_3 (V2C_548_262),
	.V (V_548)
);

VNU_3 #(quan_width) VNU549 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_111_549),
	.C2V_2 (C2V_126_549),
	.C2V_3 (C2V_268_549),
	.L (L_549),
	.V2C_1 (V2C_549_111),
	.V2C_2 (V2C_549_126),
	.V2C_3 (V2C_549_268),
	.V (V_549)
);

VNU_3 #(quan_width) VNU550 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_117_550),
	.C2V_2 (C2V_132_550),
	.C2V_3 (C2V_274_550),
	.L (L_550),
	.V2C_1 (V2C_550_117),
	.V2C_2 (V2C_550_132),
	.V2C_3 (V2C_550_274),
	.V (V_550)
);

VNU_3 #(quan_width) VNU551 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_123_551),
	.C2V_2 (C2V_138_551),
	.C2V_3 (C2V_280_551),
	.L (L_551),
	.V2C_1 (V2C_551_123),
	.V2C_2 (V2C_551_138),
	.V2C_3 (V2C_551_280),
	.V (V_551)
);

VNU_3 #(quan_width) VNU552 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_129_552),
	.C2V_2 (C2V_144_552),
	.C2V_3 (C2V_286_552),
	.L (L_552),
	.V2C_1 (V2C_552_129),
	.V2C_2 (V2C_552_144),
	.V2C_3 (V2C_552_286),
	.V (V_552)
);

VNU_3 #(quan_width) VNU553 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_553),
	.C2V_2 (C2V_135_553),
	.C2V_3 (C2V_150_553),
	.L (L_553),
	.V2C_1 (V2C_553_4),
	.V2C_2 (V2C_553_135),
	.V2C_3 (V2C_553_150),
	.V (V_553)
);

VNU_3 #(quan_width) VNU554 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_554),
	.C2V_2 (C2V_141_554),
	.C2V_3 (C2V_156_554),
	.L (L_554),
	.V2C_1 (V2C_554_10),
	.V2C_2 (V2C_554_141),
	.V2C_3 (V2C_554_156),
	.V (V_554)
);

VNU_3 #(quan_width) VNU555 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_555),
	.C2V_2 (C2V_147_555),
	.C2V_3 (C2V_162_555),
	.L (L_555),
	.V2C_1 (V2C_555_16),
	.V2C_2 (V2C_555_147),
	.V2C_3 (V2C_555_162),
	.V (V_555)
);

VNU_3 #(quan_width) VNU556 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_556),
	.C2V_2 (C2V_153_556),
	.C2V_3 (C2V_168_556),
	.L (L_556),
	.V2C_1 (V2C_556_22),
	.V2C_2 (V2C_556_153),
	.V2C_3 (V2C_556_168),
	.V (V_556)
);

VNU_3 #(quan_width) VNU557 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_557),
	.C2V_2 (C2V_159_557),
	.C2V_3 (C2V_174_557),
	.L (L_557),
	.V2C_1 (V2C_557_28),
	.V2C_2 (V2C_557_159),
	.V2C_3 (V2C_557_174),
	.V (V_557)
);

VNU_3 #(quan_width) VNU558 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_558),
	.C2V_2 (C2V_165_558),
	.C2V_3 (C2V_180_558),
	.L (L_558),
	.V2C_1 (V2C_558_34),
	.V2C_2 (V2C_558_165),
	.V2C_3 (V2C_558_180),
	.V (V_558)
);

VNU_3 #(quan_width) VNU559 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_559),
	.C2V_2 (C2V_171_559),
	.C2V_3 (C2V_186_559),
	.L (L_559),
	.V2C_1 (V2C_559_40),
	.V2C_2 (V2C_559_171),
	.V2C_3 (V2C_559_186),
	.V (V_559)
);

VNU_3 #(quan_width) VNU560 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_560),
	.C2V_2 (C2V_177_560),
	.C2V_3 (C2V_192_560),
	.L (L_560),
	.V2C_1 (V2C_560_46),
	.V2C_2 (V2C_560_177),
	.V2C_3 (V2C_560_192),
	.V (V_560)
);

VNU_3 #(quan_width) VNU561 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_561),
	.C2V_2 (C2V_183_561),
	.C2V_3 (C2V_198_561),
	.L (L_561),
	.V2C_1 (V2C_561_52),
	.V2C_2 (V2C_561_183),
	.V2C_3 (V2C_561_198),
	.V (V_561)
);

VNU_3 #(quan_width) VNU562 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_562),
	.C2V_2 (C2V_189_562),
	.C2V_3 (C2V_204_562),
	.L (L_562),
	.V2C_1 (V2C_562_58),
	.V2C_2 (V2C_562_189),
	.V2C_3 (V2C_562_204),
	.V (V_562)
);

VNU_3 #(quan_width) VNU563 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_563),
	.C2V_2 (C2V_195_563),
	.C2V_3 (C2V_210_563),
	.L (L_563),
	.V2C_1 (V2C_563_64),
	.V2C_2 (V2C_563_195),
	.V2C_3 (V2C_563_210),
	.V (V_563)
);

VNU_3 #(quan_width) VNU564 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_564),
	.C2V_2 (C2V_201_564),
	.C2V_3 (C2V_216_564),
	.L (L_564),
	.V2C_1 (V2C_564_70),
	.V2C_2 (V2C_564_201),
	.V2C_3 (V2C_564_216),
	.V (V_564)
);

VNU_3 #(quan_width) VNU565 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_565),
	.C2V_2 (C2V_207_565),
	.C2V_3 (C2V_222_565),
	.L (L_565),
	.V2C_1 (V2C_565_76),
	.V2C_2 (V2C_565_207),
	.V2C_3 (V2C_565_222),
	.V (V_565)
);

VNU_3 #(quan_width) VNU566 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_566),
	.C2V_2 (C2V_213_566),
	.C2V_3 (C2V_228_566),
	.L (L_566),
	.V2C_1 (V2C_566_82),
	.V2C_2 (V2C_566_213),
	.V2C_3 (V2C_566_228),
	.V (V_566)
);

VNU_3 #(quan_width) VNU567 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_567),
	.C2V_2 (C2V_219_567),
	.C2V_3 (C2V_234_567),
	.L (L_567),
	.V2C_1 (V2C_567_88),
	.V2C_2 (V2C_567_219),
	.V2C_3 (V2C_567_234),
	.V (V_567)
);

VNU_3 #(quan_width) VNU568 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_568),
	.C2V_2 (C2V_225_568),
	.C2V_3 (C2V_240_568),
	.L (L_568),
	.V2C_1 (V2C_568_94),
	.V2C_2 (V2C_568_225),
	.V2C_3 (V2C_568_240),
	.V (V_568)
);

VNU_3 #(quan_width) VNU569 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_569),
	.C2V_2 (C2V_231_569),
	.C2V_3 (C2V_246_569),
	.L (L_569),
	.V2C_1 (V2C_569_100),
	.V2C_2 (V2C_569_231),
	.V2C_3 (V2C_569_246),
	.V (V_569)
);

VNU_3 #(quan_width) VNU570 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_570),
	.C2V_2 (C2V_237_570),
	.C2V_3 (C2V_252_570),
	.L (L_570),
	.V2C_1 (V2C_570_106),
	.V2C_2 (V2C_570_237),
	.V2C_3 (V2C_570_252),
	.V (V_570)
);

VNU_3 #(quan_width) VNU571 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_571),
	.C2V_2 (C2V_243_571),
	.C2V_3 (C2V_258_571),
	.L (L_571),
	.V2C_1 (V2C_571_112),
	.V2C_2 (V2C_571_243),
	.V2C_3 (V2C_571_258),
	.V (V_571)
);

VNU_3 #(quan_width) VNU572 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_118_572),
	.C2V_2 (C2V_249_572),
	.C2V_3 (C2V_264_572),
	.L (L_572),
	.V2C_1 (V2C_572_118),
	.V2C_2 (V2C_572_249),
	.V2C_3 (V2C_572_264),
	.V (V_572)
);

VNU_3 #(quan_width) VNU573 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_124_573),
	.C2V_2 (C2V_255_573),
	.C2V_3 (C2V_270_573),
	.L (L_573),
	.V2C_1 (V2C_573_124),
	.V2C_2 (V2C_573_255),
	.V2C_3 (V2C_573_270),
	.V (V_573)
);

VNU_3 #(quan_width) VNU574 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_130_574),
	.C2V_2 (C2V_261_574),
	.C2V_3 (C2V_276_574),
	.L (L_574),
	.V2C_1 (V2C_574_130),
	.V2C_2 (V2C_574_261),
	.V2C_3 (V2C_574_276),
	.V (V_574)
);

VNU_3 #(quan_width) VNU575 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_136_575),
	.C2V_2 (C2V_267_575),
	.C2V_3 (C2V_282_575),
	.L (L_575),
	.V2C_1 (V2C_575_136),
	.V2C_2 (V2C_575_267),
	.V2C_3 (V2C_575_282),
	.V (V_575)
);

VNU_3 #(quan_width) VNU576 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_142_576),
	.C2V_2 (C2V_273_576),
	.C2V_3 (C2V_288_576),
	.L (L_576),
	.V2C_1 (V2C_576_142),
	.V2C_2 (V2C_576_273),
	.V2C_3 (V2C_576_288),
	.V (V_576)
);

VNU_3 #(quan_width) VNU577 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_577),
	.C2V_2 (C2V_96_577),
	.C2V_3 (C2V_225_577),
	.L (L_577),
	.V2C_1 (V2C_577_64),
	.V2C_2 (V2C_577_96),
	.V2C_3 (V2C_577_225),
	.V (V_577)
);

VNU_3 #(quan_width) VNU578 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_578),
	.C2V_2 (C2V_102_578),
	.C2V_3 (C2V_231_578),
	.L (L_578),
	.V2C_1 (V2C_578_70),
	.V2C_2 (V2C_578_102),
	.V2C_3 (V2C_578_231),
	.V (V_578)
);

VNU_3 #(quan_width) VNU579 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_579),
	.C2V_2 (C2V_108_579),
	.C2V_3 (C2V_237_579),
	.L (L_579),
	.V2C_1 (V2C_579_76),
	.V2C_2 (V2C_579_108),
	.V2C_3 (V2C_579_237),
	.V (V_579)
);

VNU_3 #(quan_width) VNU580 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_580),
	.C2V_2 (C2V_114_580),
	.C2V_3 (C2V_243_580),
	.L (L_580),
	.V2C_1 (V2C_580_82),
	.V2C_2 (V2C_580_114),
	.V2C_3 (V2C_580_243),
	.V (V_580)
);

VNU_3 #(quan_width) VNU581 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_581),
	.C2V_2 (C2V_120_581),
	.C2V_3 (C2V_249_581),
	.L (L_581),
	.V2C_1 (V2C_581_88),
	.V2C_2 (V2C_581_120),
	.V2C_3 (V2C_581_249),
	.V (V_581)
);

VNU_3 #(quan_width) VNU582 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_582),
	.C2V_2 (C2V_126_582),
	.C2V_3 (C2V_255_582),
	.L (L_582),
	.V2C_1 (V2C_582_94),
	.V2C_2 (V2C_582_126),
	.V2C_3 (V2C_582_255),
	.V (V_582)
);

VNU_3 #(quan_width) VNU583 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_583),
	.C2V_2 (C2V_132_583),
	.C2V_3 (C2V_261_583),
	.L (L_583),
	.V2C_1 (V2C_583_100),
	.V2C_2 (V2C_583_132),
	.V2C_3 (V2C_583_261),
	.V (V_583)
);

VNU_3 #(quan_width) VNU584 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_584),
	.C2V_2 (C2V_138_584),
	.C2V_3 (C2V_267_584),
	.L (L_584),
	.V2C_1 (V2C_584_106),
	.V2C_2 (V2C_584_138),
	.V2C_3 (V2C_584_267),
	.V (V_584)
);

VNU_3 #(quan_width) VNU585 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_585),
	.C2V_2 (C2V_144_585),
	.C2V_3 (C2V_273_585),
	.L (L_585),
	.V2C_1 (V2C_585_112),
	.V2C_2 (V2C_585_144),
	.V2C_3 (V2C_585_273),
	.V (V_585)
);

VNU_3 #(quan_width) VNU586 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_118_586),
	.C2V_2 (C2V_150_586),
	.C2V_3 (C2V_279_586),
	.L (L_586),
	.V2C_1 (V2C_586_118),
	.V2C_2 (V2C_586_150),
	.V2C_3 (V2C_586_279),
	.V (V_586)
);

VNU_3 #(quan_width) VNU587 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_124_587),
	.C2V_2 (C2V_156_587),
	.C2V_3 (C2V_285_587),
	.L (L_587),
	.V2C_1 (V2C_587_124),
	.V2C_2 (V2C_587_156),
	.V2C_3 (V2C_587_285),
	.V (V_587)
);

VNU_3 #(quan_width) VNU588 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_588),
	.C2V_2 (C2V_130_588),
	.C2V_3 (C2V_162_588),
	.L (L_588),
	.V2C_1 (V2C_588_3),
	.V2C_2 (V2C_588_130),
	.V2C_3 (V2C_588_162),
	.V (V_588)
);

VNU_3 #(quan_width) VNU589 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_589),
	.C2V_2 (C2V_136_589),
	.C2V_3 (C2V_168_589),
	.L (L_589),
	.V2C_1 (V2C_589_9),
	.V2C_2 (V2C_589_136),
	.V2C_3 (V2C_589_168),
	.V (V_589)
);

VNU_3 #(quan_width) VNU590 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_590),
	.C2V_2 (C2V_142_590),
	.C2V_3 (C2V_174_590),
	.L (L_590),
	.V2C_1 (V2C_590_15),
	.V2C_2 (V2C_590_142),
	.V2C_3 (V2C_590_174),
	.V (V_590)
);

VNU_3 #(quan_width) VNU591 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_591),
	.C2V_2 (C2V_148_591),
	.C2V_3 (C2V_180_591),
	.L (L_591),
	.V2C_1 (V2C_591_21),
	.V2C_2 (V2C_591_148),
	.V2C_3 (V2C_591_180),
	.V (V_591)
);

VNU_3 #(quan_width) VNU592 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_592),
	.C2V_2 (C2V_154_592),
	.C2V_3 (C2V_186_592),
	.L (L_592),
	.V2C_1 (V2C_592_27),
	.V2C_2 (V2C_592_154),
	.V2C_3 (V2C_592_186),
	.V (V_592)
);

VNU_3 #(quan_width) VNU593 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_593),
	.C2V_2 (C2V_160_593),
	.C2V_3 (C2V_192_593),
	.L (L_593),
	.V2C_1 (V2C_593_33),
	.V2C_2 (V2C_593_160),
	.V2C_3 (V2C_593_192),
	.V (V_593)
);

VNU_3 #(quan_width) VNU594 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_594),
	.C2V_2 (C2V_166_594),
	.C2V_3 (C2V_198_594),
	.L (L_594),
	.V2C_1 (V2C_594_39),
	.V2C_2 (V2C_594_166),
	.V2C_3 (V2C_594_198),
	.V (V_594)
);

VNU_3 #(quan_width) VNU595 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_595),
	.C2V_2 (C2V_172_595),
	.C2V_3 (C2V_204_595),
	.L (L_595),
	.V2C_1 (V2C_595_45),
	.V2C_2 (V2C_595_172),
	.V2C_3 (V2C_595_204),
	.V (V_595)
);

VNU_3 #(quan_width) VNU596 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_596),
	.C2V_2 (C2V_178_596),
	.C2V_3 (C2V_210_596),
	.L (L_596),
	.V2C_1 (V2C_596_51),
	.V2C_2 (V2C_596_178),
	.V2C_3 (V2C_596_210),
	.V (V_596)
);

VNU_3 #(quan_width) VNU597 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_597),
	.C2V_2 (C2V_184_597),
	.C2V_3 (C2V_216_597),
	.L (L_597),
	.V2C_1 (V2C_597_57),
	.V2C_2 (V2C_597_184),
	.V2C_3 (V2C_597_216),
	.V (V_597)
);

VNU_3 #(quan_width) VNU598 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_598),
	.C2V_2 (C2V_190_598),
	.C2V_3 (C2V_222_598),
	.L (L_598),
	.V2C_1 (V2C_598_63),
	.V2C_2 (V2C_598_190),
	.V2C_3 (V2C_598_222),
	.V (V_598)
);

VNU_3 #(quan_width) VNU599 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_599),
	.C2V_2 (C2V_196_599),
	.C2V_3 (C2V_228_599),
	.L (L_599),
	.V2C_1 (V2C_599_69),
	.V2C_2 (V2C_599_196),
	.V2C_3 (V2C_599_228),
	.V (V_599)
);

VNU_3 #(quan_width) VNU600 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_600),
	.C2V_2 (C2V_202_600),
	.C2V_3 (C2V_234_600),
	.L (L_600),
	.V2C_1 (V2C_600_75),
	.V2C_2 (V2C_600_202),
	.V2C_3 (V2C_600_234),
	.V (V_600)
);

VNU_3 #(quan_width) VNU601 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_601),
	.C2V_2 (C2V_208_601),
	.C2V_3 (C2V_240_601),
	.L (L_601),
	.V2C_1 (V2C_601_81),
	.V2C_2 (V2C_601_208),
	.V2C_3 (V2C_601_240),
	.V (V_601)
);

VNU_3 #(quan_width) VNU602 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_602),
	.C2V_2 (C2V_214_602),
	.C2V_3 (C2V_246_602),
	.L (L_602),
	.V2C_1 (V2C_602_87),
	.V2C_2 (V2C_602_214),
	.V2C_3 (V2C_602_246),
	.V (V_602)
);

VNU_3 #(quan_width) VNU603 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_93_603),
	.C2V_2 (C2V_220_603),
	.C2V_3 (C2V_252_603),
	.L (L_603),
	.V2C_1 (V2C_603_93),
	.V2C_2 (V2C_603_220),
	.V2C_3 (V2C_603_252),
	.V (V_603)
);

VNU_3 #(quan_width) VNU604 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_99_604),
	.C2V_2 (C2V_226_604),
	.C2V_3 (C2V_258_604),
	.L (L_604),
	.V2C_1 (V2C_604_99),
	.V2C_2 (V2C_604_226),
	.V2C_3 (V2C_604_258),
	.V (V_604)
);

VNU_3 #(quan_width) VNU605 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_105_605),
	.C2V_2 (C2V_232_605),
	.C2V_3 (C2V_264_605),
	.L (L_605),
	.V2C_1 (V2C_605_105),
	.V2C_2 (V2C_605_232),
	.V2C_3 (V2C_605_264),
	.V (V_605)
);

VNU_3 #(quan_width) VNU606 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_111_606),
	.C2V_2 (C2V_238_606),
	.C2V_3 (C2V_270_606),
	.L (L_606),
	.V2C_1 (V2C_606_111),
	.V2C_2 (V2C_606_238),
	.V2C_3 (V2C_606_270),
	.V (V_606)
);

VNU_3 #(quan_width) VNU607 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_117_607),
	.C2V_2 (C2V_244_607),
	.C2V_3 (C2V_276_607),
	.L (L_607),
	.V2C_1 (V2C_607_117),
	.V2C_2 (V2C_607_244),
	.V2C_3 (V2C_607_276),
	.V (V_607)
);

VNU_3 #(quan_width) VNU608 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_123_608),
	.C2V_2 (C2V_250_608),
	.C2V_3 (C2V_282_608),
	.L (L_608),
	.V2C_1 (V2C_608_123),
	.V2C_2 (V2C_608_250),
	.V2C_3 (V2C_608_282),
	.V (V_608)
);

VNU_3 #(quan_width) VNU609 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_129_609),
	.C2V_2 (C2V_256_609),
	.C2V_3 (C2V_288_609),
	.L (L_609),
	.V2C_1 (V2C_609_129),
	.V2C_2 (V2C_609_256),
	.V2C_3 (V2C_609_288),
	.V (V_609)
);

VNU_3 #(quan_width) VNU610 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_610),
	.C2V_2 (C2V_135_610),
	.C2V_3 (C2V_262_610),
	.L (L_610),
	.V2C_1 (V2C_610_6),
	.V2C_2 (V2C_610_135),
	.V2C_3 (V2C_610_262),
	.V (V_610)
);

VNU_3 #(quan_width) VNU611 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_611),
	.C2V_2 (C2V_141_611),
	.C2V_3 (C2V_268_611),
	.L (L_611),
	.V2C_1 (V2C_611_12),
	.V2C_2 (V2C_611_141),
	.V2C_3 (V2C_611_268),
	.V (V_611)
);

VNU_3 #(quan_width) VNU612 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_612),
	.C2V_2 (C2V_147_612),
	.C2V_3 (C2V_274_612),
	.L (L_612),
	.V2C_1 (V2C_612_18),
	.V2C_2 (V2C_612_147),
	.V2C_3 (V2C_612_274),
	.V (V_612)
);

VNU_3 #(quan_width) VNU613 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_613),
	.C2V_2 (C2V_153_613),
	.C2V_3 (C2V_280_613),
	.L (L_613),
	.V2C_1 (V2C_613_24),
	.V2C_2 (V2C_613_153),
	.V2C_3 (V2C_613_280),
	.V (V_613)
);

VNU_3 #(quan_width) VNU614 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_614),
	.C2V_2 (C2V_159_614),
	.C2V_3 (C2V_286_614),
	.L (L_614),
	.V2C_1 (V2C_614_30),
	.V2C_2 (V2C_614_159),
	.V2C_3 (V2C_614_286),
	.V (V_614)
);

VNU_3 #(quan_width) VNU615 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_615),
	.C2V_2 (C2V_36_615),
	.C2V_3 (C2V_165_615),
	.L (L_615),
	.V2C_1 (V2C_615_4),
	.V2C_2 (V2C_615_36),
	.V2C_3 (V2C_615_165),
	.V (V_615)
);

VNU_3 #(quan_width) VNU616 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_616),
	.C2V_2 (C2V_42_616),
	.C2V_3 (C2V_171_616),
	.L (L_616),
	.V2C_1 (V2C_616_10),
	.V2C_2 (V2C_616_42),
	.V2C_3 (V2C_616_171),
	.V (V_616)
);

VNU_3 #(quan_width) VNU617 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_617),
	.C2V_2 (C2V_48_617),
	.C2V_3 (C2V_177_617),
	.L (L_617),
	.V2C_1 (V2C_617_16),
	.V2C_2 (V2C_617_48),
	.V2C_3 (V2C_617_177),
	.V (V_617)
);

VNU_3 #(quan_width) VNU618 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_618),
	.C2V_2 (C2V_54_618),
	.C2V_3 (C2V_183_618),
	.L (L_618),
	.V2C_1 (V2C_618_22),
	.V2C_2 (V2C_618_54),
	.V2C_3 (V2C_618_183),
	.V (V_618)
);

VNU_3 #(quan_width) VNU619 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_619),
	.C2V_2 (C2V_60_619),
	.C2V_3 (C2V_189_619),
	.L (L_619),
	.V2C_1 (V2C_619_28),
	.V2C_2 (V2C_619_60),
	.V2C_3 (V2C_619_189),
	.V (V_619)
);

VNU_3 #(quan_width) VNU620 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_620),
	.C2V_2 (C2V_66_620),
	.C2V_3 (C2V_195_620),
	.L (L_620),
	.V2C_1 (V2C_620_34),
	.V2C_2 (V2C_620_66),
	.V2C_3 (V2C_620_195),
	.V (V_620)
);

VNU_3 #(quan_width) VNU621 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_621),
	.C2V_2 (C2V_72_621),
	.C2V_3 (C2V_201_621),
	.L (L_621),
	.V2C_1 (V2C_621_40),
	.V2C_2 (V2C_621_72),
	.V2C_3 (V2C_621_201),
	.V (V_621)
);

VNU_3 #(quan_width) VNU622 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_622),
	.C2V_2 (C2V_78_622),
	.C2V_3 (C2V_207_622),
	.L (L_622),
	.V2C_1 (V2C_622_46),
	.V2C_2 (V2C_622_78),
	.V2C_3 (V2C_622_207),
	.V (V_622)
);

VNU_3 #(quan_width) VNU623 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_623),
	.C2V_2 (C2V_84_623),
	.C2V_3 (C2V_213_623),
	.L (L_623),
	.V2C_1 (V2C_623_52),
	.V2C_2 (V2C_623_84),
	.V2C_3 (V2C_623_213),
	.V (V_623)
);

VNU_3 #(quan_width) VNU624 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_624),
	.C2V_2 (C2V_90_624),
	.C2V_3 (C2V_219_624),
	.L (L_624),
	.V2C_1 (V2C_624_58),
	.V2C_2 (V2C_624_90),
	.V2C_3 (V2C_624_219),
	.V (V_624)
);

VNU_3 #(quan_width) VNU625 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_625),
	.C2V_2 (C2V_57_625),
	.C2V_3 (C2V_202_625),
	.L (L_625),
	.V2C_1 (V2C_625_8),
	.V2C_2 (V2C_625_57),
	.V2C_3 (V2C_625_202),
	.V (V_625)
);

VNU_3 #(quan_width) VNU626 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_626),
	.C2V_2 (C2V_63_626),
	.C2V_3 (C2V_208_626),
	.L (L_626),
	.V2C_1 (V2C_626_14),
	.V2C_2 (V2C_626_63),
	.V2C_3 (V2C_626_208),
	.V (V_626)
);

VNU_3 #(quan_width) VNU627 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_627),
	.C2V_2 (C2V_69_627),
	.C2V_3 (C2V_214_627),
	.L (L_627),
	.V2C_1 (V2C_627_20),
	.V2C_2 (V2C_627_69),
	.V2C_3 (V2C_627_214),
	.V (V_627)
);

VNU_3 #(quan_width) VNU628 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_628),
	.C2V_2 (C2V_75_628),
	.C2V_3 (C2V_220_628),
	.L (L_628),
	.V2C_1 (V2C_628_26),
	.V2C_2 (V2C_628_75),
	.V2C_3 (V2C_628_220),
	.V (V_628)
);

VNU_3 #(quan_width) VNU629 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_629),
	.C2V_2 (C2V_81_629),
	.C2V_3 (C2V_226_629),
	.L (L_629),
	.V2C_1 (V2C_629_32),
	.V2C_2 (V2C_629_81),
	.V2C_3 (V2C_629_226),
	.V (V_629)
);

VNU_3 #(quan_width) VNU630 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_630),
	.C2V_2 (C2V_87_630),
	.C2V_3 (C2V_232_630),
	.L (L_630),
	.V2C_1 (V2C_630_38),
	.V2C_2 (V2C_630_87),
	.V2C_3 (V2C_630_232),
	.V (V_630)
);

VNU_3 #(quan_width) VNU631 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_631),
	.C2V_2 (C2V_93_631),
	.C2V_3 (C2V_238_631),
	.L (L_631),
	.V2C_1 (V2C_631_44),
	.V2C_2 (V2C_631_93),
	.V2C_3 (V2C_631_238),
	.V (V_631)
);

VNU_3 #(quan_width) VNU632 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_632),
	.C2V_2 (C2V_99_632),
	.C2V_3 (C2V_244_632),
	.L (L_632),
	.V2C_1 (V2C_632_50),
	.V2C_2 (V2C_632_99),
	.V2C_3 (V2C_632_244),
	.V (V_632)
);

VNU_3 #(quan_width) VNU633 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_633),
	.C2V_2 (C2V_105_633),
	.C2V_3 (C2V_250_633),
	.L (L_633),
	.V2C_1 (V2C_633_56),
	.V2C_2 (V2C_633_105),
	.V2C_3 (V2C_633_250),
	.V (V_633)
);

VNU_3 #(quan_width) VNU634 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_634),
	.C2V_2 (C2V_111_634),
	.C2V_3 (C2V_256_634),
	.L (L_634),
	.V2C_1 (V2C_634_62),
	.V2C_2 (V2C_634_111),
	.V2C_3 (V2C_634_256),
	.V (V_634)
);

VNU_3 #(quan_width) VNU635 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_635),
	.C2V_2 (C2V_117_635),
	.C2V_3 (C2V_262_635),
	.L (L_635),
	.V2C_1 (V2C_635_68),
	.V2C_2 (V2C_635_117),
	.V2C_3 (V2C_635_262),
	.V (V_635)
);

VNU_3 #(quan_width) VNU636 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_636),
	.C2V_2 (C2V_123_636),
	.C2V_3 (C2V_268_636),
	.L (L_636),
	.V2C_1 (V2C_636_74),
	.V2C_2 (V2C_636_123),
	.V2C_3 (V2C_636_268),
	.V (V_636)
);

VNU_3 #(quan_width) VNU637 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_80_637),
	.C2V_2 (C2V_129_637),
	.C2V_3 (C2V_274_637),
	.L (L_637),
	.V2C_1 (V2C_637_80),
	.V2C_2 (V2C_637_129),
	.V2C_3 (V2C_637_274),
	.V (V_637)
);

VNU_3 #(quan_width) VNU638 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_86_638),
	.C2V_2 (C2V_135_638),
	.C2V_3 (C2V_280_638),
	.L (L_638),
	.V2C_1 (V2C_638_86),
	.V2C_2 (V2C_638_135),
	.V2C_3 (V2C_638_280),
	.V (V_638)
);

VNU_3 #(quan_width) VNU639 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_92_639),
	.C2V_2 (C2V_141_639),
	.C2V_3 (C2V_286_639),
	.L (L_639),
	.V2C_1 (V2C_639_92),
	.V2C_2 (V2C_639_141),
	.V2C_3 (V2C_639_286),
	.V (V_639)
);

VNU_3 #(quan_width) VNU640 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_640),
	.C2V_2 (C2V_98_640),
	.C2V_3 (C2V_147_640),
	.L (L_640),
	.V2C_1 (V2C_640_4),
	.V2C_2 (V2C_640_98),
	.V2C_3 (V2C_640_147),
	.V (V_640)
);

VNU_3 #(quan_width) VNU641 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_641),
	.C2V_2 (C2V_104_641),
	.C2V_3 (C2V_153_641),
	.L (L_641),
	.V2C_1 (V2C_641_10),
	.V2C_2 (V2C_641_104),
	.V2C_3 (V2C_641_153),
	.V (V_641)
);

VNU_3 #(quan_width) VNU642 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_642),
	.C2V_2 (C2V_110_642),
	.C2V_3 (C2V_159_642),
	.L (L_642),
	.V2C_1 (V2C_642_16),
	.V2C_2 (V2C_642_110),
	.V2C_3 (V2C_642_159),
	.V (V_642)
);

VNU_3 #(quan_width) VNU643 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_643),
	.C2V_2 (C2V_116_643),
	.C2V_3 (C2V_165_643),
	.L (L_643),
	.V2C_1 (V2C_643_22),
	.V2C_2 (V2C_643_116),
	.V2C_3 (V2C_643_165),
	.V (V_643)
);

VNU_3 #(quan_width) VNU644 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_644),
	.C2V_2 (C2V_122_644),
	.C2V_3 (C2V_171_644),
	.L (L_644),
	.V2C_1 (V2C_644_28),
	.V2C_2 (V2C_644_122),
	.V2C_3 (V2C_644_171),
	.V (V_644)
);

VNU_3 #(quan_width) VNU645 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_645),
	.C2V_2 (C2V_128_645),
	.C2V_3 (C2V_177_645),
	.L (L_645),
	.V2C_1 (V2C_645_34),
	.V2C_2 (V2C_645_128),
	.V2C_3 (V2C_645_177),
	.V (V_645)
);

VNU_3 #(quan_width) VNU646 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_646),
	.C2V_2 (C2V_134_646),
	.C2V_3 (C2V_183_646),
	.L (L_646),
	.V2C_1 (V2C_646_40),
	.V2C_2 (V2C_646_134),
	.V2C_3 (V2C_646_183),
	.V (V_646)
);

VNU_3 #(quan_width) VNU647 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_647),
	.C2V_2 (C2V_140_647),
	.C2V_3 (C2V_189_647),
	.L (L_647),
	.V2C_1 (V2C_647_46),
	.V2C_2 (V2C_647_140),
	.V2C_3 (V2C_647_189),
	.V (V_647)
);

VNU_3 #(quan_width) VNU648 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_648),
	.C2V_2 (C2V_146_648),
	.C2V_3 (C2V_195_648),
	.L (L_648),
	.V2C_1 (V2C_648_52),
	.V2C_2 (V2C_648_146),
	.V2C_3 (V2C_648_195),
	.V (V_648)
);

VNU_3 #(quan_width) VNU649 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_649),
	.C2V_2 (C2V_152_649),
	.C2V_3 (C2V_201_649),
	.L (L_649),
	.V2C_1 (V2C_649_58),
	.V2C_2 (V2C_649_152),
	.V2C_3 (V2C_649_201),
	.V (V_649)
);

VNU_3 #(quan_width) VNU650 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_650),
	.C2V_2 (C2V_158_650),
	.C2V_3 (C2V_207_650),
	.L (L_650),
	.V2C_1 (V2C_650_64),
	.V2C_2 (V2C_650_158),
	.V2C_3 (V2C_650_207),
	.V (V_650)
);

VNU_3 #(quan_width) VNU651 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_651),
	.C2V_2 (C2V_164_651),
	.C2V_3 (C2V_213_651),
	.L (L_651),
	.V2C_1 (V2C_651_70),
	.V2C_2 (V2C_651_164),
	.V2C_3 (V2C_651_213),
	.V (V_651)
);

VNU_3 #(quan_width) VNU652 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_652),
	.C2V_2 (C2V_170_652),
	.C2V_3 (C2V_219_652),
	.L (L_652),
	.V2C_1 (V2C_652_76),
	.V2C_2 (V2C_652_170),
	.V2C_3 (V2C_652_219),
	.V (V_652)
);

VNU_3 #(quan_width) VNU653 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_653),
	.C2V_2 (C2V_176_653),
	.C2V_3 (C2V_225_653),
	.L (L_653),
	.V2C_1 (V2C_653_82),
	.V2C_2 (V2C_653_176),
	.V2C_3 (V2C_653_225),
	.V (V_653)
);

VNU_3 #(quan_width) VNU654 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_654),
	.C2V_2 (C2V_182_654),
	.C2V_3 (C2V_231_654),
	.L (L_654),
	.V2C_1 (V2C_654_88),
	.V2C_2 (V2C_654_182),
	.V2C_3 (V2C_654_231),
	.V (V_654)
);

VNU_3 #(quan_width) VNU655 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_655),
	.C2V_2 (C2V_188_655),
	.C2V_3 (C2V_237_655),
	.L (L_655),
	.V2C_1 (V2C_655_94),
	.V2C_2 (V2C_655_188),
	.V2C_3 (V2C_655_237),
	.V (V_655)
);

VNU_3 #(quan_width) VNU656 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_656),
	.C2V_2 (C2V_194_656),
	.C2V_3 (C2V_243_656),
	.L (L_656),
	.V2C_1 (V2C_656_100),
	.V2C_2 (V2C_656_194),
	.V2C_3 (V2C_656_243),
	.V (V_656)
);

VNU_3 #(quan_width) VNU657 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_657),
	.C2V_2 (C2V_200_657),
	.C2V_3 (C2V_249_657),
	.L (L_657),
	.V2C_1 (V2C_657_106),
	.V2C_2 (V2C_657_200),
	.V2C_3 (V2C_657_249),
	.V (V_657)
);

VNU_3 #(quan_width) VNU658 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_658),
	.C2V_2 (C2V_206_658),
	.C2V_3 (C2V_255_658),
	.L (L_658),
	.V2C_1 (V2C_658_112),
	.V2C_2 (V2C_658_206),
	.V2C_3 (V2C_658_255),
	.V (V_658)
);

VNU_3 #(quan_width) VNU659 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_118_659),
	.C2V_2 (C2V_212_659),
	.C2V_3 (C2V_261_659),
	.L (L_659),
	.V2C_1 (V2C_659_118),
	.V2C_2 (V2C_659_212),
	.V2C_3 (V2C_659_261),
	.V (V_659)
);

VNU_3 #(quan_width) VNU660 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_124_660),
	.C2V_2 (C2V_218_660),
	.C2V_3 (C2V_267_660),
	.L (L_660),
	.V2C_1 (V2C_660_124),
	.V2C_2 (V2C_660_218),
	.V2C_3 (V2C_660_267),
	.V (V_660)
);

VNU_3 #(quan_width) VNU661 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_130_661),
	.C2V_2 (C2V_224_661),
	.C2V_3 (C2V_273_661),
	.L (L_661),
	.V2C_1 (V2C_661_130),
	.V2C_2 (V2C_661_224),
	.V2C_3 (V2C_661_273),
	.V (V_661)
);

VNU_3 #(quan_width) VNU662 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_136_662),
	.C2V_2 (C2V_230_662),
	.C2V_3 (C2V_279_662),
	.L (L_662),
	.V2C_1 (V2C_662_136),
	.V2C_2 (V2C_662_230),
	.V2C_3 (V2C_662_279),
	.V (V_662)
);

VNU_3 #(quan_width) VNU663 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_142_663),
	.C2V_2 (C2V_236_663),
	.C2V_3 (C2V_285_663),
	.L (L_663),
	.V2C_1 (V2C_663_142),
	.V2C_2 (V2C_663_236),
	.V2C_3 (V2C_663_285),
	.V (V_663)
);

VNU_3 #(quan_width) VNU664 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_664),
	.C2V_2 (C2V_148_664),
	.C2V_3 (C2V_242_664),
	.L (L_664),
	.V2C_1 (V2C_664_3),
	.V2C_2 (V2C_664_148),
	.V2C_3 (V2C_664_242),
	.V (V_664)
);

VNU_3 #(quan_width) VNU665 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_665),
	.C2V_2 (C2V_154_665),
	.C2V_3 (C2V_248_665),
	.L (L_665),
	.V2C_1 (V2C_665_9),
	.V2C_2 (V2C_665_154),
	.V2C_3 (V2C_665_248),
	.V (V_665)
);

VNU_3 #(quan_width) VNU666 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_666),
	.C2V_2 (C2V_160_666),
	.C2V_3 (C2V_254_666),
	.L (L_666),
	.V2C_1 (V2C_666_15),
	.V2C_2 (V2C_666_160),
	.V2C_3 (V2C_666_254),
	.V (V_666)
);

VNU_3 #(quan_width) VNU667 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_667),
	.C2V_2 (C2V_166_667),
	.C2V_3 (C2V_260_667),
	.L (L_667),
	.V2C_1 (V2C_667_21),
	.V2C_2 (V2C_667_166),
	.V2C_3 (V2C_667_260),
	.V (V_667)
);

VNU_3 #(quan_width) VNU668 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_668),
	.C2V_2 (C2V_172_668),
	.C2V_3 (C2V_266_668),
	.L (L_668),
	.V2C_1 (V2C_668_27),
	.V2C_2 (V2C_668_172),
	.V2C_3 (V2C_668_266),
	.V (V_668)
);

VNU_3 #(quan_width) VNU669 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_669),
	.C2V_2 (C2V_178_669),
	.C2V_3 (C2V_272_669),
	.L (L_669),
	.V2C_1 (V2C_669_33),
	.V2C_2 (V2C_669_178),
	.V2C_3 (V2C_669_272),
	.V (V_669)
);

VNU_3 #(quan_width) VNU670 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_670),
	.C2V_2 (C2V_184_670),
	.C2V_3 (C2V_278_670),
	.L (L_670),
	.V2C_1 (V2C_670_39),
	.V2C_2 (V2C_670_184),
	.V2C_3 (V2C_670_278),
	.V (V_670)
);

VNU_3 #(quan_width) VNU671 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_671),
	.C2V_2 (C2V_190_671),
	.C2V_3 (C2V_284_671),
	.L (L_671),
	.V2C_1 (V2C_671_45),
	.V2C_2 (V2C_671_190),
	.V2C_3 (V2C_671_284),
	.V (V_671)
);

VNU_3 #(quan_width) VNU672 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_672),
	.C2V_2 (C2V_51_672),
	.C2V_3 (C2V_196_672),
	.L (L_672),
	.V2C_1 (V2C_672_2),
	.V2C_2 (V2C_672_51),
	.V2C_3 (V2C_672_196),
	.V (V_672)
);

VNU_3 #(quan_width) VNU673 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_214_673),
	.C2V_2 (C2V_218_673),
	.C2V_3 (C2V_287_673),
	.L (L_673),
	.V2C_1 (V2C_673_214),
	.V2C_2 (V2C_673_218),
	.V2C_3 (V2C_673_287),
	.V (V_673)
);

VNU_3 #(quan_width) VNU674 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_674),
	.C2V_2 (C2V_220_674),
	.C2V_3 (C2V_224_674),
	.L (L_674),
	.V2C_1 (V2C_674_5),
	.V2C_2 (V2C_674_220),
	.V2C_3 (V2C_674_224),
	.V (V_674)
);

VNU_3 #(quan_width) VNU675 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_675),
	.C2V_2 (C2V_226_675),
	.C2V_3 (C2V_230_675),
	.L (L_675),
	.V2C_1 (V2C_675_11),
	.V2C_2 (V2C_675_226),
	.V2C_3 (V2C_675_230),
	.V (V_675)
);

VNU_3 #(quan_width) VNU676 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_676),
	.C2V_2 (C2V_232_676),
	.C2V_3 (C2V_236_676),
	.L (L_676),
	.V2C_1 (V2C_676_17),
	.V2C_2 (V2C_676_232),
	.V2C_3 (V2C_676_236),
	.V (V_676)
);

VNU_3 #(quan_width) VNU677 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_677),
	.C2V_2 (C2V_238_677),
	.C2V_3 (C2V_242_677),
	.L (L_677),
	.V2C_1 (V2C_677_23),
	.V2C_2 (V2C_677_238),
	.V2C_3 (V2C_677_242),
	.V (V_677)
);

VNU_3 #(quan_width) VNU678 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_678),
	.C2V_2 (C2V_244_678),
	.C2V_3 (C2V_248_678),
	.L (L_678),
	.V2C_1 (V2C_678_29),
	.V2C_2 (V2C_678_244),
	.V2C_3 (V2C_678_248),
	.V (V_678)
);

VNU_3 #(quan_width) VNU679 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_679),
	.C2V_2 (C2V_250_679),
	.C2V_3 (C2V_254_679),
	.L (L_679),
	.V2C_1 (V2C_679_35),
	.V2C_2 (V2C_679_250),
	.V2C_3 (V2C_679_254),
	.V (V_679)
);

VNU_3 #(quan_width) VNU680 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_680),
	.C2V_2 (C2V_256_680),
	.C2V_3 (C2V_260_680),
	.L (L_680),
	.V2C_1 (V2C_680_41),
	.V2C_2 (V2C_680_256),
	.V2C_3 (V2C_680_260),
	.V (V_680)
);

VNU_3 #(quan_width) VNU681 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_681),
	.C2V_2 (C2V_262_681),
	.C2V_3 (C2V_266_681),
	.L (L_681),
	.V2C_1 (V2C_681_47),
	.V2C_2 (V2C_681_262),
	.V2C_3 (V2C_681_266),
	.V (V_681)
);

VNU_3 #(quan_width) VNU682 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_682),
	.C2V_2 (C2V_268_682),
	.C2V_3 (C2V_272_682),
	.L (L_682),
	.V2C_1 (V2C_682_53),
	.V2C_2 (V2C_682_268),
	.V2C_3 (V2C_682_272),
	.V (V_682)
);

VNU_3 #(quan_width) VNU683 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_59_683),
	.C2V_2 (C2V_274_683),
	.C2V_3 (C2V_278_683),
	.L (L_683),
	.V2C_1 (V2C_683_59),
	.V2C_2 (V2C_683_274),
	.V2C_3 (V2C_683_278),
	.V (V_683)
);

VNU_3 #(quan_width) VNU684 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_65_684),
	.C2V_2 (C2V_280_684),
	.C2V_3 (C2V_284_684),
	.L (L_684),
	.V2C_1 (V2C_684_65),
	.V2C_2 (V2C_684_280),
	.V2C_3 (V2C_684_284),
	.V (V_684)
);

VNU_3 #(quan_width) VNU685 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_685),
	.C2V_2 (C2V_71_685),
	.C2V_3 (C2V_286_685),
	.L (L_685),
	.V2C_1 (V2C_685_2),
	.V2C_2 (V2C_685_71),
	.V2C_3 (V2C_685_286),
	.V (V_685)
);

VNU_3 #(quan_width) VNU686 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_686),
	.C2V_2 (C2V_8_686),
	.C2V_3 (C2V_77_686),
	.L (L_686),
	.V2C_1 (V2C_686_4),
	.V2C_2 (V2C_686_8),
	.V2C_3 (V2C_686_77),
	.V (V_686)
);

VNU_3 #(quan_width) VNU687 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_687),
	.C2V_2 (C2V_14_687),
	.C2V_3 (C2V_83_687),
	.L (L_687),
	.V2C_1 (V2C_687_10),
	.V2C_2 (V2C_687_14),
	.V2C_3 (V2C_687_83),
	.V (V_687)
);

VNU_3 #(quan_width) VNU688 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_688),
	.C2V_2 (C2V_20_688),
	.C2V_3 (C2V_89_688),
	.L (L_688),
	.V2C_1 (V2C_688_16),
	.V2C_2 (V2C_688_20),
	.V2C_3 (V2C_688_89),
	.V (V_688)
);

VNU_3 #(quan_width) VNU689 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_689),
	.C2V_2 (C2V_26_689),
	.C2V_3 (C2V_95_689),
	.L (L_689),
	.V2C_1 (V2C_689_22),
	.V2C_2 (V2C_689_26),
	.V2C_3 (V2C_689_95),
	.V (V_689)
);

VNU_3 #(quan_width) VNU690 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_690),
	.C2V_2 (C2V_32_690),
	.C2V_3 (C2V_101_690),
	.L (L_690),
	.V2C_1 (V2C_690_28),
	.V2C_2 (V2C_690_32),
	.V2C_3 (V2C_690_101),
	.V (V_690)
);

VNU_3 #(quan_width) VNU691 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_691),
	.C2V_2 (C2V_38_691),
	.C2V_3 (C2V_107_691),
	.L (L_691),
	.V2C_1 (V2C_691_34),
	.V2C_2 (V2C_691_38),
	.V2C_3 (V2C_691_107),
	.V (V_691)
);

VNU_3 #(quan_width) VNU692 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_692),
	.C2V_2 (C2V_44_692),
	.C2V_3 (C2V_113_692),
	.L (L_692),
	.V2C_1 (V2C_692_40),
	.V2C_2 (V2C_692_44),
	.V2C_3 (V2C_692_113),
	.V (V_692)
);

VNU_3 #(quan_width) VNU693 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_693),
	.C2V_2 (C2V_50_693),
	.C2V_3 (C2V_119_693),
	.L (L_693),
	.V2C_1 (V2C_693_46),
	.V2C_2 (V2C_693_50),
	.V2C_3 (V2C_693_119),
	.V (V_693)
);

VNU_3 #(quan_width) VNU694 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_694),
	.C2V_2 (C2V_56_694),
	.C2V_3 (C2V_125_694),
	.L (L_694),
	.V2C_1 (V2C_694_52),
	.V2C_2 (V2C_694_56),
	.V2C_3 (V2C_694_125),
	.V (V_694)
);

VNU_3 #(quan_width) VNU695 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_695),
	.C2V_2 (C2V_62_695),
	.C2V_3 (C2V_131_695),
	.L (L_695),
	.V2C_1 (V2C_695_58),
	.V2C_2 (V2C_695_62),
	.V2C_3 (V2C_695_131),
	.V (V_695)
);

VNU_3 #(quan_width) VNU696 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_696),
	.C2V_2 (C2V_68_696),
	.C2V_3 (C2V_137_696),
	.L (L_696),
	.V2C_1 (V2C_696_64),
	.V2C_2 (V2C_696_68),
	.V2C_3 (V2C_696_137),
	.V (V_696)
);

VNU_3 #(quan_width) VNU697 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_697),
	.C2V_2 (C2V_74_697),
	.C2V_3 (C2V_143_697),
	.L (L_697),
	.V2C_1 (V2C_697_70),
	.V2C_2 (V2C_697_74),
	.V2C_3 (V2C_697_143),
	.V (V_697)
);

VNU_3 #(quan_width) VNU698 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_698),
	.C2V_2 (C2V_80_698),
	.C2V_3 (C2V_149_698),
	.L (L_698),
	.V2C_1 (V2C_698_76),
	.V2C_2 (V2C_698_80),
	.V2C_3 (V2C_698_149),
	.V (V_698)
);

VNU_3 #(quan_width) VNU699 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_699),
	.C2V_2 (C2V_86_699),
	.C2V_3 (C2V_155_699),
	.L (L_699),
	.V2C_1 (V2C_699_82),
	.V2C_2 (V2C_699_86),
	.V2C_3 (V2C_699_155),
	.V (V_699)
);

VNU_3 #(quan_width) VNU700 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_700),
	.C2V_2 (C2V_92_700),
	.C2V_3 (C2V_161_700),
	.L (L_700),
	.V2C_1 (V2C_700_88),
	.V2C_2 (V2C_700_92),
	.V2C_3 (V2C_700_161),
	.V (V_700)
);

VNU_3 #(quan_width) VNU701 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_701),
	.C2V_2 (C2V_98_701),
	.C2V_3 (C2V_167_701),
	.L (L_701),
	.V2C_1 (V2C_701_94),
	.V2C_2 (V2C_701_98),
	.V2C_3 (V2C_701_167),
	.V (V_701)
);

VNU_3 #(quan_width) VNU702 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_702),
	.C2V_2 (C2V_104_702),
	.C2V_3 (C2V_173_702),
	.L (L_702),
	.V2C_1 (V2C_702_100),
	.V2C_2 (V2C_702_104),
	.V2C_3 (V2C_702_173),
	.V (V_702)
);

VNU_3 #(quan_width) VNU703 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_703),
	.C2V_2 (C2V_110_703),
	.C2V_3 (C2V_179_703),
	.L (L_703),
	.V2C_1 (V2C_703_106),
	.V2C_2 (V2C_703_110),
	.V2C_3 (V2C_703_179),
	.V (V_703)
);

VNU_3 #(quan_width) VNU704 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_704),
	.C2V_2 (C2V_116_704),
	.C2V_3 (C2V_185_704),
	.L (L_704),
	.V2C_1 (V2C_704_112),
	.V2C_2 (V2C_704_116),
	.V2C_3 (V2C_704_185),
	.V (V_704)
);

VNU_3 #(quan_width) VNU705 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_118_705),
	.C2V_2 (C2V_122_705),
	.C2V_3 (C2V_191_705),
	.L (L_705),
	.V2C_1 (V2C_705_118),
	.V2C_2 (V2C_705_122),
	.V2C_3 (V2C_705_191),
	.V (V_705)
);

VNU_3 #(quan_width) VNU706 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_124_706),
	.C2V_2 (C2V_128_706),
	.C2V_3 (C2V_197_706),
	.L (L_706),
	.V2C_1 (V2C_706_124),
	.V2C_2 (V2C_706_128),
	.V2C_3 (V2C_706_197),
	.V (V_706)
);

VNU_3 #(quan_width) VNU707 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_130_707),
	.C2V_2 (C2V_134_707),
	.C2V_3 (C2V_203_707),
	.L (L_707),
	.V2C_1 (V2C_707_130),
	.V2C_2 (V2C_707_134),
	.V2C_3 (V2C_707_203),
	.V (V_707)
);

VNU_3 #(quan_width) VNU708 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_136_708),
	.C2V_2 (C2V_140_708),
	.C2V_3 (C2V_209_708),
	.L (L_708),
	.V2C_1 (V2C_708_136),
	.V2C_2 (V2C_708_140),
	.V2C_3 (V2C_708_209),
	.V (V_708)
);

VNU_3 #(quan_width) VNU709 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_142_709),
	.C2V_2 (C2V_146_709),
	.C2V_3 (C2V_215_709),
	.L (L_709),
	.V2C_1 (V2C_709_142),
	.V2C_2 (V2C_709_146),
	.V2C_3 (V2C_709_215),
	.V (V_709)
);

VNU_3 #(quan_width) VNU710 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_148_710),
	.C2V_2 (C2V_152_710),
	.C2V_3 (C2V_221_710),
	.L (L_710),
	.V2C_1 (V2C_710_148),
	.V2C_2 (V2C_710_152),
	.V2C_3 (V2C_710_221),
	.V (V_710)
);

VNU_3 #(quan_width) VNU711 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_154_711),
	.C2V_2 (C2V_158_711),
	.C2V_3 (C2V_227_711),
	.L (L_711),
	.V2C_1 (V2C_711_154),
	.V2C_2 (V2C_711_158),
	.V2C_3 (V2C_711_227),
	.V (V_711)
);

VNU_3 #(quan_width) VNU712 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_160_712),
	.C2V_2 (C2V_164_712),
	.C2V_3 (C2V_233_712),
	.L (L_712),
	.V2C_1 (V2C_712_160),
	.V2C_2 (V2C_712_164),
	.V2C_3 (V2C_712_233),
	.V (V_712)
);

VNU_3 #(quan_width) VNU713 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_166_713),
	.C2V_2 (C2V_170_713),
	.C2V_3 (C2V_239_713),
	.L (L_713),
	.V2C_1 (V2C_713_166),
	.V2C_2 (V2C_713_170),
	.V2C_3 (V2C_713_239),
	.V (V_713)
);

VNU_3 #(quan_width) VNU714 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_172_714),
	.C2V_2 (C2V_176_714),
	.C2V_3 (C2V_245_714),
	.L (L_714),
	.V2C_1 (V2C_714_172),
	.V2C_2 (V2C_714_176),
	.V2C_3 (V2C_714_245),
	.V (V_714)
);

VNU_3 #(quan_width) VNU715 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_178_715),
	.C2V_2 (C2V_182_715),
	.C2V_3 (C2V_251_715),
	.L (L_715),
	.V2C_1 (V2C_715_178),
	.V2C_2 (V2C_715_182),
	.V2C_3 (V2C_715_251),
	.V (V_715)
);

VNU_3 #(quan_width) VNU716 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_184_716),
	.C2V_2 (C2V_188_716),
	.C2V_3 (C2V_257_716),
	.L (L_716),
	.V2C_1 (V2C_716_184),
	.V2C_2 (V2C_716_188),
	.V2C_3 (V2C_716_257),
	.V (V_716)
);

VNU_3 #(quan_width) VNU717 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_190_717),
	.C2V_2 (C2V_194_717),
	.C2V_3 (C2V_263_717),
	.L (L_717),
	.V2C_1 (V2C_717_190),
	.V2C_2 (V2C_717_194),
	.V2C_3 (V2C_717_263),
	.V (V_717)
);

VNU_3 #(quan_width) VNU718 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_196_718),
	.C2V_2 (C2V_200_718),
	.C2V_3 (C2V_269_718),
	.L (L_718),
	.V2C_1 (V2C_718_196),
	.V2C_2 (V2C_718_200),
	.V2C_3 (V2C_718_269),
	.V (V_718)
);

VNU_3 #(quan_width) VNU719 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_202_719),
	.C2V_2 (C2V_206_719),
	.C2V_3 (C2V_275_719),
	.L (L_719),
	.V2C_1 (V2C_719_202),
	.V2C_2 (V2C_719_206),
	.V2C_3 (V2C_719_275),
	.V (V_719)
);

VNU_3 #(quan_width) VNU720 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_208_720),
	.C2V_2 (C2V_212_720),
	.C2V_3 (C2V_281_720),
	.L (L_720),
	.V2C_1 (V2C_720_208),
	.V2C_2 (V2C_720_212),
	.V2C_3 (V2C_720_281),
	.V (V_720)
);

VNU_3 #(quan_width) VNU721 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_721),
	.C2V_2 (C2V_43_721),
	.C2V_3 (C2V_191_721),
	.L (L_721),
	.V2C_1 (V2C_721_9),
	.V2C_2 (V2C_721_43),
	.V2C_3 (V2C_721_191),
	.V (V_721)
);

VNU_3 #(quan_width) VNU722 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_722),
	.C2V_2 (C2V_49_722),
	.C2V_3 (C2V_197_722),
	.L (L_722),
	.V2C_1 (V2C_722_15),
	.V2C_2 (V2C_722_49),
	.V2C_3 (V2C_722_197),
	.V (V_722)
);

VNU_3 #(quan_width) VNU723 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_723),
	.C2V_2 (C2V_55_723),
	.C2V_3 (C2V_203_723),
	.L (L_723),
	.V2C_1 (V2C_723_21),
	.V2C_2 (V2C_723_55),
	.V2C_3 (V2C_723_203),
	.V (V_723)
);

VNU_3 #(quan_width) VNU724 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_724),
	.C2V_2 (C2V_61_724),
	.C2V_3 (C2V_209_724),
	.L (L_724),
	.V2C_1 (V2C_724_27),
	.V2C_2 (V2C_724_61),
	.V2C_3 (V2C_724_209),
	.V (V_724)
);

VNU_3 #(quan_width) VNU725 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_725),
	.C2V_2 (C2V_67_725),
	.C2V_3 (C2V_215_725),
	.L (L_725),
	.V2C_1 (V2C_725_33),
	.V2C_2 (V2C_725_67),
	.V2C_3 (V2C_725_215),
	.V (V_725)
);

VNU_3 #(quan_width) VNU726 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_726),
	.C2V_2 (C2V_73_726),
	.C2V_3 (C2V_221_726),
	.L (L_726),
	.V2C_1 (V2C_726_39),
	.V2C_2 (V2C_726_73),
	.V2C_3 (V2C_726_221),
	.V (V_726)
);

VNU_3 #(quan_width) VNU727 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_727),
	.C2V_2 (C2V_79_727),
	.C2V_3 (C2V_227_727),
	.L (L_727),
	.V2C_1 (V2C_727_45),
	.V2C_2 (V2C_727_79),
	.V2C_3 (V2C_727_227),
	.V (V_727)
);

VNU_3 #(quan_width) VNU728 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_728),
	.C2V_2 (C2V_85_728),
	.C2V_3 (C2V_233_728),
	.L (L_728),
	.V2C_1 (V2C_728_51),
	.V2C_2 (V2C_728_85),
	.V2C_3 (V2C_728_233),
	.V (V_728)
);

VNU_3 #(quan_width) VNU729 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_729),
	.C2V_2 (C2V_91_729),
	.C2V_3 (C2V_239_729),
	.L (L_729),
	.V2C_1 (V2C_729_57),
	.V2C_2 (V2C_729_91),
	.V2C_3 (V2C_729_239),
	.V (V_729)
);

VNU_3 #(quan_width) VNU730 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_730),
	.C2V_2 (C2V_97_730),
	.C2V_3 (C2V_245_730),
	.L (L_730),
	.V2C_1 (V2C_730_63),
	.V2C_2 (V2C_730_97),
	.V2C_3 (V2C_730_245),
	.V (V_730)
);

VNU_3 #(quan_width) VNU731 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_731),
	.C2V_2 (C2V_103_731),
	.C2V_3 (C2V_251_731),
	.L (L_731),
	.V2C_1 (V2C_731_69),
	.V2C_2 (V2C_731_103),
	.V2C_3 (V2C_731_251),
	.V (V_731)
);

VNU_3 #(quan_width) VNU732 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_732),
	.C2V_2 (C2V_109_732),
	.C2V_3 (C2V_257_732),
	.L (L_732),
	.V2C_1 (V2C_732_75),
	.V2C_2 (V2C_732_109),
	.V2C_3 (V2C_732_257),
	.V (V_732)
);

VNU_3 #(quan_width) VNU733 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_733),
	.C2V_2 (C2V_115_733),
	.C2V_3 (C2V_263_733),
	.L (L_733),
	.V2C_1 (V2C_733_81),
	.V2C_2 (V2C_733_115),
	.V2C_3 (V2C_733_263),
	.V (V_733)
);

VNU_3 #(quan_width) VNU734 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_734),
	.C2V_2 (C2V_121_734),
	.C2V_3 (C2V_269_734),
	.L (L_734),
	.V2C_1 (V2C_734_87),
	.V2C_2 (V2C_734_121),
	.V2C_3 (V2C_734_269),
	.V (V_734)
);

VNU_3 #(quan_width) VNU735 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_93_735),
	.C2V_2 (C2V_127_735),
	.C2V_3 (C2V_275_735),
	.L (L_735),
	.V2C_1 (V2C_735_93),
	.V2C_2 (V2C_735_127),
	.V2C_3 (V2C_735_275),
	.V (V_735)
);

VNU_3 #(quan_width) VNU736 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_99_736),
	.C2V_2 (C2V_133_736),
	.C2V_3 (C2V_281_736),
	.L (L_736),
	.V2C_1 (V2C_736_99),
	.V2C_2 (V2C_736_133),
	.V2C_3 (V2C_736_281),
	.V (V_736)
);

VNU_3 #(quan_width) VNU737 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_105_737),
	.C2V_2 (C2V_139_737),
	.C2V_3 (C2V_287_737),
	.L (L_737),
	.V2C_1 (V2C_737_105),
	.V2C_2 (V2C_737_139),
	.V2C_3 (V2C_737_287),
	.V (V_737)
);

VNU_3 #(quan_width) VNU738 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_738),
	.C2V_2 (C2V_111_738),
	.C2V_3 (C2V_145_738),
	.L (L_738),
	.V2C_1 (V2C_738_5),
	.V2C_2 (V2C_738_111),
	.V2C_3 (V2C_738_145),
	.V (V_738)
);

VNU_3 #(quan_width) VNU739 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_739),
	.C2V_2 (C2V_117_739),
	.C2V_3 (C2V_151_739),
	.L (L_739),
	.V2C_1 (V2C_739_11),
	.V2C_2 (V2C_739_117),
	.V2C_3 (V2C_739_151),
	.V (V_739)
);

VNU_3 #(quan_width) VNU740 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_740),
	.C2V_2 (C2V_123_740),
	.C2V_3 (C2V_157_740),
	.L (L_740),
	.V2C_1 (V2C_740_17),
	.V2C_2 (V2C_740_123),
	.V2C_3 (V2C_740_157),
	.V (V_740)
);

VNU_3 #(quan_width) VNU741 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_741),
	.C2V_2 (C2V_129_741),
	.C2V_3 (C2V_163_741),
	.L (L_741),
	.V2C_1 (V2C_741_23),
	.V2C_2 (V2C_741_129),
	.V2C_3 (V2C_741_163),
	.V (V_741)
);

VNU_3 #(quan_width) VNU742 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_742),
	.C2V_2 (C2V_135_742),
	.C2V_3 (C2V_169_742),
	.L (L_742),
	.V2C_1 (V2C_742_29),
	.V2C_2 (V2C_742_135),
	.V2C_3 (V2C_742_169),
	.V (V_742)
);

VNU_3 #(quan_width) VNU743 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_743),
	.C2V_2 (C2V_141_743),
	.C2V_3 (C2V_175_743),
	.L (L_743),
	.V2C_1 (V2C_743_35),
	.V2C_2 (V2C_743_141),
	.V2C_3 (V2C_743_175),
	.V (V_743)
);

VNU_3 #(quan_width) VNU744 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_744),
	.C2V_2 (C2V_147_744),
	.C2V_3 (C2V_181_744),
	.L (L_744),
	.V2C_1 (V2C_744_41),
	.V2C_2 (V2C_744_147),
	.V2C_3 (V2C_744_181),
	.V (V_744)
);

VNU_3 #(quan_width) VNU745 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_745),
	.C2V_2 (C2V_153_745),
	.C2V_3 (C2V_187_745),
	.L (L_745),
	.V2C_1 (V2C_745_47),
	.V2C_2 (V2C_745_153),
	.V2C_3 (V2C_745_187),
	.V (V_745)
);

VNU_3 #(quan_width) VNU746 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_746),
	.C2V_2 (C2V_159_746),
	.C2V_3 (C2V_193_746),
	.L (L_746),
	.V2C_1 (V2C_746_53),
	.V2C_2 (V2C_746_159),
	.V2C_3 (V2C_746_193),
	.V (V_746)
);

VNU_3 #(quan_width) VNU747 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_59_747),
	.C2V_2 (C2V_165_747),
	.C2V_3 (C2V_199_747),
	.L (L_747),
	.V2C_1 (V2C_747_59),
	.V2C_2 (V2C_747_165),
	.V2C_3 (V2C_747_199),
	.V (V_747)
);

VNU_3 #(quan_width) VNU748 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_65_748),
	.C2V_2 (C2V_171_748),
	.C2V_3 (C2V_205_748),
	.L (L_748),
	.V2C_1 (V2C_748_65),
	.V2C_2 (V2C_748_171),
	.V2C_3 (V2C_748_205),
	.V (V_748)
);

VNU_3 #(quan_width) VNU749 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_71_749),
	.C2V_2 (C2V_177_749),
	.C2V_3 (C2V_211_749),
	.L (L_749),
	.V2C_1 (V2C_749_71),
	.V2C_2 (V2C_749_177),
	.V2C_3 (V2C_749_211),
	.V (V_749)
);

VNU_3 #(quan_width) VNU750 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_77_750),
	.C2V_2 (C2V_183_750),
	.C2V_3 (C2V_217_750),
	.L (L_750),
	.V2C_1 (V2C_750_77),
	.V2C_2 (V2C_750_183),
	.V2C_3 (V2C_750_217),
	.V (V_750)
);

VNU_3 #(quan_width) VNU751 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_83_751),
	.C2V_2 (C2V_189_751),
	.C2V_3 (C2V_223_751),
	.L (L_751),
	.V2C_1 (V2C_751_83),
	.V2C_2 (V2C_751_189),
	.V2C_3 (V2C_751_223),
	.V (V_751)
);

VNU_3 #(quan_width) VNU752 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_89_752),
	.C2V_2 (C2V_195_752),
	.C2V_3 (C2V_229_752),
	.L (L_752),
	.V2C_1 (V2C_752_89),
	.V2C_2 (V2C_752_195),
	.V2C_3 (V2C_752_229),
	.V (V_752)
);

VNU_3 #(quan_width) VNU753 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_95_753),
	.C2V_2 (C2V_201_753),
	.C2V_3 (C2V_235_753),
	.L (L_753),
	.V2C_1 (V2C_753_95),
	.V2C_2 (V2C_753_201),
	.V2C_3 (V2C_753_235),
	.V (V_753)
);

VNU_3 #(quan_width) VNU754 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_101_754),
	.C2V_2 (C2V_207_754),
	.C2V_3 (C2V_241_754),
	.L (L_754),
	.V2C_1 (V2C_754_101),
	.V2C_2 (V2C_754_207),
	.V2C_3 (V2C_754_241),
	.V (V_754)
);

VNU_3 #(quan_width) VNU755 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_107_755),
	.C2V_2 (C2V_213_755),
	.C2V_3 (C2V_247_755),
	.L (L_755),
	.V2C_1 (V2C_755_107),
	.V2C_2 (V2C_755_213),
	.V2C_3 (V2C_755_247),
	.V (V_755)
);

VNU_3 #(quan_width) VNU756 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_113_756),
	.C2V_2 (C2V_219_756),
	.C2V_3 (C2V_253_756),
	.L (L_756),
	.V2C_1 (V2C_756_113),
	.V2C_2 (V2C_756_219),
	.V2C_3 (V2C_756_253),
	.V (V_756)
);

VNU_3 #(quan_width) VNU757 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_119_757),
	.C2V_2 (C2V_225_757),
	.C2V_3 (C2V_259_757),
	.L (L_757),
	.V2C_1 (V2C_757_119),
	.V2C_2 (V2C_757_225),
	.V2C_3 (V2C_757_259),
	.V (V_757)
);

VNU_3 #(quan_width) VNU758 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_125_758),
	.C2V_2 (C2V_231_758),
	.C2V_3 (C2V_265_758),
	.L (L_758),
	.V2C_1 (V2C_758_125),
	.V2C_2 (V2C_758_231),
	.V2C_3 (V2C_758_265),
	.V (V_758)
);

VNU_3 #(quan_width) VNU759 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_131_759),
	.C2V_2 (C2V_237_759),
	.C2V_3 (C2V_271_759),
	.L (L_759),
	.V2C_1 (V2C_759_131),
	.V2C_2 (V2C_759_237),
	.V2C_3 (V2C_759_271),
	.V (V_759)
);

VNU_3 #(quan_width) VNU760 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_137_760),
	.C2V_2 (C2V_243_760),
	.C2V_3 (C2V_277_760),
	.L (L_760),
	.V2C_1 (V2C_760_137),
	.V2C_2 (V2C_760_243),
	.V2C_3 (V2C_760_277),
	.V (V_760)
);

VNU_3 #(quan_width) VNU761 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_143_761),
	.C2V_2 (C2V_249_761),
	.C2V_3 (C2V_283_761),
	.L (L_761),
	.V2C_1 (V2C_761_143),
	.V2C_2 (V2C_761_249),
	.V2C_3 (V2C_761_283),
	.V (V_761)
);

VNU_3 #(quan_width) VNU762 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_762),
	.C2V_2 (C2V_149_762),
	.C2V_3 (C2V_255_762),
	.L (L_762),
	.V2C_1 (V2C_762_1),
	.V2C_2 (V2C_762_149),
	.V2C_3 (V2C_762_255),
	.V (V_762)
);

VNU_3 #(quan_width) VNU763 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_763),
	.C2V_2 (C2V_155_763),
	.C2V_3 (C2V_261_763),
	.L (L_763),
	.V2C_1 (V2C_763_7),
	.V2C_2 (V2C_763_155),
	.V2C_3 (V2C_763_261),
	.V (V_763)
);

VNU_3 #(quan_width) VNU764 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_764),
	.C2V_2 (C2V_161_764),
	.C2V_3 (C2V_267_764),
	.L (L_764),
	.V2C_1 (V2C_764_13),
	.V2C_2 (V2C_764_161),
	.V2C_3 (V2C_764_267),
	.V (V_764)
);

VNU_3 #(quan_width) VNU765 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_765),
	.C2V_2 (C2V_167_765),
	.C2V_3 (C2V_273_765),
	.L (L_765),
	.V2C_1 (V2C_765_19),
	.V2C_2 (V2C_765_167),
	.V2C_3 (V2C_765_273),
	.V (V_765)
);

VNU_3 #(quan_width) VNU766 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_766),
	.C2V_2 (C2V_173_766),
	.C2V_3 (C2V_279_766),
	.L (L_766),
	.V2C_1 (V2C_766_25),
	.V2C_2 (V2C_766_173),
	.V2C_3 (V2C_766_279),
	.V (V_766)
);

VNU_3 #(quan_width) VNU767 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_767),
	.C2V_2 (C2V_179_767),
	.C2V_3 (C2V_285_767),
	.L (L_767),
	.V2C_1 (V2C_767_31),
	.V2C_2 (V2C_767_179),
	.V2C_3 (V2C_767_285),
	.V (V_767)
);

VNU_3 #(quan_width) VNU768 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_768),
	.C2V_2 (C2V_37_768),
	.C2V_3 (C2V_185_768),
	.L (L_768),
	.V2C_1 (V2C_768_3),
	.V2C_2 (V2C_768_37),
	.V2C_3 (V2C_768_185),
	.V (V_768)
);

VNU_3 #(quan_width) VNU769 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_769),
	.C2V_2 (C2V_43_769),
	.C2V_3 (C2V_155_769),
	.L (L_769),
	.V2C_1 (V2C_769_24),
	.V2C_2 (V2C_769_43),
	.V2C_3 (V2C_769_155),
	.V (V_769)
);

VNU_3 #(quan_width) VNU770 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_770),
	.C2V_2 (C2V_49_770),
	.C2V_3 (C2V_161_770),
	.L (L_770),
	.V2C_1 (V2C_770_30),
	.V2C_2 (V2C_770_49),
	.V2C_3 (V2C_770_161),
	.V (V_770)
);

VNU_3 #(quan_width) VNU771 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_771),
	.C2V_2 (C2V_55_771),
	.C2V_3 (C2V_167_771),
	.L (L_771),
	.V2C_1 (V2C_771_36),
	.V2C_2 (V2C_771_55),
	.V2C_3 (V2C_771_167),
	.V (V_771)
);

VNU_3 #(quan_width) VNU772 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_772),
	.C2V_2 (C2V_61_772),
	.C2V_3 (C2V_173_772),
	.L (L_772),
	.V2C_1 (V2C_772_42),
	.V2C_2 (V2C_772_61),
	.V2C_3 (V2C_772_173),
	.V (V_772)
);

VNU_3 #(quan_width) VNU773 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_773),
	.C2V_2 (C2V_67_773),
	.C2V_3 (C2V_179_773),
	.L (L_773),
	.V2C_1 (V2C_773_48),
	.V2C_2 (V2C_773_67),
	.V2C_3 (V2C_773_179),
	.V (V_773)
);

VNU_3 #(quan_width) VNU774 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_54_774),
	.C2V_2 (C2V_73_774),
	.C2V_3 (C2V_185_774),
	.L (L_774),
	.V2C_1 (V2C_774_54),
	.V2C_2 (V2C_774_73),
	.V2C_3 (V2C_774_185),
	.V (V_774)
);

VNU_3 #(quan_width) VNU775 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_60_775),
	.C2V_2 (C2V_79_775),
	.C2V_3 (C2V_191_775),
	.L (L_775),
	.V2C_1 (V2C_775_60),
	.V2C_2 (V2C_775_79),
	.V2C_3 (V2C_775_191),
	.V (V_775)
);

VNU_3 #(quan_width) VNU776 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_66_776),
	.C2V_2 (C2V_85_776),
	.C2V_3 (C2V_197_776),
	.L (L_776),
	.V2C_1 (V2C_776_66),
	.V2C_2 (V2C_776_85),
	.V2C_3 (V2C_776_197),
	.V (V_776)
);

VNU_3 #(quan_width) VNU777 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_72_777),
	.C2V_2 (C2V_91_777),
	.C2V_3 (C2V_203_777),
	.L (L_777),
	.V2C_1 (V2C_777_72),
	.V2C_2 (V2C_777_91),
	.V2C_3 (V2C_777_203),
	.V (V_777)
);

VNU_3 #(quan_width) VNU778 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_78_778),
	.C2V_2 (C2V_97_778),
	.C2V_3 (C2V_209_778),
	.L (L_778),
	.V2C_1 (V2C_778_78),
	.V2C_2 (V2C_778_97),
	.V2C_3 (V2C_778_209),
	.V (V_778)
);

VNU_3 #(quan_width) VNU779 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_84_779),
	.C2V_2 (C2V_103_779),
	.C2V_3 (C2V_215_779),
	.L (L_779),
	.V2C_1 (V2C_779_84),
	.V2C_2 (V2C_779_103),
	.V2C_3 (V2C_779_215),
	.V (V_779)
);

VNU_3 #(quan_width) VNU780 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_90_780),
	.C2V_2 (C2V_109_780),
	.C2V_3 (C2V_221_780),
	.L (L_780),
	.V2C_1 (V2C_780_90),
	.V2C_2 (V2C_780_109),
	.V2C_3 (V2C_780_221),
	.V (V_780)
);

VNU_3 #(quan_width) VNU781 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_96_781),
	.C2V_2 (C2V_115_781),
	.C2V_3 (C2V_227_781),
	.L (L_781),
	.V2C_1 (V2C_781_96),
	.V2C_2 (V2C_781_115),
	.V2C_3 (V2C_781_227),
	.V (V_781)
);

VNU_3 #(quan_width) VNU782 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_102_782),
	.C2V_2 (C2V_121_782),
	.C2V_3 (C2V_233_782),
	.L (L_782),
	.V2C_1 (V2C_782_102),
	.V2C_2 (V2C_782_121),
	.V2C_3 (V2C_782_233),
	.V (V_782)
);

VNU_3 #(quan_width) VNU783 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_108_783),
	.C2V_2 (C2V_127_783),
	.C2V_3 (C2V_239_783),
	.L (L_783),
	.V2C_1 (V2C_783_108),
	.V2C_2 (V2C_783_127),
	.V2C_3 (V2C_783_239),
	.V (V_783)
);

VNU_3 #(quan_width) VNU784 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_114_784),
	.C2V_2 (C2V_133_784),
	.C2V_3 (C2V_245_784),
	.L (L_784),
	.V2C_1 (V2C_784_114),
	.V2C_2 (V2C_784_133),
	.V2C_3 (V2C_784_245),
	.V (V_784)
);

VNU_3 #(quan_width) VNU785 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_120_785),
	.C2V_2 (C2V_139_785),
	.C2V_3 (C2V_251_785),
	.L (L_785),
	.V2C_1 (V2C_785_120),
	.V2C_2 (V2C_785_139),
	.V2C_3 (V2C_785_251),
	.V (V_785)
);

VNU_3 #(quan_width) VNU786 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_126_786),
	.C2V_2 (C2V_145_786),
	.C2V_3 (C2V_257_786),
	.L (L_786),
	.V2C_1 (V2C_786_126),
	.V2C_2 (V2C_786_145),
	.V2C_3 (V2C_786_257),
	.V (V_786)
);

VNU_3 #(quan_width) VNU787 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_132_787),
	.C2V_2 (C2V_151_787),
	.C2V_3 (C2V_263_787),
	.L (L_787),
	.V2C_1 (V2C_787_132),
	.V2C_2 (V2C_787_151),
	.V2C_3 (V2C_787_263),
	.V (V_787)
);

VNU_3 #(quan_width) VNU788 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_138_788),
	.C2V_2 (C2V_157_788),
	.C2V_3 (C2V_269_788),
	.L (L_788),
	.V2C_1 (V2C_788_138),
	.V2C_2 (V2C_788_157),
	.V2C_3 (V2C_788_269),
	.V (V_788)
);

VNU_3 #(quan_width) VNU789 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_144_789),
	.C2V_2 (C2V_163_789),
	.C2V_3 (C2V_275_789),
	.L (L_789),
	.V2C_1 (V2C_789_144),
	.V2C_2 (V2C_789_163),
	.V2C_3 (V2C_789_275),
	.V (V_789)
);

VNU_3 #(quan_width) VNU790 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_150_790),
	.C2V_2 (C2V_169_790),
	.C2V_3 (C2V_281_790),
	.L (L_790),
	.V2C_1 (V2C_790_150),
	.V2C_2 (V2C_790_169),
	.V2C_3 (V2C_790_281),
	.V (V_790)
);

VNU_3 #(quan_width) VNU791 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_156_791),
	.C2V_2 (C2V_175_791),
	.C2V_3 (C2V_287_791),
	.L (L_791),
	.V2C_1 (V2C_791_156),
	.V2C_2 (V2C_791_175),
	.V2C_3 (V2C_791_287),
	.V (V_791)
);

VNU_3 #(quan_width) VNU792 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_792),
	.C2V_2 (C2V_162_792),
	.C2V_3 (C2V_181_792),
	.L (L_792),
	.V2C_1 (V2C_792_5),
	.V2C_2 (V2C_792_162),
	.V2C_3 (V2C_792_181),
	.V (V_792)
);

VNU_3 #(quan_width) VNU793 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_793),
	.C2V_2 (C2V_168_793),
	.C2V_3 (C2V_187_793),
	.L (L_793),
	.V2C_1 (V2C_793_11),
	.V2C_2 (V2C_793_168),
	.V2C_3 (V2C_793_187),
	.V (V_793)
);

VNU_3 #(quan_width) VNU794 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_794),
	.C2V_2 (C2V_174_794),
	.C2V_3 (C2V_193_794),
	.L (L_794),
	.V2C_1 (V2C_794_17),
	.V2C_2 (V2C_794_174),
	.V2C_3 (V2C_794_193),
	.V (V_794)
);

VNU_3 #(quan_width) VNU795 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_795),
	.C2V_2 (C2V_180_795),
	.C2V_3 (C2V_199_795),
	.L (L_795),
	.V2C_1 (V2C_795_23),
	.V2C_2 (V2C_795_180),
	.V2C_3 (V2C_795_199),
	.V (V_795)
);

VNU_3 #(quan_width) VNU796 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_796),
	.C2V_2 (C2V_186_796),
	.C2V_3 (C2V_205_796),
	.L (L_796),
	.V2C_1 (V2C_796_29),
	.V2C_2 (V2C_796_186),
	.V2C_3 (V2C_796_205),
	.V (V_796)
);

VNU_3 #(quan_width) VNU797 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_797),
	.C2V_2 (C2V_192_797),
	.C2V_3 (C2V_211_797),
	.L (L_797),
	.V2C_1 (V2C_797_35),
	.V2C_2 (V2C_797_192),
	.V2C_3 (V2C_797_211),
	.V (V_797)
);

VNU_3 #(quan_width) VNU798 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_798),
	.C2V_2 (C2V_198_798),
	.C2V_3 (C2V_217_798),
	.L (L_798),
	.V2C_1 (V2C_798_41),
	.V2C_2 (V2C_798_198),
	.V2C_3 (V2C_798_217),
	.V (V_798)
);

VNU_3 #(quan_width) VNU799 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_799),
	.C2V_2 (C2V_204_799),
	.C2V_3 (C2V_223_799),
	.L (L_799),
	.V2C_1 (V2C_799_47),
	.V2C_2 (V2C_799_204),
	.V2C_3 (V2C_799_223),
	.V (V_799)
);

VNU_3 #(quan_width) VNU800 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_800),
	.C2V_2 (C2V_210_800),
	.C2V_3 (C2V_229_800),
	.L (L_800),
	.V2C_1 (V2C_800_53),
	.V2C_2 (V2C_800_210),
	.V2C_3 (V2C_800_229),
	.V (V_800)
);

VNU_3 #(quan_width) VNU801 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_59_801),
	.C2V_2 (C2V_216_801),
	.C2V_3 (C2V_235_801),
	.L (L_801),
	.V2C_1 (V2C_801_59),
	.V2C_2 (V2C_801_216),
	.V2C_3 (V2C_801_235),
	.V (V_801)
);

VNU_3 #(quan_width) VNU802 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_65_802),
	.C2V_2 (C2V_222_802),
	.C2V_3 (C2V_241_802),
	.L (L_802),
	.V2C_1 (V2C_802_65),
	.V2C_2 (V2C_802_222),
	.V2C_3 (V2C_802_241),
	.V (V_802)
);

VNU_3 #(quan_width) VNU803 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_71_803),
	.C2V_2 (C2V_228_803),
	.C2V_3 (C2V_247_803),
	.L (L_803),
	.V2C_1 (V2C_803_71),
	.V2C_2 (V2C_803_228),
	.V2C_3 (V2C_803_247),
	.V (V_803)
);

VNU_3 #(quan_width) VNU804 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_77_804),
	.C2V_2 (C2V_234_804),
	.C2V_3 (C2V_253_804),
	.L (L_804),
	.V2C_1 (V2C_804_77),
	.V2C_2 (V2C_804_234),
	.V2C_3 (V2C_804_253),
	.V (V_804)
);

VNU_3 #(quan_width) VNU805 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_83_805),
	.C2V_2 (C2V_240_805),
	.C2V_3 (C2V_259_805),
	.L (L_805),
	.V2C_1 (V2C_805_83),
	.V2C_2 (V2C_805_240),
	.V2C_3 (V2C_805_259),
	.V (V_805)
);

VNU_3 #(quan_width) VNU806 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_89_806),
	.C2V_2 (C2V_246_806),
	.C2V_3 (C2V_265_806),
	.L (L_806),
	.V2C_1 (V2C_806_89),
	.V2C_2 (V2C_806_246),
	.V2C_3 (V2C_806_265),
	.V (V_806)
);

VNU_3 #(quan_width) VNU807 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_95_807),
	.C2V_2 (C2V_252_807),
	.C2V_3 (C2V_271_807),
	.L (L_807),
	.V2C_1 (V2C_807_95),
	.V2C_2 (V2C_807_252),
	.V2C_3 (V2C_807_271),
	.V (V_807)
);

VNU_3 #(quan_width) VNU808 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_101_808),
	.C2V_2 (C2V_258_808),
	.C2V_3 (C2V_277_808),
	.L (L_808),
	.V2C_1 (V2C_808_101),
	.V2C_2 (V2C_808_258),
	.V2C_3 (V2C_808_277),
	.V (V_808)
);

VNU_3 #(quan_width) VNU809 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_107_809),
	.C2V_2 (C2V_264_809),
	.C2V_3 (C2V_283_809),
	.L (L_809),
	.V2C_1 (V2C_809_107),
	.V2C_2 (V2C_809_264),
	.V2C_3 (V2C_809_283),
	.V (V_809)
);

VNU_3 #(quan_width) VNU810 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_810),
	.C2V_2 (C2V_113_810),
	.C2V_3 (C2V_270_810),
	.L (L_810),
	.V2C_1 (V2C_810_1),
	.V2C_2 (V2C_810_113),
	.V2C_3 (V2C_810_270),
	.V (V_810)
);

VNU_3 #(quan_width) VNU811 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_811),
	.C2V_2 (C2V_119_811),
	.C2V_3 (C2V_276_811),
	.L (L_811),
	.V2C_1 (V2C_811_7),
	.V2C_2 (V2C_811_119),
	.V2C_3 (V2C_811_276),
	.V (V_811)
);

VNU_3 #(quan_width) VNU812 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_812),
	.C2V_2 (C2V_125_812),
	.C2V_3 (C2V_282_812),
	.L (L_812),
	.V2C_1 (V2C_812_13),
	.V2C_2 (V2C_812_125),
	.V2C_3 (V2C_812_282),
	.V (V_812)
);

VNU_3 #(quan_width) VNU813 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_813),
	.C2V_2 (C2V_131_813),
	.C2V_3 (C2V_288_813),
	.L (L_813),
	.V2C_1 (V2C_813_19),
	.V2C_2 (V2C_813_131),
	.V2C_3 (V2C_813_288),
	.V (V_813)
);

VNU_3 #(quan_width) VNU814 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_814),
	.C2V_2 (C2V_25_814),
	.C2V_3 (C2V_137_814),
	.L (L_814),
	.V2C_1 (V2C_814_6),
	.V2C_2 (V2C_814_25),
	.V2C_3 (V2C_814_137),
	.V (V_814)
);

VNU_3 #(quan_width) VNU815 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_815),
	.C2V_2 (C2V_31_815),
	.C2V_3 (C2V_143_815),
	.L (L_815),
	.V2C_1 (V2C_815_12),
	.V2C_2 (V2C_815_31),
	.V2C_3 (V2C_815_143),
	.V (V_815)
);

VNU_3 #(quan_width) VNU816 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_816),
	.C2V_2 (C2V_37_816),
	.C2V_3 (C2V_149_816),
	.L (L_816),
	.V2C_1 (V2C_816_18),
	.V2C_2 (V2C_816_37),
	.V2C_3 (V2C_816_149),
	.V (V_816)
);

VNU_3 #(quan_width) VNU817 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_817),
	.C2V_2 (C2V_74_817),
	.C2V_3 (C2V_144_817),
	.L (L_817),
	.V2C_1 (V2C_817_43),
	.V2C_2 (V2C_817_74),
	.V2C_3 (V2C_817_144),
	.V (V_817)
);

VNU_3 #(quan_width) VNU818 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_818),
	.C2V_2 (C2V_80_818),
	.C2V_3 (C2V_150_818),
	.L (L_818),
	.V2C_1 (V2C_818_49),
	.V2C_2 (V2C_818_80),
	.V2C_3 (V2C_818_150),
	.V (V_818)
);

VNU_3 #(quan_width) VNU819 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_819),
	.C2V_2 (C2V_86_819),
	.C2V_3 (C2V_156_819),
	.L (L_819),
	.V2C_1 (V2C_819_55),
	.V2C_2 (V2C_819_86),
	.V2C_3 (V2C_819_156),
	.V (V_819)
);

VNU_3 #(quan_width) VNU820 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_820),
	.C2V_2 (C2V_92_820),
	.C2V_3 (C2V_162_820),
	.L (L_820),
	.V2C_1 (V2C_820_61),
	.V2C_2 (V2C_820_92),
	.V2C_3 (V2C_820_162),
	.V (V_820)
);

VNU_3 #(quan_width) VNU821 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_821),
	.C2V_2 (C2V_98_821),
	.C2V_3 (C2V_168_821),
	.L (L_821),
	.V2C_1 (V2C_821_67),
	.V2C_2 (V2C_821_98),
	.V2C_3 (V2C_821_168),
	.V (V_821)
);

VNU_3 #(quan_width) VNU822 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_822),
	.C2V_2 (C2V_104_822),
	.C2V_3 (C2V_174_822),
	.L (L_822),
	.V2C_1 (V2C_822_73),
	.V2C_2 (V2C_822_104),
	.V2C_3 (V2C_822_174),
	.V (V_822)
);

VNU_3 #(quan_width) VNU823 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_823),
	.C2V_2 (C2V_110_823),
	.C2V_3 (C2V_180_823),
	.L (L_823),
	.V2C_1 (V2C_823_79),
	.V2C_2 (V2C_823_110),
	.V2C_3 (V2C_823_180),
	.V (V_823)
);

VNU_3 #(quan_width) VNU824 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_824),
	.C2V_2 (C2V_116_824),
	.C2V_3 (C2V_186_824),
	.L (L_824),
	.V2C_1 (V2C_824_85),
	.V2C_2 (V2C_824_116),
	.V2C_3 (V2C_824_186),
	.V (V_824)
);

VNU_3 #(quan_width) VNU825 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_91_825),
	.C2V_2 (C2V_122_825),
	.C2V_3 (C2V_192_825),
	.L (L_825),
	.V2C_1 (V2C_825_91),
	.V2C_2 (V2C_825_122),
	.V2C_3 (V2C_825_192),
	.V (V_825)
);

VNU_3 #(quan_width) VNU826 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_97_826),
	.C2V_2 (C2V_128_826),
	.C2V_3 (C2V_198_826),
	.L (L_826),
	.V2C_1 (V2C_826_97),
	.V2C_2 (V2C_826_128),
	.V2C_3 (V2C_826_198),
	.V (V_826)
);

VNU_3 #(quan_width) VNU827 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_103_827),
	.C2V_2 (C2V_134_827),
	.C2V_3 (C2V_204_827),
	.L (L_827),
	.V2C_1 (V2C_827_103),
	.V2C_2 (V2C_827_134),
	.V2C_3 (V2C_827_204),
	.V (V_827)
);

VNU_3 #(quan_width) VNU828 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_109_828),
	.C2V_2 (C2V_140_828),
	.C2V_3 (C2V_210_828),
	.L (L_828),
	.V2C_1 (V2C_828_109),
	.V2C_2 (V2C_828_140),
	.V2C_3 (V2C_828_210),
	.V (V_828)
);

VNU_3 #(quan_width) VNU829 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_115_829),
	.C2V_2 (C2V_146_829),
	.C2V_3 (C2V_216_829),
	.L (L_829),
	.V2C_1 (V2C_829_115),
	.V2C_2 (V2C_829_146),
	.V2C_3 (V2C_829_216),
	.V (V_829)
);

VNU_3 #(quan_width) VNU830 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_121_830),
	.C2V_2 (C2V_152_830),
	.C2V_3 (C2V_222_830),
	.L (L_830),
	.V2C_1 (V2C_830_121),
	.V2C_2 (V2C_830_152),
	.V2C_3 (V2C_830_222),
	.V (V_830)
);

VNU_3 #(quan_width) VNU831 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_127_831),
	.C2V_2 (C2V_158_831),
	.C2V_3 (C2V_228_831),
	.L (L_831),
	.V2C_1 (V2C_831_127),
	.V2C_2 (V2C_831_158),
	.V2C_3 (V2C_831_228),
	.V (V_831)
);

VNU_3 #(quan_width) VNU832 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_133_832),
	.C2V_2 (C2V_164_832),
	.C2V_3 (C2V_234_832),
	.L (L_832),
	.V2C_1 (V2C_832_133),
	.V2C_2 (V2C_832_164),
	.V2C_3 (V2C_832_234),
	.V (V_832)
);

VNU_3 #(quan_width) VNU833 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_139_833),
	.C2V_2 (C2V_170_833),
	.C2V_3 (C2V_240_833),
	.L (L_833),
	.V2C_1 (V2C_833_139),
	.V2C_2 (V2C_833_170),
	.V2C_3 (V2C_833_240),
	.V (V_833)
);

VNU_3 #(quan_width) VNU834 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_145_834),
	.C2V_2 (C2V_176_834),
	.C2V_3 (C2V_246_834),
	.L (L_834),
	.V2C_1 (V2C_834_145),
	.V2C_2 (V2C_834_176),
	.V2C_3 (V2C_834_246),
	.V (V_834)
);

VNU_3 #(quan_width) VNU835 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_151_835),
	.C2V_2 (C2V_182_835),
	.C2V_3 (C2V_252_835),
	.L (L_835),
	.V2C_1 (V2C_835_151),
	.V2C_2 (V2C_835_182),
	.V2C_3 (V2C_835_252),
	.V (V_835)
);

VNU_3 #(quan_width) VNU836 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_157_836),
	.C2V_2 (C2V_188_836),
	.C2V_3 (C2V_258_836),
	.L (L_836),
	.V2C_1 (V2C_836_157),
	.V2C_2 (V2C_836_188),
	.V2C_3 (V2C_836_258),
	.V (V_836)
);

VNU_3 #(quan_width) VNU837 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_163_837),
	.C2V_2 (C2V_194_837),
	.C2V_3 (C2V_264_837),
	.L (L_837),
	.V2C_1 (V2C_837_163),
	.V2C_2 (V2C_837_194),
	.V2C_3 (V2C_837_264),
	.V (V_837)
);

VNU_3 #(quan_width) VNU838 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_169_838),
	.C2V_2 (C2V_200_838),
	.C2V_3 (C2V_270_838),
	.L (L_838),
	.V2C_1 (V2C_838_169),
	.V2C_2 (V2C_838_200),
	.V2C_3 (V2C_838_270),
	.V (V_838)
);

VNU_3 #(quan_width) VNU839 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_175_839),
	.C2V_2 (C2V_206_839),
	.C2V_3 (C2V_276_839),
	.L (L_839),
	.V2C_1 (V2C_839_175),
	.V2C_2 (V2C_839_206),
	.V2C_3 (V2C_839_276),
	.V (V_839)
);

VNU_3 #(quan_width) VNU840 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_181_840),
	.C2V_2 (C2V_212_840),
	.C2V_3 (C2V_282_840),
	.L (L_840),
	.V2C_1 (V2C_840_181),
	.V2C_2 (V2C_840_212),
	.V2C_3 (V2C_840_282),
	.V (V_840)
);

VNU_3 #(quan_width) VNU841 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_187_841),
	.C2V_2 (C2V_218_841),
	.C2V_3 (C2V_288_841),
	.L (L_841),
	.V2C_1 (V2C_841_187),
	.V2C_2 (V2C_841_218),
	.V2C_3 (V2C_841_288),
	.V (V_841)
);

VNU_3 #(quan_width) VNU842 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_842),
	.C2V_2 (C2V_193_842),
	.C2V_3 (C2V_224_842),
	.L (L_842),
	.V2C_1 (V2C_842_6),
	.V2C_2 (V2C_842_193),
	.V2C_3 (V2C_842_224),
	.V (V_842)
);

VNU_3 #(quan_width) VNU843 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_843),
	.C2V_2 (C2V_199_843),
	.C2V_3 (C2V_230_843),
	.L (L_843),
	.V2C_1 (V2C_843_12),
	.V2C_2 (V2C_843_199),
	.V2C_3 (V2C_843_230),
	.V (V_843)
);

VNU_3 #(quan_width) VNU844 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_844),
	.C2V_2 (C2V_205_844),
	.C2V_3 (C2V_236_844),
	.L (L_844),
	.V2C_1 (V2C_844_18),
	.V2C_2 (V2C_844_205),
	.V2C_3 (V2C_844_236),
	.V (V_844)
);

VNU_3 #(quan_width) VNU845 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_845),
	.C2V_2 (C2V_211_845),
	.C2V_3 (C2V_242_845),
	.L (L_845),
	.V2C_1 (V2C_845_24),
	.V2C_2 (V2C_845_211),
	.V2C_3 (V2C_845_242),
	.V (V_845)
);

VNU_3 #(quan_width) VNU846 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_846),
	.C2V_2 (C2V_217_846),
	.C2V_3 (C2V_248_846),
	.L (L_846),
	.V2C_1 (V2C_846_30),
	.V2C_2 (V2C_846_217),
	.V2C_3 (V2C_846_248),
	.V (V_846)
);

VNU_3 #(quan_width) VNU847 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_847),
	.C2V_2 (C2V_223_847),
	.C2V_3 (C2V_254_847),
	.L (L_847),
	.V2C_1 (V2C_847_36),
	.V2C_2 (V2C_847_223),
	.V2C_3 (V2C_847_254),
	.V (V_847)
);

VNU_3 #(quan_width) VNU848 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_848),
	.C2V_2 (C2V_229_848),
	.C2V_3 (C2V_260_848),
	.L (L_848),
	.V2C_1 (V2C_848_42),
	.V2C_2 (V2C_848_229),
	.V2C_3 (V2C_848_260),
	.V (V_848)
);

VNU_3 #(quan_width) VNU849 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_849),
	.C2V_2 (C2V_235_849),
	.C2V_3 (C2V_266_849),
	.L (L_849),
	.V2C_1 (V2C_849_48),
	.V2C_2 (V2C_849_235),
	.V2C_3 (V2C_849_266),
	.V (V_849)
);

VNU_3 #(quan_width) VNU850 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_54_850),
	.C2V_2 (C2V_241_850),
	.C2V_3 (C2V_272_850),
	.L (L_850),
	.V2C_1 (V2C_850_54),
	.V2C_2 (V2C_850_241),
	.V2C_3 (V2C_850_272),
	.V (V_850)
);

VNU_3 #(quan_width) VNU851 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_60_851),
	.C2V_2 (C2V_247_851),
	.C2V_3 (C2V_278_851),
	.L (L_851),
	.V2C_1 (V2C_851_60),
	.V2C_2 (V2C_851_247),
	.V2C_3 (V2C_851_278),
	.V (V_851)
);

VNU_3 #(quan_width) VNU852 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_66_852),
	.C2V_2 (C2V_253_852),
	.C2V_3 (C2V_284_852),
	.L (L_852),
	.V2C_1 (V2C_852_66),
	.V2C_2 (V2C_852_253),
	.V2C_3 (V2C_852_284),
	.V (V_852)
);

VNU_3 #(quan_width) VNU853 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_853),
	.C2V_2 (C2V_72_853),
	.C2V_3 (C2V_259_853),
	.L (L_853),
	.V2C_1 (V2C_853_2),
	.V2C_2 (V2C_853_72),
	.V2C_3 (V2C_853_259),
	.V (V_853)
);

VNU_3 #(quan_width) VNU854 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_854),
	.C2V_2 (C2V_78_854),
	.C2V_3 (C2V_265_854),
	.L (L_854),
	.V2C_1 (V2C_854_8),
	.V2C_2 (V2C_854_78),
	.V2C_3 (V2C_854_265),
	.V (V_854)
);

VNU_3 #(quan_width) VNU855 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_855),
	.C2V_2 (C2V_84_855),
	.C2V_3 (C2V_271_855),
	.L (L_855),
	.V2C_1 (V2C_855_14),
	.V2C_2 (V2C_855_84),
	.V2C_3 (V2C_855_271),
	.V (V_855)
);

VNU_3 #(quan_width) VNU856 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_856),
	.C2V_2 (C2V_90_856),
	.C2V_3 (C2V_277_856),
	.L (L_856),
	.V2C_1 (V2C_856_20),
	.V2C_2 (V2C_856_90),
	.V2C_3 (V2C_856_277),
	.V (V_856)
);

VNU_3 #(quan_width) VNU857 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_857),
	.C2V_2 (C2V_96_857),
	.C2V_3 (C2V_283_857),
	.L (L_857),
	.V2C_1 (V2C_857_26),
	.V2C_2 (V2C_857_96),
	.V2C_3 (V2C_857_283),
	.V (V_857)
);

VNU_3 #(quan_width) VNU858 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_858),
	.C2V_2 (C2V_32_858),
	.C2V_3 (C2V_102_858),
	.L (L_858),
	.V2C_1 (V2C_858_1),
	.V2C_2 (V2C_858_32),
	.V2C_3 (V2C_858_102),
	.V (V_858)
);

VNU_3 #(quan_width) VNU859 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_859),
	.C2V_2 (C2V_38_859),
	.C2V_3 (C2V_108_859),
	.L (L_859),
	.V2C_1 (V2C_859_7),
	.V2C_2 (V2C_859_38),
	.V2C_3 (V2C_859_108),
	.V (V_859)
);

VNU_3 #(quan_width) VNU860 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_860),
	.C2V_2 (C2V_44_860),
	.C2V_3 (C2V_114_860),
	.L (L_860),
	.V2C_1 (V2C_860_13),
	.V2C_2 (V2C_860_44),
	.V2C_3 (V2C_860_114),
	.V (V_860)
);

VNU_3 #(quan_width) VNU861 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_861),
	.C2V_2 (C2V_50_861),
	.C2V_3 (C2V_120_861),
	.L (L_861),
	.V2C_1 (V2C_861_19),
	.V2C_2 (V2C_861_50),
	.V2C_3 (V2C_861_120),
	.V (V_861)
);

VNU_3 #(quan_width) VNU862 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_862),
	.C2V_2 (C2V_56_862),
	.C2V_3 (C2V_126_862),
	.L (L_862),
	.V2C_1 (V2C_862_25),
	.V2C_2 (V2C_862_56),
	.V2C_3 (V2C_862_126),
	.V (V_862)
);

VNU_3 #(quan_width) VNU863 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_863),
	.C2V_2 (C2V_62_863),
	.C2V_3 (C2V_132_863),
	.L (L_863),
	.V2C_1 (V2C_863_31),
	.V2C_2 (V2C_863_62),
	.V2C_3 (V2C_863_132),
	.V (V_863)
);

VNU_3 #(quan_width) VNU864 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_864),
	.C2V_2 (C2V_68_864),
	.C2V_3 (C2V_138_864),
	.L (L_864),
	.V2C_1 (V2C_864_37),
	.V2C_2 (V2C_864_68),
	.V2C_3 (V2C_864_138),
	.V (V_864)
);

VNU_6 #(quan_width) VNU865 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_865),
	.C2V_2 (C2V_85_865),
	.C2V_3 (C2V_87_865),
	.C2V_4 (C2V_110_865),
	.C2V_5 (C2V_234_865),
	.C2V_6 (C2V_263_865),
	.L (L_865),
	.V2C_1 (V2C_865_64),
	.V2C_2 (V2C_865_85),
	.V2C_3 (V2C_865_87),
	.V2C_4 (V2C_865_110),
	.V2C_5 (V2C_865_234),
	.V2C_6 (V2C_865_263),
	.V (V_865)
);

VNU_6 #(quan_width) VNU866 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_866),
	.C2V_2 (C2V_91_866),
	.C2V_3 (C2V_93_866),
	.C2V_4 (C2V_116_866),
	.C2V_5 (C2V_240_866),
	.C2V_6 (C2V_269_866),
	.L (L_866),
	.V2C_1 (V2C_866_70),
	.V2C_2 (V2C_866_91),
	.V2C_3 (V2C_866_93),
	.V2C_4 (V2C_866_116),
	.V2C_5 (V2C_866_240),
	.V2C_6 (V2C_866_269),
	.V (V_866)
);

VNU_6 #(quan_width) VNU867 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_867),
	.C2V_2 (C2V_97_867),
	.C2V_3 (C2V_99_867),
	.C2V_4 (C2V_122_867),
	.C2V_5 (C2V_246_867),
	.C2V_6 (C2V_275_867),
	.L (L_867),
	.V2C_1 (V2C_867_76),
	.V2C_2 (V2C_867_97),
	.V2C_3 (V2C_867_99),
	.V2C_4 (V2C_867_122),
	.V2C_5 (V2C_867_246),
	.V2C_6 (V2C_867_275),
	.V (V_867)
);

VNU_6 #(quan_width) VNU868 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_868),
	.C2V_2 (C2V_103_868),
	.C2V_3 (C2V_105_868),
	.C2V_4 (C2V_128_868),
	.C2V_5 (C2V_252_868),
	.C2V_6 (C2V_281_868),
	.L (L_868),
	.V2C_1 (V2C_868_82),
	.V2C_2 (V2C_868_103),
	.V2C_3 (V2C_868_105),
	.V2C_4 (V2C_868_128),
	.V2C_5 (V2C_868_252),
	.V2C_6 (V2C_868_281),
	.V (V_868)
);

VNU_6 #(quan_width) VNU869 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_869),
	.C2V_2 (C2V_109_869),
	.C2V_3 (C2V_111_869),
	.C2V_4 (C2V_134_869),
	.C2V_5 (C2V_258_869),
	.C2V_6 (C2V_287_869),
	.L (L_869),
	.V2C_1 (V2C_869_88),
	.V2C_2 (V2C_869_109),
	.V2C_3 (V2C_869_111),
	.V2C_4 (V2C_869_134),
	.V2C_5 (V2C_869_258),
	.V2C_6 (V2C_869_287),
	.V (V_869)
);

VNU_6 #(quan_width) VNU870 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_870),
	.C2V_2 (C2V_94_870),
	.C2V_3 (C2V_115_870),
	.C2V_4 (C2V_117_870),
	.C2V_5 (C2V_140_870),
	.C2V_6 (C2V_264_870),
	.L (L_870),
	.V2C_1 (V2C_870_5),
	.V2C_2 (V2C_870_94),
	.V2C_3 (V2C_870_115),
	.V2C_4 (V2C_870_117),
	.V2C_5 (V2C_870_140),
	.V2C_6 (V2C_870_264),
	.V (V_870)
);

VNU_6 #(quan_width) VNU871 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_871),
	.C2V_2 (C2V_100_871),
	.C2V_3 (C2V_121_871),
	.C2V_4 (C2V_123_871),
	.C2V_5 (C2V_146_871),
	.C2V_6 (C2V_270_871),
	.L (L_871),
	.V2C_1 (V2C_871_11),
	.V2C_2 (V2C_871_100),
	.V2C_3 (V2C_871_121),
	.V2C_4 (V2C_871_123),
	.V2C_5 (V2C_871_146),
	.V2C_6 (V2C_871_270),
	.V (V_871)
);

VNU_6 #(quan_width) VNU872 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_872),
	.C2V_2 (C2V_106_872),
	.C2V_3 (C2V_127_872),
	.C2V_4 (C2V_129_872),
	.C2V_5 (C2V_152_872),
	.C2V_6 (C2V_276_872),
	.L (L_872),
	.V2C_1 (V2C_872_17),
	.V2C_2 (V2C_872_106),
	.V2C_3 (V2C_872_127),
	.V2C_4 (V2C_872_129),
	.V2C_5 (V2C_872_152),
	.V2C_6 (V2C_872_276),
	.V (V_872)
);

VNU_6 #(quan_width) VNU873 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_873),
	.C2V_2 (C2V_112_873),
	.C2V_3 (C2V_133_873),
	.C2V_4 (C2V_135_873),
	.C2V_5 (C2V_158_873),
	.C2V_6 (C2V_282_873),
	.L (L_873),
	.V2C_1 (V2C_873_23),
	.V2C_2 (V2C_873_112),
	.V2C_3 (V2C_873_133),
	.V2C_4 (V2C_873_135),
	.V2C_5 (V2C_873_158),
	.V2C_6 (V2C_873_282),
	.V (V_873)
);

VNU_6 #(quan_width) VNU874 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_874),
	.C2V_2 (C2V_118_874),
	.C2V_3 (C2V_139_874),
	.C2V_4 (C2V_141_874),
	.C2V_5 (C2V_164_874),
	.C2V_6 (C2V_288_874),
	.L (L_874),
	.V2C_1 (V2C_874_29),
	.V2C_2 (V2C_874_118),
	.V2C_3 (V2C_874_139),
	.V2C_4 (V2C_874_141),
	.V2C_5 (V2C_874_164),
	.V2C_6 (V2C_874_288),
	.V (V_874)
);

VNU_6 #(quan_width) VNU875 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_875),
	.C2V_2 (C2V_35_875),
	.C2V_3 (C2V_124_875),
	.C2V_4 (C2V_145_875),
	.C2V_5 (C2V_147_875),
	.C2V_6 (C2V_170_875),
	.L (L_875),
	.V2C_1 (V2C_875_6),
	.V2C_2 (V2C_875_35),
	.V2C_3 (V2C_875_124),
	.V2C_4 (V2C_875_145),
	.V2C_5 (V2C_875_147),
	.V2C_6 (V2C_875_170),
	.V (V_875)
);

VNU_6 #(quan_width) VNU876 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_876),
	.C2V_2 (C2V_41_876),
	.C2V_3 (C2V_130_876),
	.C2V_4 (C2V_151_876),
	.C2V_5 (C2V_153_876),
	.C2V_6 (C2V_176_876),
	.L (L_876),
	.V2C_1 (V2C_876_12),
	.V2C_2 (V2C_876_41),
	.V2C_3 (V2C_876_130),
	.V2C_4 (V2C_876_151),
	.V2C_5 (V2C_876_153),
	.V2C_6 (V2C_876_176),
	.V (V_876)
);

VNU_6 #(quan_width) VNU877 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_877),
	.C2V_2 (C2V_47_877),
	.C2V_3 (C2V_136_877),
	.C2V_4 (C2V_157_877),
	.C2V_5 (C2V_159_877),
	.C2V_6 (C2V_182_877),
	.L (L_877),
	.V2C_1 (V2C_877_18),
	.V2C_2 (V2C_877_47),
	.V2C_3 (V2C_877_136),
	.V2C_4 (V2C_877_157),
	.V2C_5 (V2C_877_159),
	.V2C_6 (V2C_877_182),
	.V (V_877)
);

VNU_6 #(quan_width) VNU878 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_878),
	.C2V_2 (C2V_53_878),
	.C2V_3 (C2V_142_878),
	.C2V_4 (C2V_163_878),
	.C2V_5 (C2V_165_878),
	.C2V_6 (C2V_188_878),
	.L (L_878),
	.V2C_1 (V2C_878_24),
	.V2C_2 (V2C_878_53),
	.V2C_3 (V2C_878_142),
	.V2C_4 (V2C_878_163),
	.V2C_5 (V2C_878_165),
	.V2C_6 (V2C_878_188),
	.V (V_878)
);

VNU_6 #(quan_width) VNU879 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_879),
	.C2V_2 (C2V_59_879),
	.C2V_3 (C2V_148_879),
	.C2V_4 (C2V_169_879),
	.C2V_5 (C2V_171_879),
	.C2V_6 (C2V_194_879),
	.L (L_879),
	.V2C_1 (V2C_879_30),
	.V2C_2 (V2C_879_59),
	.V2C_3 (V2C_879_148),
	.V2C_4 (V2C_879_169),
	.V2C_5 (V2C_879_171),
	.V2C_6 (V2C_879_194),
	.V (V_879)
);

VNU_6 #(quan_width) VNU880 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_880),
	.C2V_2 (C2V_65_880),
	.C2V_3 (C2V_154_880),
	.C2V_4 (C2V_175_880),
	.C2V_5 (C2V_177_880),
	.C2V_6 (C2V_200_880),
	.L (L_880),
	.V2C_1 (V2C_880_36),
	.V2C_2 (V2C_880_65),
	.V2C_3 (V2C_880_154),
	.V2C_4 (V2C_880_175),
	.V2C_5 (V2C_880_177),
	.V2C_6 (V2C_880_200),
	.V (V_880)
);

VNU_6 #(quan_width) VNU881 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_881),
	.C2V_2 (C2V_71_881),
	.C2V_3 (C2V_160_881),
	.C2V_4 (C2V_181_881),
	.C2V_5 (C2V_183_881),
	.C2V_6 (C2V_206_881),
	.L (L_881),
	.V2C_1 (V2C_881_42),
	.V2C_2 (V2C_881_71),
	.V2C_3 (V2C_881_160),
	.V2C_4 (V2C_881_181),
	.V2C_5 (V2C_881_183),
	.V2C_6 (V2C_881_206),
	.V (V_881)
);

VNU_6 #(quan_width) VNU882 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_882),
	.C2V_2 (C2V_77_882),
	.C2V_3 (C2V_166_882),
	.C2V_4 (C2V_187_882),
	.C2V_5 (C2V_189_882),
	.C2V_6 (C2V_212_882),
	.L (L_882),
	.V2C_1 (V2C_882_48),
	.V2C_2 (V2C_882_77),
	.V2C_3 (V2C_882_166),
	.V2C_4 (V2C_882_187),
	.V2C_5 (V2C_882_189),
	.V2C_6 (V2C_882_212),
	.V (V_882)
);

VNU_6 #(quan_width) VNU883 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_54_883),
	.C2V_2 (C2V_83_883),
	.C2V_3 (C2V_172_883),
	.C2V_4 (C2V_193_883),
	.C2V_5 (C2V_195_883),
	.C2V_6 (C2V_218_883),
	.L (L_883),
	.V2C_1 (V2C_883_54),
	.V2C_2 (V2C_883_83),
	.V2C_3 (V2C_883_172),
	.V2C_4 (V2C_883_193),
	.V2C_5 (V2C_883_195),
	.V2C_6 (V2C_883_218),
	.V (V_883)
);

VNU_6 #(quan_width) VNU884 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_60_884),
	.C2V_2 (C2V_89_884),
	.C2V_3 (C2V_178_884),
	.C2V_4 (C2V_199_884),
	.C2V_5 (C2V_201_884),
	.C2V_6 (C2V_224_884),
	.L (L_884),
	.V2C_1 (V2C_884_60),
	.V2C_2 (V2C_884_89),
	.V2C_3 (V2C_884_178),
	.V2C_4 (V2C_884_199),
	.V2C_5 (V2C_884_201),
	.V2C_6 (V2C_884_224),
	.V (V_884)
);

VNU_6 #(quan_width) VNU885 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_66_885),
	.C2V_2 (C2V_95_885),
	.C2V_3 (C2V_184_885),
	.C2V_4 (C2V_205_885),
	.C2V_5 (C2V_207_885),
	.C2V_6 (C2V_230_885),
	.L (L_885),
	.V2C_1 (V2C_885_66),
	.V2C_2 (V2C_885_95),
	.V2C_3 (V2C_885_184),
	.V2C_4 (V2C_885_205),
	.V2C_5 (V2C_885_207),
	.V2C_6 (V2C_885_230),
	.V (V_885)
);

VNU_6 #(quan_width) VNU886 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_72_886),
	.C2V_2 (C2V_101_886),
	.C2V_3 (C2V_190_886),
	.C2V_4 (C2V_211_886),
	.C2V_5 (C2V_213_886),
	.C2V_6 (C2V_236_886),
	.L (L_886),
	.V2C_1 (V2C_886_72),
	.V2C_2 (V2C_886_101),
	.V2C_3 (V2C_886_190),
	.V2C_4 (V2C_886_211),
	.V2C_5 (V2C_886_213),
	.V2C_6 (V2C_886_236),
	.V (V_886)
);

VNU_6 #(quan_width) VNU887 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_78_887),
	.C2V_2 (C2V_107_887),
	.C2V_3 (C2V_196_887),
	.C2V_4 (C2V_217_887),
	.C2V_5 (C2V_219_887),
	.C2V_6 (C2V_242_887),
	.L (L_887),
	.V2C_1 (V2C_887_78),
	.V2C_2 (V2C_887_107),
	.V2C_3 (V2C_887_196),
	.V2C_4 (V2C_887_217),
	.V2C_5 (V2C_887_219),
	.V2C_6 (V2C_887_242),
	.V (V_887)
);

VNU_6 #(quan_width) VNU888 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_84_888),
	.C2V_2 (C2V_113_888),
	.C2V_3 (C2V_202_888),
	.C2V_4 (C2V_223_888),
	.C2V_5 (C2V_225_888),
	.C2V_6 (C2V_248_888),
	.L (L_888),
	.V2C_1 (V2C_888_84),
	.V2C_2 (V2C_888_113),
	.V2C_3 (V2C_888_202),
	.V2C_4 (V2C_888_223),
	.V2C_5 (V2C_888_225),
	.V2C_6 (V2C_888_248),
	.V (V_888)
);

VNU_6 #(quan_width) VNU889 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_90_889),
	.C2V_2 (C2V_119_889),
	.C2V_3 (C2V_208_889),
	.C2V_4 (C2V_229_889),
	.C2V_5 (C2V_231_889),
	.C2V_6 (C2V_254_889),
	.L (L_889),
	.V2C_1 (V2C_889_90),
	.V2C_2 (V2C_889_119),
	.V2C_3 (V2C_889_208),
	.V2C_4 (V2C_889_229),
	.V2C_5 (V2C_889_231),
	.V2C_6 (V2C_889_254),
	.V (V_889)
);

VNU_6 #(quan_width) VNU890 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_96_890),
	.C2V_2 (C2V_125_890),
	.C2V_3 (C2V_214_890),
	.C2V_4 (C2V_235_890),
	.C2V_5 (C2V_237_890),
	.C2V_6 (C2V_260_890),
	.L (L_890),
	.V2C_1 (V2C_890_96),
	.V2C_2 (V2C_890_125),
	.V2C_3 (V2C_890_214),
	.V2C_4 (V2C_890_235),
	.V2C_5 (V2C_890_237),
	.V2C_6 (V2C_890_260),
	.V (V_890)
);

VNU_6 #(quan_width) VNU891 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_102_891),
	.C2V_2 (C2V_131_891),
	.C2V_3 (C2V_220_891),
	.C2V_4 (C2V_241_891),
	.C2V_5 (C2V_243_891),
	.C2V_6 (C2V_266_891),
	.L (L_891),
	.V2C_1 (V2C_891_102),
	.V2C_2 (V2C_891_131),
	.V2C_3 (V2C_891_220),
	.V2C_4 (V2C_891_241),
	.V2C_5 (V2C_891_243),
	.V2C_6 (V2C_891_266),
	.V (V_891)
);

VNU_6 #(quan_width) VNU892 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_108_892),
	.C2V_2 (C2V_137_892),
	.C2V_3 (C2V_226_892),
	.C2V_4 (C2V_247_892),
	.C2V_5 (C2V_249_892),
	.C2V_6 (C2V_272_892),
	.L (L_892),
	.V2C_1 (V2C_892_108),
	.V2C_2 (V2C_892_137),
	.V2C_3 (V2C_892_226),
	.V2C_4 (V2C_892_247),
	.V2C_5 (V2C_892_249),
	.V2C_6 (V2C_892_272),
	.V (V_892)
);

VNU_6 #(quan_width) VNU893 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_114_893),
	.C2V_2 (C2V_143_893),
	.C2V_3 (C2V_232_893),
	.C2V_4 (C2V_253_893),
	.C2V_5 (C2V_255_893),
	.C2V_6 (C2V_278_893),
	.L (L_893),
	.V2C_1 (V2C_893_114),
	.V2C_2 (V2C_893_143),
	.V2C_3 (V2C_893_232),
	.V2C_4 (V2C_893_253),
	.V2C_5 (V2C_893_255),
	.V2C_6 (V2C_893_278),
	.V (V_893)
);

VNU_6 #(quan_width) VNU894 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_120_894),
	.C2V_2 (C2V_149_894),
	.C2V_3 (C2V_238_894),
	.C2V_4 (C2V_259_894),
	.C2V_5 (C2V_261_894),
	.C2V_6 (C2V_284_894),
	.L (L_894),
	.V2C_1 (V2C_894_120),
	.V2C_2 (V2C_894_149),
	.V2C_3 (V2C_894_238),
	.V2C_4 (V2C_894_259),
	.V2C_5 (V2C_894_261),
	.V2C_6 (V2C_894_284),
	.V (V_894)
);

VNU_6 #(quan_width) VNU895 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_895),
	.C2V_2 (C2V_126_895),
	.C2V_3 (C2V_155_895),
	.C2V_4 (C2V_244_895),
	.C2V_5 (C2V_265_895),
	.C2V_6 (C2V_267_895),
	.L (L_895),
	.V2C_1 (V2C_895_2),
	.V2C_2 (V2C_895_126),
	.V2C_3 (V2C_895_155),
	.V2C_4 (V2C_895_244),
	.V2C_5 (V2C_895_265),
	.V2C_6 (V2C_895_267),
	.V (V_895)
);

VNU_6 #(quan_width) VNU896 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_896),
	.C2V_2 (C2V_132_896),
	.C2V_3 (C2V_161_896),
	.C2V_4 (C2V_250_896),
	.C2V_5 (C2V_271_896),
	.C2V_6 (C2V_273_896),
	.L (L_896),
	.V2C_1 (V2C_896_8),
	.V2C_2 (V2C_896_132),
	.V2C_3 (V2C_896_161),
	.V2C_4 (V2C_896_250),
	.V2C_5 (V2C_896_271),
	.V2C_6 (V2C_896_273),
	.V (V_896)
);

VNU_6 #(quan_width) VNU897 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_897),
	.C2V_2 (C2V_138_897),
	.C2V_3 (C2V_167_897),
	.C2V_4 (C2V_256_897),
	.C2V_5 (C2V_277_897),
	.C2V_6 (C2V_279_897),
	.L (L_897),
	.V2C_1 (V2C_897_14),
	.V2C_2 (V2C_897_138),
	.V2C_3 (V2C_897_167),
	.V2C_4 (V2C_897_256),
	.V2C_5 (V2C_897_277),
	.V2C_6 (V2C_897_279),
	.V (V_897)
);

VNU_6 #(quan_width) VNU898 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_898),
	.C2V_2 (C2V_144_898),
	.C2V_3 (C2V_173_898),
	.C2V_4 (C2V_262_898),
	.C2V_5 (C2V_283_898),
	.C2V_6 (C2V_285_898),
	.L (L_898),
	.V2C_1 (V2C_898_20),
	.V2C_2 (V2C_898_144),
	.V2C_3 (V2C_898_173),
	.V2C_4 (V2C_898_262),
	.V2C_5 (V2C_898_283),
	.V2C_6 (V2C_898_285),
	.V (V_898)
);

VNU_6 #(quan_width) VNU899 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_899),
	.C2V_2 (C2V_3_899),
	.C2V_3 (C2V_26_899),
	.C2V_4 (C2V_150_899),
	.C2V_5 (C2V_179_899),
	.C2V_6 (C2V_268_899),
	.L (L_899),
	.V2C_1 (V2C_899_1),
	.V2C_2 (V2C_899_3),
	.V2C_3 (V2C_899_26),
	.V2C_4 (V2C_899_150),
	.V2C_5 (V2C_899_179),
	.V2C_6 (V2C_899_268),
	.V (V_899)
);

VNU_6 #(quan_width) VNU900 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_900),
	.C2V_2 (C2V_9_900),
	.C2V_3 (C2V_32_900),
	.C2V_4 (C2V_156_900),
	.C2V_5 (C2V_185_900),
	.C2V_6 (C2V_274_900),
	.L (L_900),
	.V2C_1 (V2C_900_7),
	.V2C_2 (V2C_900_9),
	.V2C_3 (V2C_900_32),
	.V2C_4 (V2C_900_156),
	.V2C_5 (V2C_900_185),
	.V2C_6 (V2C_900_274),
	.V (V_900)
);

VNU_6 #(quan_width) VNU901 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_901),
	.C2V_2 (C2V_15_901),
	.C2V_3 (C2V_38_901),
	.C2V_4 (C2V_162_901),
	.C2V_5 (C2V_191_901),
	.C2V_6 (C2V_280_901),
	.L (L_901),
	.V2C_1 (V2C_901_13),
	.V2C_2 (V2C_901_15),
	.V2C_3 (V2C_901_38),
	.V2C_4 (V2C_901_162),
	.V2C_5 (V2C_901_191),
	.V2C_6 (V2C_901_280),
	.V (V_901)
);

VNU_6 #(quan_width) VNU902 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_902),
	.C2V_2 (C2V_21_902),
	.C2V_3 (C2V_44_902),
	.C2V_4 (C2V_168_902),
	.C2V_5 (C2V_197_902),
	.C2V_6 (C2V_286_902),
	.L (L_902),
	.V2C_1 (V2C_902_19),
	.V2C_2 (V2C_902_21),
	.V2C_3 (V2C_902_44),
	.V2C_4 (V2C_902_168),
	.V2C_5 (V2C_902_197),
	.V2C_6 (V2C_902_286),
	.V (V_902)
);

VNU_6 #(quan_width) VNU903 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_903),
	.C2V_2 (C2V_25_903),
	.C2V_3 (C2V_27_903),
	.C2V_4 (C2V_50_903),
	.C2V_5 (C2V_174_903),
	.C2V_6 (C2V_203_903),
	.L (L_903),
	.V2C_1 (V2C_903_4),
	.V2C_2 (V2C_903_25),
	.V2C_3 (V2C_903_27),
	.V2C_4 (V2C_903_50),
	.V2C_5 (V2C_903_174),
	.V2C_6 (V2C_903_203),
	.V (V_903)
);

VNU_6 #(quan_width) VNU904 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_904),
	.C2V_2 (C2V_31_904),
	.C2V_3 (C2V_33_904),
	.C2V_4 (C2V_56_904),
	.C2V_5 (C2V_180_904),
	.C2V_6 (C2V_209_904),
	.L (L_904),
	.V2C_1 (V2C_904_10),
	.V2C_2 (V2C_904_31),
	.V2C_3 (V2C_904_33),
	.V2C_4 (V2C_904_56),
	.V2C_5 (V2C_904_180),
	.V2C_6 (V2C_904_209),
	.V (V_904)
);

VNU_6 #(quan_width) VNU905 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_905),
	.C2V_2 (C2V_37_905),
	.C2V_3 (C2V_39_905),
	.C2V_4 (C2V_62_905),
	.C2V_5 (C2V_186_905),
	.C2V_6 (C2V_215_905),
	.L (L_905),
	.V2C_1 (V2C_905_16),
	.V2C_2 (V2C_905_37),
	.V2C_3 (V2C_905_39),
	.V2C_4 (V2C_905_62),
	.V2C_5 (V2C_905_186),
	.V2C_6 (V2C_905_215),
	.V (V_905)
);

VNU_6 #(quan_width) VNU906 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_906),
	.C2V_2 (C2V_43_906),
	.C2V_3 (C2V_45_906),
	.C2V_4 (C2V_68_906),
	.C2V_5 (C2V_192_906),
	.C2V_6 (C2V_221_906),
	.L (L_906),
	.V2C_1 (V2C_906_22),
	.V2C_2 (V2C_906_43),
	.V2C_3 (V2C_906_45),
	.V2C_4 (V2C_906_68),
	.V2C_5 (V2C_906_192),
	.V2C_6 (V2C_906_221),
	.V (V_906)
);

VNU_6 #(quan_width) VNU907 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_907),
	.C2V_2 (C2V_49_907),
	.C2V_3 (C2V_51_907),
	.C2V_4 (C2V_74_907),
	.C2V_5 (C2V_198_907),
	.C2V_6 (C2V_227_907),
	.L (L_907),
	.V2C_1 (V2C_907_28),
	.V2C_2 (V2C_907_49),
	.V2C_3 (V2C_907_51),
	.V2C_4 (V2C_907_74),
	.V2C_5 (V2C_907_198),
	.V2C_6 (V2C_907_227),
	.V (V_907)
);

VNU_6 #(quan_width) VNU908 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_908),
	.C2V_2 (C2V_55_908),
	.C2V_3 (C2V_57_908),
	.C2V_4 (C2V_80_908),
	.C2V_5 (C2V_204_908),
	.C2V_6 (C2V_233_908),
	.L (L_908),
	.V2C_1 (V2C_908_34),
	.V2C_2 (V2C_908_55),
	.V2C_3 (V2C_908_57),
	.V2C_4 (V2C_908_80),
	.V2C_5 (V2C_908_204),
	.V2C_6 (V2C_908_233),
	.V (V_908)
);

VNU_6 #(quan_width) VNU909 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_909),
	.C2V_2 (C2V_61_909),
	.C2V_3 (C2V_63_909),
	.C2V_4 (C2V_86_909),
	.C2V_5 (C2V_210_909),
	.C2V_6 (C2V_239_909),
	.L (L_909),
	.V2C_1 (V2C_909_40),
	.V2C_2 (V2C_909_61),
	.V2C_3 (V2C_909_63),
	.V2C_4 (V2C_909_86),
	.V2C_5 (V2C_909_210),
	.V2C_6 (V2C_909_239),
	.V (V_909)
);

VNU_6 #(quan_width) VNU910 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_910),
	.C2V_2 (C2V_67_910),
	.C2V_3 (C2V_69_910),
	.C2V_4 (C2V_92_910),
	.C2V_5 (C2V_216_910),
	.C2V_6 (C2V_245_910),
	.L (L_910),
	.V2C_1 (V2C_910_46),
	.V2C_2 (V2C_910_67),
	.V2C_3 (V2C_910_69),
	.V2C_4 (V2C_910_92),
	.V2C_5 (V2C_910_216),
	.V2C_6 (V2C_910_245),
	.V (V_910)
);

VNU_6 #(quan_width) VNU911 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_911),
	.C2V_2 (C2V_73_911),
	.C2V_3 (C2V_75_911),
	.C2V_4 (C2V_98_911),
	.C2V_5 (C2V_222_911),
	.C2V_6 (C2V_251_911),
	.L (L_911),
	.V2C_1 (V2C_911_52),
	.V2C_2 (V2C_911_73),
	.V2C_3 (V2C_911_75),
	.V2C_4 (V2C_911_98),
	.V2C_5 (V2C_911_222),
	.V2C_6 (V2C_911_251),
	.V (V_911)
);

VNU_6 #(quan_width) VNU912 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_912),
	.C2V_2 (C2V_79_912),
	.C2V_3 (C2V_81_912),
	.C2V_4 (C2V_104_912),
	.C2V_5 (C2V_228_912),
	.C2V_6 (C2V_257_912),
	.L (L_912),
	.V2C_1 (V2C_912_58),
	.V2C_2 (V2C_912_79),
	.V2C_3 (V2C_912_81),
	.V2C_4 (V2C_912_104),
	.V2C_5 (V2C_912_228),
	.V2C_6 (V2C_912_257),
	.V (V_912)
);

VNU_6 #(quan_width) VNU913 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_913),
	.C2V_2 (C2V_111_913),
	.C2V_3 (C2V_127_913),
	.C2V_4 (C2V_150_913),
	.C2V_5 (C2V_208_913),
	.C2V_6 (C2V_263_913),
	.L (L_913),
	.V2C_1 (V2C_913_20),
	.V2C_2 (V2C_913_111),
	.V2C_3 (V2C_913_127),
	.V2C_4 (V2C_913_150),
	.V2C_5 (V2C_913_208),
	.V2C_6 (V2C_913_263),
	.V (V_913)
);

VNU_6 #(quan_width) VNU914 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_914),
	.C2V_2 (C2V_117_914),
	.C2V_3 (C2V_133_914),
	.C2V_4 (C2V_156_914),
	.C2V_5 (C2V_214_914),
	.C2V_6 (C2V_269_914),
	.L (L_914),
	.V2C_1 (V2C_914_26),
	.V2C_2 (V2C_914_117),
	.V2C_3 (V2C_914_133),
	.V2C_4 (V2C_914_156),
	.V2C_5 (V2C_914_214),
	.V2C_6 (V2C_914_269),
	.V (V_914)
);

VNU_6 #(quan_width) VNU915 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_915),
	.C2V_2 (C2V_123_915),
	.C2V_3 (C2V_139_915),
	.C2V_4 (C2V_162_915),
	.C2V_5 (C2V_220_915),
	.C2V_6 (C2V_275_915),
	.L (L_915),
	.V2C_1 (V2C_915_32),
	.V2C_2 (V2C_915_123),
	.V2C_3 (V2C_915_139),
	.V2C_4 (V2C_915_162),
	.V2C_5 (V2C_915_220),
	.V2C_6 (V2C_915_275),
	.V (V_915)
);

VNU_6 #(quan_width) VNU916 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_916),
	.C2V_2 (C2V_129_916),
	.C2V_3 (C2V_145_916),
	.C2V_4 (C2V_168_916),
	.C2V_5 (C2V_226_916),
	.C2V_6 (C2V_281_916),
	.L (L_916),
	.V2C_1 (V2C_916_38),
	.V2C_2 (V2C_916_129),
	.V2C_3 (V2C_916_145),
	.V2C_4 (V2C_916_168),
	.V2C_5 (V2C_916_226),
	.V2C_6 (V2C_916_281),
	.V (V_916)
);

VNU_6 #(quan_width) VNU917 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_917),
	.C2V_2 (C2V_135_917),
	.C2V_3 (C2V_151_917),
	.C2V_4 (C2V_174_917),
	.C2V_5 (C2V_232_917),
	.C2V_6 (C2V_287_917),
	.L (L_917),
	.V2C_1 (V2C_917_44),
	.V2C_2 (V2C_917_135),
	.V2C_3 (V2C_917_151),
	.V2C_4 (V2C_917_174),
	.V2C_5 (V2C_917_232),
	.V2C_6 (V2C_917_287),
	.V (V_917)
);

VNU_6 #(quan_width) VNU918 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_918),
	.C2V_2 (C2V_50_918),
	.C2V_3 (C2V_141_918),
	.C2V_4 (C2V_157_918),
	.C2V_5 (C2V_180_918),
	.C2V_6 (C2V_238_918),
	.L (L_918),
	.V2C_1 (V2C_918_5),
	.V2C_2 (V2C_918_50),
	.V2C_3 (V2C_918_141),
	.V2C_4 (V2C_918_157),
	.V2C_5 (V2C_918_180),
	.V2C_6 (V2C_918_238),
	.V (V_918)
);

VNU_6 #(quan_width) VNU919 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_919),
	.C2V_2 (C2V_56_919),
	.C2V_3 (C2V_147_919),
	.C2V_4 (C2V_163_919),
	.C2V_5 (C2V_186_919),
	.C2V_6 (C2V_244_919),
	.L (L_919),
	.V2C_1 (V2C_919_11),
	.V2C_2 (V2C_919_56),
	.V2C_3 (V2C_919_147),
	.V2C_4 (V2C_919_163),
	.V2C_5 (V2C_919_186),
	.V2C_6 (V2C_919_244),
	.V (V_919)
);

VNU_6 #(quan_width) VNU920 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_920),
	.C2V_2 (C2V_62_920),
	.C2V_3 (C2V_153_920),
	.C2V_4 (C2V_169_920),
	.C2V_5 (C2V_192_920),
	.C2V_6 (C2V_250_920),
	.L (L_920),
	.V2C_1 (V2C_920_17),
	.V2C_2 (V2C_920_62),
	.V2C_3 (V2C_920_153),
	.V2C_4 (V2C_920_169),
	.V2C_5 (V2C_920_192),
	.V2C_6 (V2C_920_250),
	.V (V_920)
);

VNU_6 #(quan_width) VNU921 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_921),
	.C2V_2 (C2V_68_921),
	.C2V_3 (C2V_159_921),
	.C2V_4 (C2V_175_921),
	.C2V_5 (C2V_198_921),
	.C2V_6 (C2V_256_921),
	.L (L_921),
	.V2C_1 (V2C_921_23),
	.V2C_2 (V2C_921_68),
	.V2C_3 (V2C_921_159),
	.V2C_4 (V2C_921_175),
	.V2C_5 (V2C_921_198),
	.V2C_6 (V2C_921_256),
	.V (V_921)
);

VNU_6 #(quan_width) VNU922 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_922),
	.C2V_2 (C2V_74_922),
	.C2V_3 (C2V_165_922),
	.C2V_4 (C2V_181_922),
	.C2V_5 (C2V_204_922),
	.C2V_6 (C2V_262_922),
	.L (L_922),
	.V2C_1 (V2C_922_29),
	.V2C_2 (V2C_922_74),
	.V2C_3 (V2C_922_165),
	.V2C_4 (V2C_922_181),
	.V2C_5 (V2C_922_204),
	.V2C_6 (V2C_922_262),
	.V (V_922)
);

VNU_6 #(quan_width) VNU923 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_923),
	.C2V_2 (C2V_80_923),
	.C2V_3 (C2V_171_923),
	.C2V_4 (C2V_187_923),
	.C2V_5 (C2V_210_923),
	.C2V_6 (C2V_268_923),
	.L (L_923),
	.V2C_1 (V2C_923_35),
	.V2C_2 (V2C_923_80),
	.V2C_3 (V2C_923_171),
	.V2C_4 (V2C_923_187),
	.V2C_5 (V2C_923_210),
	.V2C_6 (V2C_923_268),
	.V (V_923)
);

VNU_6 #(quan_width) VNU924 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_924),
	.C2V_2 (C2V_86_924),
	.C2V_3 (C2V_177_924),
	.C2V_4 (C2V_193_924),
	.C2V_5 (C2V_216_924),
	.C2V_6 (C2V_274_924),
	.L (L_924),
	.V2C_1 (V2C_924_41),
	.V2C_2 (V2C_924_86),
	.V2C_3 (V2C_924_177),
	.V2C_4 (V2C_924_193),
	.V2C_5 (V2C_924_216),
	.V2C_6 (V2C_924_274),
	.V (V_924)
);

VNU_6 #(quan_width) VNU925 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_925),
	.C2V_2 (C2V_92_925),
	.C2V_3 (C2V_183_925),
	.C2V_4 (C2V_199_925),
	.C2V_5 (C2V_222_925),
	.C2V_6 (C2V_280_925),
	.L (L_925),
	.V2C_1 (V2C_925_47),
	.V2C_2 (V2C_925_92),
	.V2C_3 (V2C_925_183),
	.V2C_4 (V2C_925_199),
	.V2C_5 (V2C_925_222),
	.V2C_6 (V2C_925_280),
	.V (V_925)
);

VNU_6 #(quan_width) VNU926 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_926),
	.C2V_2 (C2V_98_926),
	.C2V_3 (C2V_189_926),
	.C2V_4 (C2V_205_926),
	.C2V_5 (C2V_228_926),
	.C2V_6 (C2V_286_926),
	.L (L_926),
	.V2C_1 (V2C_926_53),
	.V2C_2 (V2C_926_98),
	.V2C_3 (V2C_926_189),
	.V2C_4 (V2C_926_205),
	.V2C_5 (V2C_926_228),
	.V2C_6 (V2C_926_286),
	.V (V_926)
);

VNU_6 #(quan_width) VNU927 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_927),
	.C2V_2 (C2V_59_927),
	.C2V_3 (C2V_104_927),
	.C2V_4 (C2V_195_927),
	.C2V_5 (C2V_211_927),
	.C2V_6 (C2V_234_927),
	.L (L_927),
	.V2C_1 (V2C_927_4),
	.V2C_2 (V2C_927_59),
	.V2C_3 (V2C_927_104),
	.V2C_4 (V2C_927_195),
	.V2C_5 (V2C_927_211),
	.V2C_6 (V2C_927_234),
	.V (V_927)
);

VNU_6 #(quan_width) VNU928 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_928),
	.C2V_2 (C2V_65_928),
	.C2V_3 (C2V_110_928),
	.C2V_4 (C2V_201_928),
	.C2V_5 (C2V_217_928),
	.C2V_6 (C2V_240_928),
	.L (L_928),
	.V2C_1 (V2C_928_10),
	.V2C_2 (V2C_928_65),
	.V2C_3 (V2C_928_110),
	.V2C_4 (V2C_928_201),
	.V2C_5 (V2C_928_217),
	.V2C_6 (V2C_928_240),
	.V (V_928)
);

VNU_6 #(quan_width) VNU929 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_929),
	.C2V_2 (C2V_71_929),
	.C2V_3 (C2V_116_929),
	.C2V_4 (C2V_207_929),
	.C2V_5 (C2V_223_929),
	.C2V_6 (C2V_246_929),
	.L (L_929),
	.V2C_1 (V2C_929_16),
	.V2C_2 (V2C_929_71),
	.V2C_3 (V2C_929_116),
	.V2C_4 (V2C_929_207),
	.V2C_5 (V2C_929_223),
	.V2C_6 (V2C_929_246),
	.V (V_929)
);

VNU_6 #(quan_width) VNU930 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_930),
	.C2V_2 (C2V_77_930),
	.C2V_3 (C2V_122_930),
	.C2V_4 (C2V_213_930),
	.C2V_5 (C2V_229_930),
	.C2V_6 (C2V_252_930),
	.L (L_930),
	.V2C_1 (V2C_930_22),
	.V2C_2 (V2C_930_77),
	.V2C_3 (V2C_930_122),
	.V2C_4 (V2C_930_213),
	.V2C_5 (V2C_930_229),
	.V2C_6 (V2C_930_252),
	.V (V_930)
);

VNU_6 #(quan_width) VNU931 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_931),
	.C2V_2 (C2V_83_931),
	.C2V_3 (C2V_128_931),
	.C2V_4 (C2V_219_931),
	.C2V_5 (C2V_235_931),
	.C2V_6 (C2V_258_931),
	.L (L_931),
	.V2C_1 (V2C_931_28),
	.V2C_2 (V2C_931_83),
	.V2C_3 (V2C_931_128),
	.V2C_4 (V2C_931_219),
	.V2C_5 (V2C_931_235),
	.V2C_6 (V2C_931_258),
	.V (V_931)
);

VNU_6 #(quan_width) VNU932 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_932),
	.C2V_2 (C2V_89_932),
	.C2V_3 (C2V_134_932),
	.C2V_4 (C2V_225_932),
	.C2V_5 (C2V_241_932),
	.C2V_6 (C2V_264_932),
	.L (L_932),
	.V2C_1 (V2C_932_34),
	.V2C_2 (V2C_932_89),
	.V2C_3 (V2C_932_134),
	.V2C_4 (V2C_932_225),
	.V2C_5 (V2C_932_241),
	.V2C_6 (V2C_932_264),
	.V (V_932)
);

VNU_6 #(quan_width) VNU933 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_933),
	.C2V_2 (C2V_95_933),
	.C2V_3 (C2V_140_933),
	.C2V_4 (C2V_231_933),
	.C2V_5 (C2V_247_933),
	.C2V_6 (C2V_270_933),
	.L (L_933),
	.V2C_1 (V2C_933_40),
	.V2C_2 (V2C_933_95),
	.V2C_3 (V2C_933_140),
	.V2C_4 (V2C_933_231),
	.V2C_5 (V2C_933_247),
	.V2C_6 (V2C_933_270),
	.V (V_933)
);

VNU_6 #(quan_width) VNU934 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_934),
	.C2V_2 (C2V_101_934),
	.C2V_3 (C2V_146_934),
	.C2V_4 (C2V_237_934),
	.C2V_5 (C2V_253_934),
	.C2V_6 (C2V_276_934),
	.L (L_934),
	.V2C_1 (V2C_934_46),
	.V2C_2 (V2C_934_101),
	.V2C_3 (V2C_934_146),
	.V2C_4 (V2C_934_237),
	.V2C_5 (V2C_934_253),
	.V2C_6 (V2C_934_276),
	.V (V_934)
);

VNU_6 #(quan_width) VNU935 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_935),
	.C2V_2 (C2V_107_935),
	.C2V_3 (C2V_152_935),
	.C2V_4 (C2V_243_935),
	.C2V_5 (C2V_259_935),
	.C2V_6 (C2V_282_935),
	.L (L_935),
	.V2C_1 (V2C_935_52),
	.V2C_2 (V2C_935_107),
	.V2C_3 (V2C_935_152),
	.V2C_4 (V2C_935_243),
	.V2C_5 (V2C_935_259),
	.V2C_6 (V2C_935_282),
	.V (V_935)
);

VNU_6 #(quan_width) VNU936 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_936),
	.C2V_2 (C2V_113_936),
	.C2V_3 (C2V_158_936),
	.C2V_4 (C2V_249_936),
	.C2V_5 (C2V_265_936),
	.C2V_6 (C2V_288_936),
	.L (L_936),
	.V2C_1 (V2C_936_58),
	.V2C_2 (V2C_936_113),
	.V2C_3 (V2C_936_158),
	.V2C_4 (V2C_936_249),
	.V2C_5 (V2C_936_265),
	.V2C_6 (V2C_936_288),
	.V (V_936)
);

VNU_6 #(quan_width) VNU937 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_937),
	.C2V_2 (C2V_64_937),
	.C2V_3 (C2V_119_937),
	.C2V_4 (C2V_164_937),
	.C2V_5 (C2V_255_937),
	.C2V_6 (C2V_271_937),
	.L (L_937),
	.V2C_1 (V2C_937_6),
	.V2C_2 (V2C_937_64),
	.V2C_3 (V2C_937_119),
	.V2C_4 (V2C_937_164),
	.V2C_5 (V2C_937_255),
	.V2C_6 (V2C_937_271),
	.V (V_937)
);

VNU_6 #(quan_width) VNU938 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_938),
	.C2V_2 (C2V_70_938),
	.C2V_3 (C2V_125_938),
	.C2V_4 (C2V_170_938),
	.C2V_5 (C2V_261_938),
	.C2V_6 (C2V_277_938),
	.L (L_938),
	.V2C_1 (V2C_938_12),
	.V2C_2 (V2C_938_70),
	.V2C_3 (V2C_938_125),
	.V2C_4 (V2C_938_170),
	.V2C_5 (V2C_938_261),
	.V2C_6 (V2C_938_277),
	.V (V_938)
);

VNU_6 #(quan_width) VNU939 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_939),
	.C2V_2 (C2V_76_939),
	.C2V_3 (C2V_131_939),
	.C2V_4 (C2V_176_939),
	.C2V_5 (C2V_267_939),
	.C2V_6 (C2V_283_939),
	.L (L_939),
	.V2C_1 (V2C_939_18),
	.V2C_2 (V2C_939_76),
	.V2C_3 (V2C_939_131),
	.V2C_4 (V2C_939_176),
	.V2C_5 (V2C_939_267),
	.V2C_6 (V2C_939_283),
	.V (V_939)
);

VNU_6 #(quan_width) VNU940 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_940),
	.C2V_2 (C2V_24_940),
	.C2V_3 (C2V_82_940),
	.C2V_4 (C2V_137_940),
	.C2V_5 (C2V_182_940),
	.C2V_6 (C2V_273_940),
	.L (L_940),
	.V2C_1 (V2C_940_1),
	.V2C_2 (V2C_940_24),
	.V2C_3 (V2C_940_82),
	.V2C_4 (V2C_940_137),
	.V2C_5 (V2C_940_182),
	.V2C_6 (V2C_940_273),
	.V (V_940)
);

VNU_6 #(quan_width) VNU941 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_941),
	.C2V_2 (C2V_30_941),
	.C2V_3 (C2V_88_941),
	.C2V_4 (C2V_143_941),
	.C2V_5 (C2V_188_941),
	.C2V_6 (C2V_279_941),
	.L (L_941),
	.V2C_1 (V2C_941_7),
	.V2C_2 (V2C_941_30),
	.V2C_3 (V2C_941_88),
	.V2C_4 (V2C_941_143),
	.V2C_5 (V2C_941_188),
	.V2C_6 (V2C_941_279),
	.V (V_941)
);

VNU_6 #(quan_width) VNU942 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_942),
	.C2V_2 (C2V_36_942),
	.C2V_3 (C2V_94_942),
	.C2V_4 (C2V_149_942),
	.C2V_5 (C2V_194_942),
	.C2V_6 (C2V_285_942),
	.L (L_942),
	.V2C_1 (V2C_942_13),
	.V2C_2 (V2C_942_36),
	.V2C_3 (V2C_942_94),
	.V2C_4 (V2C_942_149),
	.V2C_5 (V2C_942_194),
	.V2C_6 (V2C_942_285),
	.V (V_942)
);

VNU_6 #(quan_width) VNU943 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_943),
	.C2V_2 (C2V_19_943),
	.C2V_3 (C2V_42_943),
	.C2V_4 (C2V_100_943),
	.C2V_5 (C2V_155_943),
	.C2V_6 (C2V_200_943),
	.L (L_943),
	.V2C_1 (V2C_943_3),
	.V2C_2 (V2C_943_19),
	.V2C_3 (V2C_943_42),
	.V2C_4 (V2C_943_100),
	.V2C_5 (V2C_943_155),
	.V2C_6 (V2C_943_200),
	.V (V_943)
);

VNU_6 #(quan_width) VNU944 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_944),
	.C2V_2 (C2V_25_944),
	.C2V_3 (C2V_48_944),
	.C2V_4 (C2V_106_944),
	.C2V_5 (C2V_161_944),
	.C2V_6 (C2V_206_944),
	.L (L_944),
	.V2C_1 (V2C_944_9),
	.V2C_2 (V2C_944_25),
	.V2C_3 (V2C_944_48),
	.V2C_4 (V2C_944_106),
	.V2C_5 (V2C_944_161),
	.V2C_6 (V2C_944_206),
	.V (V_944)
);

VNU_6 #(quan_width) VNU945 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_945),
	.C2V_2 (C2V_31_945),
	.C2V_3 (C2V_54_945),
	.C2V_4 (C2V_112_945),
	.C2V_5 (C2V_167_945),
	.C2V_6 (C2V_212_945),
	.L (L_945),
	.V2C_1 (V2C_945_15),
	.V2C_2 (V2C_945_31),
	.V2C_3 (V2C_945_54),
	.V2C_4 (V2C_945_112),
	.V2C_5 (V2C_945_167),
	.V2C_6 (V2C_945_212),
	.V (V_945)
);

VNU_6 #(quan_width) VNU946 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_946),
	.C2V_2 (C2V_37_946),
	.C2V_3 (C2V_60_946),
	.C2V_4 (C2V_118_946),
	.C2V_5 (C2V_173_946),
	.C2V_6 (C2V_218_946),
	.L (L_946),
	.V2C_1 (V2C_946_21),
	.V2C_2 (V2C_946_37),
	.V2C_3 (V2C_946_60),
	.V2C_4 (V2C_946_118),
	.V2C_5 (V2C_946_173),
	.V2C_6 (V2C_946_218),
	.V (V_946)
);

VNU_6 #(quan_width) VNU947 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_947),
	.C2V_2 (C2V_43_947),
	.C2V_3 (C2V_66_947),
	.C2V_4 (C2V_124_947),
	.C2V_5 (C2V_179_947),
	.C2V_6 (C2V_224_947),
	.L (L_947),
	.V2C_1 (V2C_947_27),
	.V2C_2 (V2C_947_43),
	.V2C_3 (V2C_947_66),
	.V2C_4 (V2C_947_124),
	.V2C_5 (V2C_947_179),
	.V2C_6 (V2C_947_224),
	.V (V_947)
);

VNU_6 #(quan_width) VNU948 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_948),
	.C2V_2 (C2V_49_948),
	.C2V_3 (C2V_72_948),
	.C2V_4 (C2V_130_948),
	.C2V_5 (C2V_185_948),
	.C2V_6 (C2V_230_948),
	.L (L_948),
	.V2C_1 (V2C_948_33),
	.V2C_2 (V2C_948_49),
	.V2C_3 (V2C_948_72),
	.V2C_4 (V2C_948_130),
	.V2C_5 (V2C_948_185),
	.V2C_6 (V2C_948_230),
	.V (V_948)
);

VNU_6 #(quan_width) VNU949 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_949),
	.C2V_2 (C2V_55_949),
	.C2V_3 (C2V_78_949),
	.C2V_4 (C2V_136_949),
	.C2V_5 (C2V_191_949),
	.C2V_6 (C2V_236_949),
	.L (L_949),
	.V2C_1 (V2C_949_39),
	.V2C_2 (V2C_949_55),
	.V2C_3 (V2C_949_78),
	.V2C_4 (V2C_949_136),
	.V2C_5 (V2C_949_191),
	.V2C_6 (V2C_949_236),
	.V (V_949)
);

VNU_6 #(quan_width) VNU950 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_950),
	.C2V_2 (C2V_61_950),
	.C2V_3 (C2V_84_950),
	.C2V_4 (C2V_142_950),
	.C2V_5 (C2V_197_950),
	.C2V_6 (C2V_242_950),
	.L (L_950),
	.V2C_1 (V2C_950_45),
	.V2C_2 (V2C_950_61),
	.V2C_3 (V2C_950_84),
	.V2C_4 (V2C_950_142),
	.V2C_5 (V2C_950_197),
	.V2C_6 (V2C_950_242),
	.V (V_950)
);

VNU_6 #(quan_width) VNU951 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_951),
	.C2V_2 (C2V_67_951),
	.C2V_3 (C2V_90_951),
	.C2V_4 (C2V_148_951),
	.C2V_5 (C2V_203_951),
	.C2V_6 (C2V_248_951),
	.L (L_951),
	.V2C_1 (V2C_951_51),
	.V2C_2 (V2C_951_67),
	.V2C_3 (V2C_951_90),
	.V2C_4 (V2C_951_148),
	.V2C_5 (V2C_951_203),
	.V2C_6 (V2C_951_248),
	.V (V_951)
);

VNU_6 #(quan_width) VNU952 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_952),
	.C2V_2 (C2V_73_952),
	.C2V_3 (C2V_96_952),
	.C2V_4 (C2V_154_952),
	.C2V_5 (C2V_209_952),
	.C2V_6 (C2V_254_952),
	.L (L_952),
	.V2C_1 (V2C_952_57),
	.V2C_2 (V2C_952_73),
	.V2C_3 (V2C_952_96),
	.V2C_4 (V2C_952_154),
	.V2C_5 (V2C_952_209),
	.V2C_6 (V2C_952_254),
	.V (V_952)
);

VNU_6 #(quan_width) VNU953 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_953),
	.C2V_2 (C2V_79_953),
	.C2V_3 (C2V_102_953),
	.C2V_4 (C2V_160_953),
	.C2V_5 (C2V_215_953),
	.C2V_6 (C2V_260_953),
	.L (L_953),
	.V2C_1 (V2C_953_63),
	.V2C_2 (V2C_953_79),
	.V2C_3 (V2C_953_102),
	.V2C_4 (V2C_953_160),
	.V2C_5 (V2C_953_215),
	.V2C_6 (V2C_953_260),
	.V (V_953)
);

VNU_6 #(quan_width) VNU954 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_954),
	.C2V_2 (C2V_85_954),
	.C2V_3 (C2V_108_954),
	.C2V_4 (C2V_166_954),
	.C2V_5 (C2V_221_954),
	.C2V_6 (C2V_266_954),
	.L (L_954),
	.V2C_1 (V2C_954_69),
	.V2C_2 (V2C_954_85),
	.V2C_3 (V2C_954_108),
	.V2C_4 (V2C_954_166),
	.V2C_5 (V2C_954_221),
	.V2C_6 (V2C_954_266),
	.V (V_954)
);

VNU_6 #(quan_width) VNU955 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_955),
	.C2V_2 (C2V_91_955),
	.C2V_3 (C2V_114_955),
	.C2V_4 (C2V_172_955),
	.C2V_5 (C2V_227_955),
	.C2V_6 (C2V_272_955),
	.L (L_955),
	.V2C_1 (V2C_955_75),
	.V2C_2 (V2C_955_91),
	.V2C_3 (V2C_955_114),
	.V2C_4 (V2C_955_172),
	.V2C_5 (V2C_955_227),
	.V2C_6 (V2C_955_272),
	.V (V_955)
);

VNU_6 #(quan_width) VNU956 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_956),
	.C2V_2 (C2V_97_956),
	.C2V_3 (C2V_120_956),
	.C2V_4 (C2V_178_956),
	.C2V_5 (C2V_233_956),
	.C2V_6 (C2V_278_956),
	.L (L_956),
	.V2C_1 (V2C_956_81),
	.V2C_2 (V2C_956_97),
	.V2C_3 (V2C_956_120),
	.V2C_4 (V2C_956_178),
	.V2C_5 (V2C_956_233),
	.V2C_6 (V2C_956_278),
	.V (V_956)
);

VNU_6 #(quan_width) VNU957 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_957),
	.C2V_2 (C2V_103_957),
	.C2V_3 (C2V_126_957),
	.C2V_4 (C2V_184_957),
	.C2V_5 (C2V_239_957),
	.C2V_6 (C2V_284_957),
	.L (L_957),
	.V2C_1 (V2C_957_87),
	.V2C_2 (V2C_957_103),
	.V2C_3 (V2C_957_126),
	.V2C_4 (V2C_957_184),
	.V2C_5 (V2C_957_239),
	.V2C_6 (V2C_957_284),
	.V (V_957)
);

VNU_6 #(quan_width) VNU958 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_958),
	.C2V_2 (C2V_93_958),
	.C2V_3 (C2V_109_958),
	.C2V_4 (C2V_132_958),
	.C2V_5 (C2V_190_958),
	.C2V_6 (C2V_245_958),
	.L (L_958),
	.V2C_1 (V2C_958_2),
	.V2C_2 (V2C_958_93),
	.V2C_3 (V2C_958_109),
	.V2C_4 (V2C_958_132),
	.V2C_5 (V2C_958_190),
	.V2C_6 (V2C_958_245),
	.V (V_958)
);

VNU_6 #(quan_width) VNU959 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_959),
	.C2V_2 (C2V_99_959),
	.C2V_3 (C2V_115_959),
	.C2V_4 (C2V_138_959),
	.C2V_5 (C2V_196_959),
	.C2V_6 (C2V_251_959),
	.L (L_959),
	.V2C_1 (V2C_959_8),
	.V2C_2 (V2C_959_99),
	.V2C_3 (V2C_959_115),
	.V2C_4 (V2C_959_138),
	.V2C_5 (V2C_959_196),
	.V2C_6 (V2C_959_251),
	.V (V_959)
);

VNU_6 #(quan_width) VNU960 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_960),
	.C2V_2 (C2V_105_960),
	.C2V_3 (C2V_121_960),
	.C2V_4 (C2V_144_960),
	.C2V_5 (C2V_202_960),
	.C2V_6 (C2V_257_960),
	.L (L_960),
	.V2C_1 (V2C_960_14),
	.V2C_2 (V2C_960_105),
	.V2C_3 (V2C_960_121),
	.V2C_4 (V2C_960_144),
	.V2C_5 (V2C_960_202),
	.V2C_6 (V2C_960_257),
	.V (V_960)
);

VNU_6 #(quan_width) VNU961 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_961),
	.C2V_2 (C2V_122_961),
	.C2V_3 (C2V_211_961),
	.C2V_4 (C2V_228_961),
	.C2V_5 (C2V_249_961),
	.C2V_6 (C2V_280_961),
	.L (L_961),
	.V2C_1 (V2C_961_5),
	.V2C_2 (V2C_961_122),
	.V2C_3 (V2C_961_211),
	.V2C_4 (V2C_961_228),
	.V2C_5 (V2C_961_249),
	.V2C_6 (V2C_961_280),
	.V (V_961)
);

VNU_6 #(quan_width) VNU962 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_962),
	.C2V_2 (C2V_128_962),
	.C2V_3 (C2V_217_962),
	.C2V_4 (C2V_234_962),
	.C2V_5 (C2V_255_962),
	.C2V_6 (C2V_286_962),
	.L (L_962),
	.V2C_1 (V2C_962_11),
	.V2C_2 (V2C_962_128),
	.V2C_3 (V2C_962_217),
	.V2C_4 (V2C_962_234),
	.V2C_5 (V2C_962_255),
	.V2C_6 (V2C_962_286),
	.V (V_962)
);

VNU_6 #(quan_width) VNU963 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_963),
	.C2V_2 (C2V_17_963),
	.C2V_3 (C2V_134_963),
	.C2V_4 (C2V_223_963),
	.C2V_5 (C2V_240_963),
	.C2V_6 (C2V_261_963),
	.L (L_963),
	.V2C_1 (V2C_963_4),
	.V2C_2 (V2C_963_17),
	.V2C_3 (V2C_963_134),
	.V2C_4 (V2C_963_223),
	.V2C_5 (V2C_963_240),
	.V2C_6 (V2C_963_261),
	.V (V_963)
);

VNU_6 #(quan_width) VNU964 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_964),
	.C2V_2 (C2V_23_964),
	.C2V_3 (C2V_140_964),
	.C2V_4 (C2V_229_964),
	.C2V_5 (C2V_246_964),
	.C2V_6 (C2V_267_964),
	.L (L_964),
	.V2C_1 (V2C_964_10),
	.V2C_2 (V2C_964_23),
	.V2C_3 (V2C_964_140),
	.V2C_4 (V2C_964_229),
	.V2C_5 (V2C_964_246),
	.V2C_6 (V2C_964_267),
	.V (V_964)
);

VNU_6 #(quan_width) VNU965 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_965),
	.C2V_2 (C2V_29_965),
	.C2V_3 (C2V_146_965),
	.C2V_4 (C2V_235_965),
	.C2V_5 (C2V_252_965),
	.C2V_6 (C2V_273_965),
	.L (L_965),
	.V2C_1 (V2C_965_16),
	.V2C_2 (V2C_965_29),
	.V2C_3 (V2C_965_146),
	.V2C_4 (V2C_965_235),
	.V2C_5 (V2C_965_252),
	.V2C_6 (V2C_965_273),
	.V (V_965)
);

VNU_6 #(quan_width) VNU966 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_966),
	.C2V_2 (C2V_35_966),
	.C2V_3 (C2V_152_966),
	.C2V_4 (C2V_241_966),
	.C2V_5 (C2V_258_966),
	.C2V_6 (C2V_279_966),
	.L (L_966),
	.V2C_1 (V2C_966_22),
	.V2C_2 (V2C_966_35),
	.V2C_3 (V2C_966_152),
	.V2C_4 (V2C_966_241),
	.V2C_5 (V2C_966_258),
	.V2C_6 (V2C_966_279),
	.V (V_966)
);

VNU_6 #(quan_width) VNU967 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_967),
	.C2V_2 (C2V_41_967),
	.C2V_3 (C2V_158_967),
	.C2V_4 (C2V_247_967),
	.C2V_5 (C2V_264_967),
	.C2V_6 (C2V_285_967),
	.L (L_967),
	.V2C_1 (V2C_967_28),
	.V2C_2 (V2C_967_41),
	.V2C_3 (V2C_967_158),
	.V2C_4 (V2C_967_247),
	.V2C_5 (V2C_967_264),
	.V2C_6 (V2C_967_285),
	.V (V_967)
);

VNU_6 #(quan_width) VNU968 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_968),
	.C2V_2 (C2V_34_968),
	.C2V_3 (C2V_47_968),
	.C2V_4 (C2V_164_968),
	.C2V_5 (C2V_253_968),
	.C2V_6 (C2V_270_968),
	.L (L_968),
	.V2C_1 (V2C_968_3),
	.V2C_2 (V2C_968_34),
	.V2C_3 (V2C_968_47),
	.V2C_4 (V2C_968_164),
	.V2C_5 (V2C_968_253),
	.V2C_6 (V2C_968_270),
	.V (V_968)
);

VNU_6 #(quan_width) VNU969 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_969),
	.C2V_2 (C2V_40_969),
	.C2V_3 (C2V_53_969),
	.C2V_4 (C2V_170_969),
	.C2V_5 (C2V_259_969),
	.C2V_6 (C2V_276_969),
	.L (L_969),
	.V2C_1 (V2C_969_9),
	.V2C_2 (V2C_969_40),
	.V2C_3 (V2C_969_53),
	.V2C_4 (V2C_969_170),
	.V2C_5 (V2C_969_259),
	.V2C_6 (V2C_969_276),
	.V (V_969)
);

VNU_6 #(quan_width) VNU970 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_970),
	.C2V_2 (C2V_46_970),
	.C2V_3 (C2V_59_970),
	.C2V_4 (C2V_176_970),
	.C2V_5 (C2V_265_970),
	.C2V_6 (C2V_282_970),
	.L (L_970),
	.V2C_1 (V2C_970_15),
	.V2C_2 (V2C_970_46),
	.V2C_3 (V2C_970_59),
	.V2C_4 (V2C_970_176),
	.V2C_5 (V2C_970_265),
	.V2C_6 (V2C_970_282),
	.V (V_970)
);

VNU_6 #(quan_width) VNU971 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_971),
	.C2V_2 (C2V_52_971),
	.C2V_3 (C2V_65_971),
	.C2V_4 (C2V_182_971),
	.C2V_5 (C2V_271_971),
	.C2V_6 (C2V_288_971),
	.L (L_971),
	.V2C_1 (V2C_971_21),
	.V2C_2 (V2C_971_52),
	.V2C_3 (V2C_971_65),
	.V2C_4 (V2C_971_182),
	.V2C_5 (V2C_971_271),
	.V2C_6 (V2C_971_288),
	.V (V_971)
);

VNU_6 #(quan_width) VNU972 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_972),
	.C2V_2 (C2V_27_972),
	.C2V_3 (C2V_58_972),
	.C2V_4 (C2V_71_972),
	.C2V_5 (C2V_188_972),
	.C2V_6 (C2V_277_972),
	.L (L_972),
	.V2C_1 (V2C_972_6),
	.V2C_2 (V2C_972_27),
	.V2C_3 (V2C_972_58),
	.V2C_4 (V2C_972_71),
	.V2C_5 (V2C_972_188),
	.V2C_6 (V2C_972_277),
	.V (V_972)
);

VNU_6 #(quan_width) VNU973 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_973),
	.C2V_2 (C2V_33_973),
	.C2V_3 (C2V_64_973),
	.C2V_4 (C2V_77_973),
	.C2V_5 (C2V_194_973),
	.C2V_6 (C2V_283_973),
	.L (L_973),
	.V2C_1 (V2C_973_12),
	.V2C_2 (V2C_973_33),
	.V2C_3 (V2C_973_64),
	.V2C_4 (V2C_973_77),
	.V2C_5 (V2C_973_194),
	.V2C_6 (V2C_973_283),
	.V (V_973)
);

VNU_6 #(quan_width) VNU974 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_974),
	.C2V_2 (C2V_18_974),
	.C2V_3 (C2V_39_974),
	.C2V_4 (C2V_70_974),
	.C2V_5 (C2V_83_974),
	.C2V_6 (C2V_200_974),
	.L (L_974),
	.V2C_1 (V2C_974_1),
	.V2C_2 (V2C_974_18),
	.V2C_3 (V2C_974_39),
	.V2C_4 (V2C_974_70),
	.V2C_5 (V2C_974_83),
	.V2C_6 (V2C_974_200),
	.V (V_974)
);

VNU_6 #(quan_width) VNU975 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_975),
	.C2V_2 (C2V_24_975),
	.C2V_3 (C2V_45_975),
	.C2V_4 (C2V_76_975),
	.C2V_5 (C2V_89_975),
	.C2V_6 (C2V_206_975),
	.L (L_975),
	.V2C_1 (V2C_975_7),
	.V2C_2 (V2C_975_24),
	.V2C_3 (V2C_975_45),
	.V2C_4 (V2C_975_76),
	.V2C_5 (V2C_975_89),
	.V2C_6 (V2C_975_206),
	.V (V_975)
);

VNU_6 #(quan_width) VNU976 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_976),
	.C2V_2 (C2V_30_976),
	.C2V_3 (C2V_51_976),
	.C2V_4 (C2V_82_976),
	.C2V_5 (C2V_95_976),
	.C2V_6 (C2V_212_976),
	.L (L_976),
	.V2C_1 (V2C_976_13),
	.V2C_2 (V2C_976_30),
	.V2C_3 (V2C_976_51),
	.V2C_4 (V2C_976_82),
	.V2C_5 (V2C_976_95),
	.V2C_6 (V2C_976_212),
	.V (V_976)
);

VNU_6 #(quan_width) VNU977 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_977),
	.C2V_2 (C2V_36_977),
	.C2V_3 (C2V_57_977),
	.C2V_4 (C2V_88_977),
	.C2V_5 (C2V_101_977),
	.C2V_6 (C2V_218_977),
	.L (L_977),
	.V2C_1 (V2C_977_19),
	.V2C_2 (V2C_977_36),
	.V2C_3 (V2C_977_57),
	.V2C_4 (V2C_977_88),
	.V2C_5 (V2C_977_101),
	.V2C_6 (V2C_977_218),
	.V (V_977)
);

VNU_6 #(quan_width) VNU978 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_978),
	.C2V_2 (C2V_42_978),
	.C2V_3 (C2V_63_978),
	.C2V_4 (C2V_94_978),
	.C2V_5 (C2V_107_978),
	.C2V_6 (C2V_224_978),
	.L (L_978),
	.V2C_1 (V2C_978_25),
	.V2C_2 (V2C_978_42),
	.V2C_3 (V2C_978_63),
	.V2C_4 (V2C_978_94),
	.V2C_5 (V2C_978_107),
	.V2C_6 (V2C_978_224),
	.V (V_978)
);

VNU_6 #(quan_width) VNU979 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_979),
	.C2V_2 (C2V_48_979),
	.C2V_3 (C2V_69_979),
	.C2V_4 (C2V_100_979),
	.C2V_5 (C2V_113_979),
	.C2V_6 (C2V_230_979),
	.L (L_979),
	.V2C_1 (V2C_979_31),
	.V2C_2 (V2C_979_48),
	.V2C_3 (V2C_979_69),
	.V2C_4 (V2C_979_100),
	.V2C_5 (V2C_979_113),
	.V2C_6 (V2C_979_230),
	.V (V_979)
);

VNU_6 #(quan_width) VNU980 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_980),
	.C2V_2 (C2V_54_980),
	.C2V_3 (C2V_75_980),
	.C2V_4 (C2V_106_980),
	.C2V_5 (C2V_119_980),
	.C2V_6 (C2V_236_980),
	.L (L_980),
	.V2C_1 (V2C_980_37),
	.V2C_2 (V2C_980_54),
	.V2C_3 (V2C_980_75),
	.V2C_4 (V2C_980_106),
	.V2C_5 (V2C_980_119),
	.V2C_6 (V2C_980_236),
	.V (V_980)
);

VNU_6 #(quan_width) VNU981 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_981),
	.C2V_2 (C2V_60_981),
	.C2V_3 (C2V_81_981),
	.C2V_4 (C2V_112_981),
	.C2V_5 (C2V_125_981),
	.C2V_6 (C2V_242_981),
	.L (L_981),
	.V2C_1 (V2C_981_43),
	.V2C_2 (V2C_981_60),
	.V2C_3 (V2C_981_81),
	.V2C_4 (V2C_981_112),
	.V2C_5 (V2C_981_125),
	.V2C_6 (V2C_981_242),
	.V (V_981)
);

VNU_6 #(quan_width) VNU982 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_982),
	.C2V_2 (C2V_66_982),
	.C2V_3 (C2V_87_982),
	.C2V_4 (C2V_118_982),
	.C2V_5 (C2V_131_982),
	.C2V_6 (C2V_248_982),
	.L (L_982),
	.V2C_1 (V2C_982_49),
	.V2C_2 (V2C_982_66),
	.V2C_3 (V2C_982_87),
	.V2C_4 (V2C_982_118),
	.V2C_5 (V2C_982_131),
	.V2C_6 (V2C_982_248),
	.V (V_982)
);

VNU_6 #(quan_width) VNU983 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_983),
	.C2V_2 (C2V_72_983),
	.C2V_3 (C2V_93_983),
	.C2V_4 (C2V_124_983),
	.C2V_5 (C2V_137_983),
	.C2V_6 (C2V_254_983),
	.L (L_983),
	.V2C_1 (V2C_983_55),
	.V2C_2 (V2C_983_72),
	.V2C_3 (V2C_983_93),
	.V2C_4 (V2C_983_124),
	.V2C_5 (V2C_983_137),
	.V2C_6 (V2C_983_254),
	.V (V_983)
);

VNU_6 #(quan_width) VNU984 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_984),
	.C2V_2 (C2V_78_984),
	.C2V_3 (C2V_99_984),
	.C2V_4 (C2V_130_984),
	.C2V_5 (C2V_143_984),
	.C2V_6 (C2V_260_984),
	.L (L_984),
	.V2C_1 (V2C_984_61),
	.V2C_2 (V2C_984_78),
	.V2C_3 (V2C_984_99),
	.V2C_4 (V2C_984_130),
	.V2C_5 (V2C_984_143),
	.V2C_6 (V2C_984_260),
	.V (V_984)
);

VNU_6 #(quan_width) VNU985 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_985),
	.C2V_2 (C2V_84_985),
	.C2V_3 (C2V_105_985),
	.C2V_4 (C2V_136_985),
	.C2V_5 (C2V_149_985),
	.C2V_6 (C2V_266_985),
	.L (L_985),
	.V2C_1 (V2C_985_67),
	.V2C_2 (V2C_985_84),
	.V2C_3 (V2C_985_105),
	.V2C_4 (V2C_985_136),
	.V2C_5 (V2C_985_149),
	.V2C_6 (V2C_985_266),
	.V (V_985)
);

VNU_6 #(quan_width) VNU986 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_986),
	.C2V_2 (C2V_90_986),
	.C2V_3 (C2V_111_986),
	.C2V_4 (C2V_142_986),
	.C2V_5 (C2V_155_986),
	.C2V_6 (C2V_272_986),
	.L (L_986),
	.V2C_1 (V2C_986_73),
	.V2C_2 (V2C_986_90),
	.V2C_3 (V2C_986_111),
	.V2C_4 (V2C_986_142),
	.V2C_5 (V2C_986_155),
	.V2C_6 (V2C_986_272),
	.V (V_986)
);

VNU_6 #(quan_width) VNU987 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_987),
	.C2V_2 (C2V_96_987),
	.C2V_3 (C2V_117_987),
	.C2V_4 (C2V_148_987),
	.C2V_5 (C2V_161_987),
	.C2V_6 (C2V_278_987),
	.L (L_987),
	.V2C_1 (V2C_987_79),
	.V2C_2 (V2C_987_96),
	.V2C_3 (V2C_987_117),
	.V2C_4 (V2C_987_148),
	.V2C_5 (V2C_987_161),
	.V2C_6 (V2C_987_278),
	.V (V_987)
);

VNU_6 #(quan_width) VNU988 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_988),
	.C2V_2 (C2V_102_988),
	.C2V_3 (C2V_123_988),
	.C2V_4 (C2V_154_988),
	.C2V_5 (C2V_167_988),
	.C2V_6 (C2V_284_988),
	.L (L_988),
	.V2C_1 (V2C_988_85),
	.V2C_2 (V2C_988_102),
	.V2C_3 (V2C_988_123),
	.V2C_4 (V2C_988_154),
	.V2C_5 (V2C_988_167),
	.V2C_6 (V2C_988_284),
	.V (V_988)
);

VNU_6 #(quan_width) VNU989 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_989),
	.C2V_2 (C2V_91_989),
	.C2V_3 (C2V_108_989),
	.C2V_4 (C2V_129_989),
	.C2V_5 (C2V_160_989),
	.C2V_6 (C2V_173_989),
	.L (L_989),
	.V2C_1 (V2C_989_2),
	.V2C_2 (V2C_989_91),
	.V2C_3 (V2C_989_108),
	.V2C_4 (V2C_989_129),
	.V2C_5 (V2C_989_160),
	.V2C_6 (V2C_989_173),
	.V (V_989)
);

VNU_6 #(quan_width) VNU990 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_990),
	.C2V_2 (C2V_97_990),
	.C2V_3 (C2V_114_990),
	.C2V_4 (C2V_135_990),
	.C2V_5 (C2V_166_990),
	.C2V_6 (C2V_179_990),
	.L (L_990),
	.V2C_1 (V2C_990_8),
	.V2C_2 (V2C_990_97),
	.V2C_3 (V2C_990_114),
	.V2C_4 (V2C_990_135),
	.V2C_5 (V2C_990_166),
	.V2C_6 (V2C_990_179),
	.V (V_990)
);

VNU_6 #(quan_width) VNU991 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_991),
	.C2V_2 (C2V_103_991),
	.C2V_3 (C2V_120_991),
	.C2V_4 (C2V_141_991),
	.C2V_5 (C2V_172_991),
	.C2V_6 (C2V_185_991),
	.L (L_991),
	.V2C_1 (V2C_991_14),
	.V2C_2 (V2C_991_103),
	.V2C_3 (V2C_991_120),
	.V2C_4 (V2C_991_141),
	.V2C_5 (V2C_991_172),
	.V2C_6 (V2C_991_185),
	.V (V_991)
);

VNU_6 #(quan_width) VNU992 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_992),
	.C2V_2 (C2V_109_992),
	.C2V_3 (C2V_126_992),
	.C2V_4 (C2V_147_992),
	.C2V_5 (C2V_178_992),
	.C2V_6 (C2V_191_992),
	.L (L_992),
	.V2C_1 (V2C_992_20),
	.V2C_2 (V2C_992_109),
	.V2C_3 (V2C_992_126),
	.V2C_4 (V2C_992_147),
	.V2C_5 (V2C_992_178),
	.V2C_6 (V2C_992_191),
	.V (V_992)
);

VNU_6 #(quan_width) VNU993 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_993),
	.C2V_2 (C2V_115_993),
	.C2V_3 (C2V_132_993),
	.C2V_4 (C2V_153_993),
	.C2V_5 (C2V_184_993),
	.C2V_6 (C2V_197_993),
	.L (L_993),
	.V2C_1 (V2C_993_26),
	.V2C_2 (V2C_993_115),
	.V2C_3 (V2C_993_132),
	.V2C_4 (V2C_993_153),
	.V2C_5 (V2C_993_184),
	.V2C_6 (V2C_993_197),
	.V (V_993)
);

VNU_6 #(quan_width) VNU994 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_994),
	.C2V_2 (C2V_121_994),
	.C2V_3 (C2V_138_994),
	.C2V_4 (C2V_159_994),
	.C2V_5 (C2V_190_994),
	.C2V_6 (C2V_203_994),
	.L (L_994),
	.V2C_1 (V2C_994_32),
	.V2C_2 (V2C_994_121),
	.V2C_3 (V2C_994_138),
	.V2C_4 (V2C_994_159),
	.V2C_5 (V2C_994_190),
	.V2C_6 (V2C_994_203),
	.V (V_994)
);

VNU_6 #(quan_width) VNU995 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_995),
	.C2V_2 (C2V_127_995),
	.C2V_3 (C2V_144_995),
	.C2V_4 (C2V_165_995),
	.C2V_5 (C2V_196_995),
	.C2V_6 (C2V_209_995),
	.L (L_995),
	.V2C_1 (V2C_995_38),
	.V2C_2 (V2C_995_127),
	.V2C_3 (V2C_995_144),
	.V2C_4 (V2C_995_165),
	.V2C_5 (V2C_995_196),
	.V2C_6 (V2C_995_209),
	.V (V_995)
);

VNU_6 #(quan_width) VNU996 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_996),
	.C2V_2 (C2V_133_996),
	.C2V_3 (C2V_150_996),
	.C2V_4 (C2V_171_996),
	.C2V_5 (C2V_202_996),
	.C2V_6 (C2V_215_996),
	.L (L_996),
	.V2C_1 (V2C_996_44),
	.V2C_2 (V2C_996_133),
	.V2C_3 (V2C_996_150),
	.V2C_4 (V2C_996_171),
	.V2C_5 (V2C_996_202),
	.V2C_6 (V2C_996_215),
	.V (V_996)
);

VNU_6 #(quan_width) VNU997 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_997),
	.C2V_2 (C2V_139_997),
	.C2V_3 (C2V_156_997),
	.C2V_4 (C2V_177_997),
	.C2V_5 (C2V_208_997),
	.C2V_6 (C2V_221_997),
	.L (L_997),
	.V2C_1 (V2C_997_50),
	.V2C_2 (V2C_997_139),
	.V2C_3 (V2C_997_156),
	.V2C_4 (V2C_997_177),
	.V2C_5 (V2C_997_208),
	.V2C_6 (V2C_997_221),
	.V (V_997)
);

VNU_6 #(quan_width) VNU998 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_998),
	.C2V_2 (C2V_145_998),
	.C2V_3 (C2V_162_998),
	.C2V_4 (C2V_183_998),
	.C2V_5 (C2V_214_998),
	.C2V_6 (C2V_227_998),
	.L (L_998),
	.V2C_1 (V2C_998_56),
	.V2C_2 (V2C_998_145),
	.V2C_3 (V2C_998_162),
	.V2C_4 (V2C_998_183),
	.V2C_5 (V2C_998_214),
	.V2C_6 (V2C_998_227),
	.V (V_998)
);

VNU_6 #(quan_width) VNU999 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_999),
	.C2V_2 (C2V_151_999),
	.C2V_3 (C2V_168_999),
	.C2V_4 (C2V_189_999),
	.C2V_5 (C2V_220_999),
	.C2V_6 (C2V_233_999),
	.L (L_999),
	.V2C_1 (V2C_999_62),
	.V2C_2 (V2C_999_151),
	.V2C_3 (V2C_999_168),
	.V2C_4 (V2C_999_189),
	.V2C_5 (V2C_999_220),
	.V2C_6 (V2C_999_233),
	.V (V_999)
);

VNU_6 #(quan_width) VNU1000 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_1000),
	.C2V_2 (C2V_157_1000),
	.C2V_3 (C2V_174_1000),
	.C2V_4 (C2V_195_1000),
	.C2V_5 (C2V_226_1000),
	.C2V_6 (C2V_239_1000),
	.L (L_1000),
	.V2C_1 (V2C_1000_68),
	.V2C_2 (V2C_1000_157),
	.V2C_3 (V2C_1000_174),
	.V2C_4 (V2C_1000_195),
	.V2C_5 (V2C_1000_226),
	.V2C_6 (V2C_1000_239),
	.V (V_1000)
);

VNU_6 #(quan_width) VNU1001 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_1001),
	.C2V_2 (C2V_163_1001),
	.C2V_3 (C2V_180_1001),
	.C2V_4 (C2V_201_1001),
	.C2V_5 (C2V_232_1001),
	.C2V_6 (C2V_245_1001),
	.L (L_1001),
	.V2C_1 (V2C_1001_74),
	.V2C_2 (V2C_1001_163),
	.V2C_3 (V2C_1001_180),
	.V2C_4 (V2C_1001_201),
	.V2C_5 (V2C_1001_232),
	.V2C_6 (V2C_1001_245),
	.V (V_1001)
);

VNU_6 #(quan_width) VNU1002 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_80_1002),
	.C2V_2 (C2V_169_1002),
	.C2V_3 (C2V_186_1002),
	.C2V_4 (C2V_207_1002),
	.C2V_5 (C2V_238_1002),
	.C2V_6 (C2V_251_1002),
	.L (L_1002),
	.V2C_1 (V2C_1002_80),
	.V2C_2 (V2C_1002_169),
	.V2C_3 (V2C_1002_186),
	.V2C_4 (V2C_1002_207),
	.V2C_5 (V2C_1002_238),
	.V2C_6 (V2C_1002_251),
	.V (V_1002)
);

VNU_6 #(quan_width) VNU1003 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_86_1003),
	.C2V_2 (C2V_175_1003),
	.C2V_3 (C2V_192_1003),
	.C2V_4 (C2V_213_1003),
	.C2V_5 (C2V_244_1003),
	.C2V_6 (C2V_257_1003),
	.L (L_1003),
	.V2C_1 (V2C_1003_86),
	.V2C_2 (V2C_1003_175),
	.V2C_3 (V2C_1003_192),
	.V2C_4 (V2C_1003_213),
	.V2C_5 (V2C_1003_244),
	.V2C_6 (V2C_1003_257),
	.V (V_1003)
);

VNU_6 #(quan_width) VNU1004 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_92_1004),
	.C2V_2 (C2V_181_1004),
	.C2V_3 (C2V_198_1004),
	.C2V_4 (C2V_219_1004),
	.C2V_5 (C2V_250_1004),
	.C2V_6 (C2V_263_1004),
	.L (L_1004),
	.V2C_1 (V2C_1004_92),
	.V2C_2 (V2C_1004_181),
	.V2C_3 (V2C_1004_198),
	.V2C_4 (V2C_1004_219),
	.V2C_5 (V2C_1004_250),
	.V2C_6 (V2C_1004_263),
	.V (V_1004)
);

VNU_6 #(quan_width) VNU1005 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_98_1005),
	.C2V_2 (C2V_187_1005),
	.C2V_3 (C2V_204_1005),
	.C2V_4 (C2V_225_1005),
	.C2V_5 (C2V_256_1005),
	.C2V_6 (C2V_269_1005),
	.L (L_1005),
	.V2C_1 (V2C_1005_98),
	.V2C_2 (V2C_1005_187),
	.V2C_3 (V2C_1005_204),
	.V2C_4 (V2C_1005_225),
	.V2C_5 (V2C_1005_256),
	.V2C_6 (V2C_1005_269),
	.V (V_1005)
);

VNU_6 #(quan_width) VNU1006 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_104_1006),
	.C2V_2 (C2V_193_1006),
	.C2V_3 (C2V_210_1006),
	.C2V_4 (C2V_231_1006),
	.C2V_5 (C2V_262_1006),
	.C2V_6 (C2V_275_1006),
	.L (L_1006),
	.V2C_1 (V2C_1006_104),
	.V2C_2 (V2C_1006_193),
	.V2C_3 (V2C_1006_210),
	.V2C_4 (V2C_1006_231),
	.V2C_5 (V2C_1006_262),
	.V2C_6 (V2C_1006_275),
	.V (V_1006)
);

VNU_6 #(quan_width) VNU1007 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_110_1007),
	.C2V_2 (C2V_199_1007),
	.C2V_3 (C2V_216_1007),
	.C2V_4 (C2V_237_1007),
	.C2V_5 (C2V_268_1007),
	.C2V_6 (C2V_281_1007),
	.L (L_1007),
	.V2C_1 (V2C_1007_110),
	.V2C_2 (V2C_1007_199),
	.V2C_3 (V2C_1007_216),
	.V2C_4 (V2C_1007_237),
	.V2C_5 (V2C_1007_268),
	.V2C_6 (V2C_1007_281),
	.V (V_1007)
);

VNU_6 #(quan_width) VNU1008 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_116_1008),
	.C2V_2 (C2V_205_1008),
	.C2V_3 (C2V_222_1008),
	.C2V_4 (C2V_243_1008),
	.C2V_5 (C2V_274_1008),
	.C2V_6 (C2V_287_1008),
	.L (L_1008),
	.V2C_1 (V2C_1008_116),
	.V2C_2 (V2C_1008_205),
	.V2C_3 (V2C_1008_222),
	.V2C_4 (V2C_1008_243),
	.V2C_5 (V2C_1008_274),
	.V2C_6 (V2C_1008_287),
	.V (V_1008)
);

VNU_6 #(quan_width) VNU1009 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_1009),
	.C2V_2 (C2V_114_1009),
	.C2V_3 (C2V_177_1009),
	.C2V_4 (C2V_218_1009),
	.C2V_5 (C2V_265_1009),
	.C2V_6 (C2V_269_1009),
	.L (L_1009),
	.V2C_1 (V2C_1009_100),
	.V2C_2 (V2C_1009_114),
	.V2C_3 (V2C_1009_177),
	.V2C_4 (V2C_1009_218),
	.V2C_5 (V2C_1009_265),
	.V2C_6 (V2C_1009_269),
	.V (V_1009)
);

VNU_6 #(quan_width) VNU1010 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_1010),
	.C2V_2 (C2V_120_1010),
	.C2V_3 (C2V_183_1010),
	.C2V_4 (C2V_224_1010),
	.C2V_5 (C2V_271_1010),
	.C2V_6 (C2V_275_1010),
	.L (L_1010),
	.V2C_1 (V2C_1010_106),
	.V2C_2 (V2C_1010_120),
	.V2C_3 (V2C_1010_183),
	.V2C_4 (V2C_1010_224),
	.V2C_5 (V2C_1010_271),
	.V2C_6 (V2C_1010_275),
	.V (V_1010)
);

VNU_6 #(quan_width) VNU1011 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_1011),
	.C2V_2 (C2V_126_1011),
	.C2V_3 (C2V_189_1011),
	.C2V_4 (C2V_230_1011),
	.C2V_5 (C2V_277_1011),
	.C2V_6 (C2V_281_1011),
	.L (L_1011),
	.V2C_1 (V2C_1011_112),
	.V2C_2 (V2C_1011_126),
	.V2C_3 (V2C_1011_189),
	.V2C_4 (V2C_1011_230),
	.V2C_5 (V2C_1011_277),
	.V2C_6 (V2C_1011_281),
	.V (V_1011)
);

VNU_6 #(quan_width) VNU1012 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_118_1012),
	.C2V_2 (C2V_132_1012),
	.C2V_3 (C2V_195_1012),
	.C2V_4 (C2V_236_1012),
	.C2V_5 (C2V_283_1012),
	.C2V_6 (C2V_287_1012),
	.L (L_1012),
	.V2C_1 (V2C_1012_118),
	.V2C_2 (V2C_1012_132),
	.V2C_3 (V2C_1012_195),
	.V2C_4 (V2C_1012_236),
	.V2C_5 (V2C_1012_283),
	.V2C_6 (V2C_1012_287),
	.V (V_1012)
);

VNU_6 #(quan_width) VNU1013 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_1013),
	.C2V_2 (C2V_5_1013),
	.C2V_3 (C2V_124_1013),
	.C2V_4 (C2V_138_1013),
	.C2V_5 (C2V_201_1013),
	.C2V_6 (C2V_242_1013),
	.L (L_1013),
	.V2C_1 (V2C_1013_1),
	.V2C_2 (V2C_1013_5),
	.V2C_3 (V2C_1013_124),
	.V2C_4 (V2C_1013_138),
	.V2C_5 (V2C_1013_201),
	.V2C_6 (V2C_1013_242),
	.V (V_1013)
);

VNU_6 #(quan_width) VNU1014 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_1014),
	.C2V_2 (C2V_11_1014),
	.C2V_3 (C2V_130_1014),
	.C2V_4 (C2V_144_1014),
	.C2V_5 (C2V_207_1014),
	.C2V_6 (C2V_248_1014),
	.L (L_1014),
	.V2C_1 (V2C_1014_7),
	.V2C_2 (V2C_1014_11),
	.V2C_3 (V2C_1014_130),
	.V2C_4 (V2C_1014_144),
	.V2C_5 (V2C_1014_207),
	.V2C_6 (V2C_1014_248),
	.V (V_1014)
);

VNU_6 #(quan_width) VNU1015 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_1015),
	.C2V_2 (C2V_17_1015),
	.C2V_3 (C2V_136_1015),
	.C2V_4 (C2V_150_1015),
	.C2V_5 (C2V_213_1015),
	.C2V_6 (C2V_254_1015),
	.L (L_1015),
	.V2C_1 (V2C_1015_13),
	.V2C_2 (V2C_1015_17),
	.V2C_3 (V2C_1015_136),
	.V2C_4 (V2C_1015_150),
	.V2C_5 (V2C_1015_213),
	.V2C_6 (V2C_1015_254),
	.V (V_1015)
);

VNU_6 #(quan_width) VNU1016 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_1016),
	.C2V_2 (C2V_23_1016),
	.C2V_3 (C2V_142_1016),
	.C2V_4 (C2V_156_1016),
	.C2V_5 (C2V_219_1016),
	.C2V_6 (C2V_260_1016),
	.L (L_1016),
	.V2C_1 (V2C_1016_19),
	.V2C_2 (V2C_1016_23),
	.V2C_3 (V2C_1016_142),
	.V2C_4 (V2C_1016_156),
	.V2C_5 (V2C_1016_219),
	.V2C_6 (V2C_1016_260),
	.V (V_1016)
);

VNU_6 #(quan_width) VNU1017 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_1017),
	.C2V_2 (C2V_29_1017),
	.C2V_3 (C2V_148_1017),
	.C2V_4 (C2V_162_1017),
	.C2V_5 (C2V_225_1017),
	.C2V_6 (C2V_266_1017),
	.L (L_1017),
	.V2C_1 (V2C_1017_25),
	.V2C_2 (V2C_1017_29),
	.V2C_3 (V2C_1017_148),
	.V2C_4 (V2C_1017_162),
	.V2C_5 (V2C_1017_225),
	.V2C_6 (V2C_1017_266),
	.V (V_1017)
);

VNU_6 #(quan_width) VNU1018 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_1018),
	.C2V_2 (C2V_35_1018),
	.C2V_3 (C2V_154_1018),
	.C2V_4 (C2V_168_1018),
	.C2V_5 (C2V_231_1018),
	.C2V_6 (C2V_272_1018),
	.L (L_1018),
	.V2C_1 (V2C_1018_31),
	.V2C_2 (V2C_1018_35),
	.V2C_3 (V2C_1018_154),
	.V2C_4 (V2C_1018_168),
	.V2C_5 (V2C_1018_231),
	.V2C_6 (V2C_1018_272),
	.V (V_1018)
);

VNU_6 #(quan_width) VNU1019 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_1019),
	.C2V_2 (C2V_41_1019),
	.C2V_3 (C2V_160_1019),
	.C2V_4 (C2V_174_1019),
	.C2V_5 (C2V_237_1019),
	.C2V_6 (C2V_278_1019),
	.L (L_1019),
	.V2C_1 (V2C_1019_37),
	.V2C_2 (V2C_1019_41),
	.V2C_3 (V2C_1019_160),
	.V2C_4 (V2C_1019_174),
	.V2C_5 (V2C_1019_237),
	.V2C_6 (V2C_1019_278),
	.V (V_1019)
);

VNU_6 #(quan_width) VNU1020 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_1020),
	.C2V_2 (C2V_47_1020),
	.C2V_3 (C2V_166_1020),
	.C2V_4 (C2V_180_1020),
	.C2V_5 (C2V_243_1020),
	.C2V_6 (C2V_284_1020),
	.L (L_1020),
	.V2C_1 (V2C_1020_43),
	.V2C_2 (V2C_1020_47),
	.V2C_3 (V2C_1020_166),
	.V2C_4 (V2C_1020_180),
	.V2C_5 (V2C_1020_243),
	.V2C_6 (V2C_1020_284),
	.V (V_1020)
);

VNU_6 #(quan_width) VNU1021 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_1021),
	.C2V_2 (C2V_49_1021),
	.C2V_3 (C2V_53_1021),
	.C2V_4 (C2V_172_1021),
	.C2V_5 (C2V_186_1021),
	.C2V_6 (C2V_249_1021),
	.L (L_1021),
	.V2C_1 (V2C_1021_2),
	.V2C_2 (V2C_1021_49),
	.V2C_3 (V2C_1021_53),
	.V2C_4 (V2C_1021_172),
	.V2C_5 (V2C_1021_186),
	.V2C_6 (V2C_1021_249),
	.V (V_1021)
);

VNU_6 #(quan_width) VNU1022 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_1022),
	.C2V_2 (C2V_55_1022),
	.C2V_3 (C2V_59_1022),
	.C2V_4 (C2V_178_1022),
	.C2V_5 (C2V_192_1022),
	.C2V_6 (C2V_255_1022),
	.L (L_1022),
	.V2C_1 (V2C_1022_8),
	.V2C_2 (V2C_1022_55),
	.V2C_3 (V2C_1022_59),
	.V2C_4 (V2C_1022_178),
	.V2C_5 (V2C_1022_192),
	.V2C_6 (V2C_1022_255),
	.V (V_1022)
);

VNU_6 #(quan_width) VNU1023 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_1023),
	.C2V_2 (C2V_61_1023),
	.C2V_3 (C2V_65_1023),
	.C2V_4 (C2V_184_1023),
	.C2V_5 (C2V_198_1023),
	.C2V_6 (C2V_261_1023),
	.L (L_1023),
	.V2C_1 (V2C_1023_14),
	.V2C_2 (V2C_1023_61),
	.V2C_3 (V2C_1023_65),
	.V2C_4 (V2C_1023_184),
	.V2C_5 (V2C_1023_198),
	.V2C_6 (V2C_1023_261),
	.V (V_1023)
);

VNU_6 #(quan_width) VNU1024 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_1024),
	.C2V_2 (C2V_67_1024),
	.C2V_3 (C2V_71_1024),
	.C2V_4 (C2V_190_1024),
	.C2V_5 (C2V_204_1024),
	.C2V_6 (C2V_267_1024),
	.L (L_1024),
	.V2C_1 (V2C_1024_20),
	.V2C_2 (V2C_1024_67),
	.V2C_3 (V2C_1024_71),
	.V2C_4 (V2C_1024_190),
	.V2C_5 (V2C_1024_204),
	.V2C_6 (V2C_1024_267),
	.V (V_1024)
);

VNU_6 #(quan_width) VNU1025 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_1025),
	.C2V_2 (C2V_73_1025),
	.C2V_3 (C2V_77_1025),
	.C2V_4 (C2V_196_1025),
	.C2V_5 (C2V_210_1025),
	.C2V_6 (C2V_273_1025),
	.L (L_1025),
	.V2C_1 (V2C_1025_26),
	.V2C_2 (V2C_1025_73),
	.V2C_3 (V2C_1025_77),
	.V2C_4 (V2C_1025_196),
	.V2C_5 (V2C_1025_210),
	.V2C_6 (V2C_1025_273),
	.V (V_1025)
);

VNU_6 #(quan_width) VNU1026 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_1026),
	.C2V_2 (C2V_79_1026),
	.C2V_3 (C2V_83_1026),
	.C2V_4 (C2V_202_1026),
	.C2V_5 (C2V_216_1026),
	.C2V_6 (C2V_279_1026),
	.L (L_1026),
	.V2C_1 (V2C_1026_32),
	.V2C_2 (V2C_1026_79),
	.V2C_3 (V2C_1026_83),
	.V2C_4 (V2C_1026_202),
	.V2C_5 (V2C_1026_216),
	.V2C_6 (V2C_1026_279),
	.V (V_1026)
);

VNU_6 #(quan_width) VNU1027 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_1027),
	.C2V_2 (C2V_85_1027),
	.C2V_3 (C2V_89_1027),
	.C2V_4 (C2V_208_1027),
	.C2V_5 (C2V_222_1027),
	.C2V_6 (C2V_285_1027),
	.L (L_1027),
	.V2C_1 (V2C_1027_38),
	.V2C_2 (V2C_1027_85),
	.V2C_3 (V2C_1027_89),
	.V2C_4 (V2C_1027_208),
	.V2C_5 (V2C_1027_222),
	.V2C_6 (V2C_1027_285),
	.V (V_1027)
);

VNU_6 #(quan_width) VNU1028 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_1028),
	.C2V_2 (C2V_44_1028),
	.C2V_3 (C2V_91_1028),
	.C2V_4 (C2V_95_1028),
	.C2V_5 (C2V_214_1028),
	.C2V_6 (C2V_228_1028),
	.L (L_1028),
	.V2C_1 (V2C_1028_3),
	.V2C_2 (V2C_1028_44),
	.V2C_3 (V2C_1028_91),
	.V2C_4 (V2C_1028_95),
	.V2C_5 (V2C_1028_214),
	.V2C_6 (V2C_1028_228),
	.V (V_1028)
);

VNU_6 #(quan_width) VNU1029 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_1029),
	.C2V_2 (C2V_50_1029),
	.C2V_3 (C2V_97_1029),
	.C2V_4 (C2V_101_1029),
	.C2V_5 (C2V_220_1029),
	.C2V_6 (C2V_234_1029),
	.L (L_1029),
	.V2C_1 (V2C_1029_9),
	.V2C_2 (V2C_1029_50),
	.V2C_3 (V2C_1029_97),
	.V2C_4 (V2C_1029_101),
	.V2C_5 (V2C_1029_220),
	.V2C_6 (V2C_1029_234),
	.V (V_1029)
);

VNU_6 #(quan_width) VNU1030 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_1030),
	.C2V_2 (C2V_56_1030),
	.C2V_3 (C2V_103_1030),
	.C2V_4 (C2V_107_1030),
	.C2V_5 (C2V_226_1030),
	.C2V_6 (C2V_240_1030),
	.L (L_1030),
	.V2C_1 (V2C_1030_15),
	.V2C_2 (V2C_1030_56),
	.V2C_3 (V2C_1030_103),
	.V2C_4 (V2C_1030_107),
	.V2C_5 (V2C_1030_226),
	.V2C_6 (V2C_1030_240),
	.V (V_1030)
);

VNU_6 #(quan_width) VNU1031 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_1031),
	.C2V_2 (C2V_62_1031),
	.C2V_3 (C2V_109_1031),
	.C2V_4 (C2V_113_1031),
	.C2V_5 (C2V_232_1031),
	.C2V_6 (C2V_246_1031),
	.L (L_1031),
	.V2C_1 (V2C_1031_21),
	.V2C_2 (V2C_1031_62),
	.V2C_3 (V2C_1031_109),
	.V2C_4 (V2C_1031_113),
	.V2C_5 (V2C_1031_232),
	.V2C_6 (V2C_1031_246),
	.V (V_1031)
);

VNU_6 #(quan_width) VNU1032 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_1032),
	.C2V_2 (C2V_68_1032),
	.C2V_3 (C2V_115_1032),
	.C2V_4 (C2V_119_1032),
	.C2V_5 (C2V_238_1032),
	.C2V_6 (C2V_252_1032),
	.L (L_1032),
	.V2C_1 (V2C_1032_27),
	.V2C_2 (V2C_1032_68),
	.V2C_3 (V2C_1032_115),
	.V2C_4 (V2C_1032_119),
	.V2C_5 (V2C_1032_238),
	.V2C_6 (V2C_1032_252),
	.V (V_1032)
);

VNU_6 #(quan_width) VNU1033 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_1033),
	.C2V_2 (C2V_74_1033),
	.C2V_3 (C2V_121_1033),
	.C2V_4 (C2V_125_1033),
	.C2V_5 (C2V_244_1033),
	.C2V_6 (C2V_258_1033),
	.L (L_1033),
	.V2C_1 (V2C_1033_33),
	.V2C_2 (V2C_1033_74),
	.V2C_3 (V2C_1033_121),
	.V2C_4 (V2C_1033_125),
	.V2C_5 (V2C_1033_244),
	.V2C_6 (V2C_1033_258),
	.V (V_1033)
);

VNU_6 #(quan_width) VNU1034 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_1034),
	.C2V_2 (C2V_80_1034),
	.C2V_3 (C2V_127_1034),
	.C2V_4 (C2V_131_1034),
	.C2V_5 (C2V_250_1034),
	.C2V_6 (C2V_264_1034),
	.L (L_1034),
	.V2C_1 (V2C_1034_39),
	.V2C_2 (V2C_1034_80),
	.V2C_3 (V2C_1034_127),
	.V2C_4 (V2C_1034_131),
	.V2C_5 (V2C_1034_250),
	.V2C_6 (V2C_1034_264),
	.V (V_1034)
);

VNU_6 #(quan_width) VNU1035 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_1035),
	.C2V_2 (C2V_86_1035),
	.C2V_3 (C2V_133_1035),
	.C2V_4 (C2V_137_1035),
	.C2V_5 (C2V_256_1035),
	.C2V_6 (C2V_270_1035),
	.L (L_1035),
	.V2C_1 (V2C_1035_45),
	.V2C_2 (V2C_1035_86),
	.V2C_3 (V2C_1035_133),
	.V2C_4 (V2C_1035_137),
	.V2C_5 (V2C_1035_256),
	.V2C_6 (V2C_1035_270),
	.V (V_1035)
);

VNU_6 #(quan_width) VNU1036 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_1036),
	.C2V_2 (C2V_92_1036),
	.C2V_3 (C2V_139_1036),
	.C2V_4 (C2V_143_1036),
	.C2V_5 (C2V_262_1036),
	.C2V_6 (C2V_276_1036),
	.L (L_1036),
	.V2C_1 (V2C_1036_51),
	.V2C_2 (V2C_1036_92),
	.V2C_3 (V2C_1036_139),
	.V2C_4 (V2C_1036_143),
	.V2C_5 (V2C_1036_262),
	.V2C_6 (V2C_1036_276),
	.V (V_1036)
);

VNU_6 #(quan_width) VNU1037 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_1037),
	.C2V_2 (C2V_98_1037),
	.C2V_3 (C2V_145_1037),
	.C2V_4 (C2V_149_1037),
	.C2V_5 (C2V_268_1037),
	.C2V_6 (C2V_282_1037),
	.L (L_1037),
	.V2C_1 (V2C_1037_57),
	.V2C_2 (V2C_1037_98),
	.V2C_3 (V2C_1037_145),
	.V2C_4 (V2C_1037_149),
	.V2C_5 (V2C_1037_268),
	.V2C_6 (V2C_1037_282),
	.V (V_1037)
);

VNU_6 #(quan_width) VNU1038 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_1038),
	.C2V_2 (C2V_104_1038),
	.C2V_3 (C2V_151_1038),
	.C2V_4 (C2V_155_1038),
	.C2V_5 (C2V_274_1038),
	.C2V_6 (C2V_288_1038),
	.L (L_1038),
	.V2C_1 (V2C_1038_63),
	.V2C_2 (V2C_1038_104),
	.V2C_3 (V2C_1038_151),
	.V2C_4 (V2C_1038_155),
	.V2C_5 (V2C_1038_274),
	.V2C_6 (V2C_1038_288),
	.V (V_1038)
);

VNU_6 #(quan_width) VNU1039 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_1039),
	.C2V_2 (C2V_69_1039),
	.C2V_3 (C2V_110_1039),
	.C2V_4 (C2V_157_1039),
	.C2V_5 (C2V_161_1039),
	.C2V_6 (C2V_280_1039),
	.L (L_1039),
	.V2C_1 (V2C_1039_6),
	.V2C_2 (V2C_1039_69),
	.V2C_3 (V2C_1039_110),
	.V2C_4 (V2C_1039_157),
	.V2C_5 (V2C_1039_161),
	.V2C_6 (V2C_1039_280),
	.V (V_1039)
);

VNU_6 #(quan_width) VNU1040 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_1040),
	.C2V_2 (C2V_75_1040),
	.C2V_3 (C2V_116_1040),
	.C2V_4 (C2V_163_1040),
	.C2V_5 (C2V_167_1040),
	.C2V_6 (C2V_286_1040),
	.L (L_1040),
	.V2C_1 (V2C_1040_12),
	.V2C_2 (V2C_1040_75),
	.V2C_3 (V2C_1040_116),
	.V2C_4 (V2C_1040_163),
	.V2C_5 (V2C_1040_167),
	.V2C_6 (V2C_1040_286),
	.V (V_1040)
);

VNU_6 #(quan_width) VNU1041 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_1041),
	.C2V_2 (C2V_18_1041),
	.C2V_3 (C2V_81_1041),
	.C2V_4 (C2V_122_1041),
	.C2V_5 (C2V_169_1041),
	.C2V_6 (C2V_173_1041),
	.L (L_1041),
	.V2C_1 (V2C_1041_4),
	.V2C_2 (V2C_1041_18),
	.V2C_3 (V2C_1041_81),
	.V2C_4 (V2C_1041_122),
	.V2C_5 (V2C_1041_169),
	.V2C_6 (V2C_1041_173),
	.V (V_1041)
);

VNU_6 #(quan_width) VNU1042 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_1042),
	.C2V_2 (C2V_24_1042),
	.C2V_3 (C2V_87_1042),
	.C2V_4 (C2V_128_1042),
	.C2V_5 (C2V_175_1042),
	.C2V_6 (C2V_179_1042),
	.L (L_1042),
	.V2C_1 (V2C_1042_10),
	.V2C_2 (V2C_1042_24),
	.V2C_3 (V2C_1042_87),
	.V2C_4 (V2C_1042_128),
	.V2C_5 (V2C_1042_175),
	.V2C_6 (V2C_1042_179),
	.V (V_1042)
);

VNU_6 #(quan_width) VNU1043 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_1043),
	.C2V_2 (C2V_30_1043),
	.C2V_3 (C2V_93_1043),
	.C2V_4 (C2V_134_1043),
	.C2V_5 (C2V_181_1043),
	.C2V_6 (C2V_185_1043),
	.L (L_1043),
	.V2C_1 (V2C_1043_16),
	.V2C_2 (V2C_1043_30),
	.V2C_3 (V2C_1043_93),
	.V2C_4 (V2C_1043_134),
	.V2C_5 (V2C_1043_181),
	.V2C_6 (V2C_1043_185),
	.V (V_1043)
);

VNU_6 #(quan_width) VNU1044 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_1044),
	.C2V_2 (C2V_36_1044),
	.C2V_3 (C2V_99_1044),
	.C2V_4 (C2V_140_1044),
	.C2V_5 (C2V_187_1044),
	.C2V_6 (C2V_191_1044),
	.L (L_1044),
	.V2C_1 (V2C_1044_22),
	.V2C_2 (V2C_1044_36),
	.V2C_3 (V2C_1044_99),
	.V2C_4 (V2C_1044_140),
	.V2C_5 (V2C_1044_187),
	.V2C_6 (V2C_1044_191),
	.V (V_1044)
);

VNU_6 #(quan_width) VNU1045 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_1045),
	.C2V_2 (C2V_42_1045),
	.C2V_3 (C2V_105_1045),
	.C2V_4 (C2V_146_1045),
	.C2V_5 (C2V_193_1045),
	.C2V_6 (C2V_197_1045),
	.L (L_1045),
	.V2C_1 (V2C_1045_28),
	.V2C_2 (V2C_1045_42),
	.V2C_3 (V2C_1045_105),
	.V2C_4 (V2C_1045_146),
	.V2C_5 (V2C_1045_193),
	.V2C_6 (V2C_1045_197),
	.V (V_1045)
);

VNU_6 #(quan_width) VNU1046 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_1046),
	.C2V_2 (C2V_48_1046),
	.C2V_3 (C2V_111_1046),
	.C2V_4 (C2V_152_1046),
	.C2V_5 (C2V_199_1046),
	.C2V_6 (C2V_203_1046),
	.L (L_1046),
	.V2C_1 (V2C_1046_34),
	.V2C_2 (V2C_1046_48),
	.V2C_3 (V2C_1046_111),
	.V2C_4 (V2C_1046_152),
	.V2C_5 (V2C_1046_199),
	.V2C_6 (V2C_1046_203),
	.V (V_1046)
);

VNU_6 #(quan_width) VNU1047 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_1047),
	.C2V_2 (C2V_54_1047),
	.C2V_3 (C2V_117_1047),
	.C2V_4 (C2V_158_1047),
	.C2V_5 (C2V_205_1047),
	.C2V_6 (C2V_209_1047),
	.L (L_1047),
	.V2C_1 (V2C_1047_40),
	.V2C_2 (V2C_1047_54),
	.V2C_3 (V2C_1047_117),
	.V2C_4 (V2C_1047_158),
	.V2C_5 (V2C_1047_205),
	.V2C_6 (V2C_1047_209),
	.V (V_1047)
);

VNU_6 #(quan_width) VNU1048 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_1048),
	.C2V_2 (C2V_60_1048),
	.C2V_3 (C2V_123_1048),
	.C2V_4 (C2V_164_1048),
	.C2V_5 (C2V_211_1048),
	.C2V_6 (C2V_215_1048),
	.L (L_1048),
	.V2C_1 (V2C_1048_46),
	.V2C_2 (V2C_1048_60),
	.V2C_3 (V2C_1048_123),
	.V2C_4 (V2C_1048_164),
	.V2C_5 (V2C_1048_211),
	.V2C_6 (V2C_1048_215),
	.V (V_1048)
);

VNU_6 #(quan_width) VNU1049 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_1049),
	.C2V_2 (C2V_66_1049),
	.C2V_3 (C2V_129_1049),
	.C2V_4 (C2V_170_1049),
	.C2V_5 (C2V_217_1049),
	.C2V_6 (C2V_221_1049),
	.L (L_1049),
	.V2C_1 (V2C_1049_52),
	.V2C_2 (V2C_1049_66),
	.V2C_3 (V2C_1049_129),
	.V2C_4 (V2C_1049_170),
	.V2C_5 (V2C_1049_217),
	.V2C_6 (V2C_1049_221),
	.V (V_1049)
);

VNU_6 #(quan_width) VNU1050 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_1050),
	.C2V_2 (C2V_72_1050),
	.C2V_3 (C2V_135_1050),
	.C2V_4 (C2V_176_1050),
	.C2V_5 (C2V_223_1050),
	.C2V_6 (C2V_227_1050),
	.L (L_1050),
	.V2C_1 (V2C_1050_58),
	.V2C_2 (V2C_1050_72),
	.V2C_3 (V2C_1050_135),
	.V2C_4 (V2C_1050_176),
	.V2C_5 (V2C_1050_223),
	.V2C_6 (V2C_1050_227),
	.V (V_1050)
);

VNU_6 #(quan_width) VNU1051 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_1051),
	.C2V_2 (C2V_78_1051),
	.C2V_3 (C2V_141_1051),
	.C2V_4 (C2V_182_1051),
	.C2V_5 (C2V_229_1051),
	.C2V_6 (C2V_233_1051),
	.L (L_1051),
	.V2C_1 (V2C_1051_64),
	.V2C_2 (V2C_1051_78),
	.V2C_3 (V2C_1051_141),
	.V2C_4 (V2C_1051_182),
	.V2C_5 (V2C_1051_229),
	.V2C_6 (V2C_1051_233),
	.V (V_1051)
);

VNU_6 #(quan_width) VNU1052 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_1052),
	.C2V_2 (C2V_84_1052),
	.C2V_3 (C2V_147_1052),
	.C2V_4 (C2V_188_1052),
	.C2V_5 (C2V_235_1052),
	.C2V_6 (C2V_239_1052),
	.L (L_1052),
	.V2C_1 (V2C_1052_70),
	.V2C_2 (V2C_1052_84),
	.V2C_3 (V2C_1052_147),
	.V2C_4 (V2C_1052_188),
	.V2C_5 (V2C_1052_235),
	.V2C_6 (V2C_1052_239),
	.V (V_1052)
);

VNU_6 #(quan_width) VNU1053 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_1053),
	.C2V_2 (C2V_90_1053),
	.C2V_3 (C2V_153_1053),
	.C2V_4 (C2V_194_1053),
	.C2V_5 (C2V_241_1053),
	.C2V_6 (C2V_245_1053),
	.L (L_1053),
	.V2C_1 (V2C_1053_76),
	.V2C_2 (V2C_1053_90),
	.V2C_3 (V2C_1053_153),
	.V2C_4 (V2C_1053_194),
	.V2C_5 (V2C_1053_241),
	.V2C_6 (V2C_1053_245),
	.V (V_1053)
);

VNU_6 #(quan_width) VNU1054 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_1054),
	.C2V_2 (C2V_96_1054),
	.C2V_3 (C2V_159_1054),
	.C2V_4 (C2V_200_1054),
	.C2V_5 (C2V_247_1054),
	.C2V_6 (C2V_251_1054),
	.L (L_1054),
	.V2C_1 (V2C_1054_82),
	.V2C_2 (V2C_1054_96),
	.V2C_3 (V2C_1054_159),
	.V2C_4 (V2C_1054_200),
	.V2C_5 (V2C_1054_247),
	.V2C_6 (V2C_1054_251),
	.V (V_1054)
);

VNU_6 #(quan_width) VNU1055 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_1055),
	.C2V_2 (C2V_102_1055),
	.C2V_3 (C2V_165_1055),
	.C2V_4 (C2V_206_1055),
	.C2V_5 (C2V_253_1055),
	.C2V_6 (C2V_257_1055),
	.L (L_1055),
	.V2C_1 (V2C_1055_88),
	.V2C_2 (V2C_1055_102),
	.V2C_3 (V2C_1055_165),
	.V2C_4 (V2C_1055_206),
	.V2C_5 (V2C_1055_253),
	.V2C_6 (V2C_1055_257),
	.V (V_1055)
);

VNU_6 #(quan_width) VNU1056 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_1056),
	.C2V_2 (C2V_108_1056),
	.C2V_3 (C2V_171_1056),
	.C2V_4 (C2V_212_1056),
	.C2V_5 (C2V_259_1056),
	.C2V_6 (C2V_263_1056),
	.L (L_1056),
	.V2C_1 (V2C_1056_94),
	.V2C_2 (V2C_1056_108),
	.V2C_3 (V2C_1056_171),
	.V2C_4 (V2C_1056_212),
	.V2C_5 (V2C_1056_259),
	.V2C_6 (V2C_1056_263),
	.V (V_1056)
);

VNU_6 #(quan_width) VNU1057 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_1057),
	.C2V_2 (C2V_104_1057),
	.C2V_3 (C2V_109_1057),
	.C2V_4 (C2V_226_1057),
	.C2V_5 (C2V_263_1057),
	.C2V_6 (C2V_285_1057),
	.L (L_1057),
	.V2C_1 (V2C_1057_18),
	.V2C_2 (V2C_1057_104),
	.V2C_3 (V2C_1057_109),
	.V2C_4 (V2C_1057_226),
	.V2C_5 (V2C_1057_263),
	.V2C_6 (V2C_1057_285),
	.V (V_1057)
);

VNU_6 #(quan_width) VNU1058 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_1058),
	.C2V_2 (C2V_24_1058),
	.C2V_3 (C2V_110_1058),
	.C2V_4 (C2V_115_1058),
	.C2V_5 (C2V_232_1058),
	.C2V_6 (C2V_269_1058),
	.L (L_1058),
	.V2C_1 (V2C_1058_3),
	.V2C_2 (V2C_1058_24),
	.V2C_3 (V2C_1058_110),
	.V2C_4 (V2C_1058_115),
	.V2C_5 (V2C_1058_232),
	.V2C_6 (V2C_1058_269),
	.V (V_1058)
);

VNU_6 #(quan_width) VNU1059 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_1059),
	.C2V_2 (C2V_30_1059),
	.C2V_3 (C2V_116_1059),
	.C2V_4 (C2V_121_1059),
	.C2V_5 (C2V_238_1059),
	.C2V_6 (C2V_275_1059),
	.L (L_1059),
	.V2C_1 (V2C_1059_9),
	.V2C_2 (V2C_1059_30),
	.V2C_3 (V2C_1059_116),
	.V2C_4 (V2C_1059_121),
	.V2C_5 (V2C_1059_238),
	.V2C_6 (V2C_1059_275),
	.V (V_1059)
);

VNU_6 #(quan_width) VNU1060 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_1060),
	.C2V_2 (C2V_36_1060),
	.C2V_3 (C2V_122_1060),
	.C2V_4 (C2V_127_1060),
	.C2V_5 (C2V_244_1060),
	.C2V_6 (C2V_281_1060),
	.L (L_1060),
	.V2C_1 (V2C_1060_15),
	.V2C_2 (V2C_1060_36),
	.V2C_3 (V2C_1060_122),
	.V2C_4 (V2C_1060_127),
	.V2C_5 (V2C_1060_244),
	.V2C_6 (V2C_1060_281),
	.V (V_1060)
);

VNU_6 #(quan_width) VNU1061 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_1061),
	.C2V_2 (C2V_42_1061),
	.C2V_3 (C2V_128_1061),
	.C2V_4 (C2V_133_1061),
	.C2V_5 (C2V_250_1061),
	.C2V_6 (C2V_287_1061),
	.L (L_1061),
	.V2C_1 (V2C_1061_21),
	.V2C_2 (V2C_1061_42),
	.V2C_3 (V2C_1061_128),
	.V2C_4 (V2C_1061_133),
	.V2C_5 (V2C_1061_250),
	.V2C_6 (V2C_1061_287),
	.V (V_1061)
);

VNU_6 #(quan_width) VNU1062 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_1062),
	.C2V_2 (C2V_27_1062),
	.C2V_3 (C2V_48_1062),
	.C2V_4 (C2V_134_1062),
	.C2V_5 (C2V_139_1062),
	.C2V_6 (C2V_256_1062),
	.L (L_1062),
	.V2C_1 (V2C_1062_5),
	.V2C_2 (V2C_1062_27),
	.V2C_3 (V2C_1062_48),
	.V2C_4 (V2C_1062_134),
	.V2C_5 (V2C_1062_139),
	.V2C_6 (V2C_1062_256),
	.V (V_1062)
);

VNU_6 #(quan_width) VNU1063 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_1063),
	.C2V_2 (C2V_33_1063),
	.C2V_3 (C2V_54_1063),
	.C2V_4 (C2V_140_1063),
	.C2V_5 (C2V_145_1063),
	.C2V_6 (C2V_262_1063),
	.L (L_1063),
	.V2C_1 (V2C_1063_11),
	.V2C_2 (V2C_1063_33),
	.V2C_3 (V2C_1063_54),
	.V2C_4 (V2C_1063_140),
	.V2C_5 (V2C_1063_145),
	.V2C_6 (V2C_1063_262),
	.V (V_1063)
);

VNU_6 #(quan_width) VNU1064 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_1064),
	.C2V_2 (C2V_39_1064),
	.C2V_3 (C2V_60_1064),
	.C2V_4 (C2V_146_1064),
	.C2V_5 (C2V_151_1064),
	.C2V_6 (C2V_268_1064),
	.L (L_1064),
	.V2C_1 (V2C_1064_17),
	.V2C_2 (V2C_1064_39),
	.V2C_3 (V2C_1064_60),
	.V2C_4 (V2C_1064_146),
	.V2C_5 (V2C_1064_151),
	.V2C_6 (V2C_1064_268),
	.V (V_1064)
);

VNU_6 #(quan_width) VNU1065 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_1065),
	.C2V_2 (C2V_45_1065),
	.C2V_3 (C2V_66_1065),
	.C2V_4 (C2V_152_1065),
	.C2V_5 (C2V_157_1065),
	.C2V_6 (C2V_274_1065),
	.L (L_1065),
	.V2C_1 (V2C_1065_23),
	.V2C_2 (V2C_1065_45),
	.V2C_3 (V2C_1065_66),
	.V2C_4 (V2C_1065_152),
	.V2C_5 (V2C_1065_157),
	.V2C_6 (V2C_1065_274),
	.V (V_1065)
);

VNU_6 #(quan_width) VNU1066 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_1066),
	.C2V_2 (C2V_51_1066),
	.C2V_3 (C2V_72_1066),
	.C2V_4 (C2V_158_1066),
	.C2V_5 (C2V_163_1066),
	.C2V_6 (C2V_280_1066),
	.L (L_1066),
	.V2C_1 (V2C_1066_29),
	.V2C_2 (V2C_1066_51),
	.V2C_3 (V2C_1066_72),
	.V2C_4 (V2C_1066_158),
	.V2C_5 (V2C_1066_163),
	.V2C_6 (V2C_1066_280),
	.V (V_1066)
);

VNU_6 #(quan_width) VNU1067 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_1067),
	.C2V_2 (C2V_57_1067),
	.C2V_3 (C2V_78_1067),
	.C2V_4 (C2V_164_1067),
	.C2V_5 (C2V_169_1067),
	.C2V_6 (C2V_286_1067),
	.L (L_1067),
	.V2C_1 (V2C_1067_35),
	.V2C_2 (V2C_1067_57),
	.V2C_3 (V2C_1067_78),
	.V2C_4 (V2C_1067_164),
	.V2C_5 (V2C_1067_169),
	.V2C_6 (V2C_1067_286),
	.V (V_1067)
);

VNU_6 #(quan_width) VNU1068 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_1068),
	.C2V_2 (C2V_41_1068),
	.C2V_3 (C2V_63_1068),
	.C2V_4 (C2V_84_1068),
	.C2V_5 (C2V_170_1068),
	.C2V_6 (C2V_175_1068),
	.L (L_1068),
	.V2C_1 (V2C_1068_4),
	.V2C_2 (V2C_1068_41),
	.V2C_3 (V2C_1068_63),
	.V2C_4 (V2C_1068_84),
	.V2C_5 (V2C_1068_170),
	.V2C_6 (V2C_1068_175),
	.V (V_1068)
);

VNU_6 #(quan_width) VNU1069 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_1069),
	.C2V_2 (C2V_47_1069),
	.C2V_3 (C2V_69_1069),
	.C2V_4 (C2V_90_1069),
	.C2V_5 (C2V_176_1069),
	.C2V_6 (C2V_181_1069),
	.L (L_1069),
	.V2C_1 (V2C_1069_10),
	.V2C_2 (V2C_1069_47),
	.V2C_3 (V2C_1069_69),
	.V2C_4 (V2C_1069_90),
	.V2C_5 (V2C_1069_176),
	.V2C_6 (V2C_1069_181),
	.V (V_1069)
);

VNU_6 #(quan_width) VNU1070 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_1070),
	.C2V_2 (C2V_53_1070),
	.C2V_3 (C2V_75_1070),
	.C2V_4 (C2V_96_1070),
	.C2V_5 (C2V_182_1070),
	.C2V_6 (C2V_187_1070),
	.L (L_1070),
	.V2C_1 (V2C_1070_16),
	.V2C_2 (V2C_1070_53),
	.V2C_3 (V2C_1070_75),
	.V2C_4 (V2C_1070_96),
	.V2C_5 (V2C_1070_182),
	.V2C_6 (V2C_1070_187),
	.V (V_1070)
);

VNU_6 #(quan_width) VNU1071 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_1071),
	.C2V_2 (C2V_59_1071),
	.C2V_3 (C2V_81_1071),
	.C2V_4 (C2V_102_1071),
	.C2V_5 (C2V_188_1071),
	.C2V_6 (C2V_193_1071),
	.L (L_1071),
	.V2C_1 (V2C_1071_22),
	.V2C_2 (V2C_1071_59),
	.V2C_3 (V2C_1071_81),
	.V2C_4 (V2C_1071_102),
	.V2C_5 (V2C_1071_188),
	.V2C_6 (V2C_1071_193),
	.V (V_1071)
);

VNU_6 #(quan_width) VNU1072 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_1072),
	.C2V_2 (C2V_65_1072),
	.C2V_3 (C2V_87_1072),
	.C2V_4 (C2V_108_1072),
	.C2V_5 (C2V_194_1072),
	.C2V_6 (C2V_199_1072),
	.L (L_1072),
	.V2C_1 (V2C_1072_28),
	.V2C_2 (V2C_1072_65),
	.V2C_3 (V2C_1072_87),
	.V2C_4 (V2C_1072_108),
	.V2C_5 (V2C_1072_194),
	.V2C_6 (V2C_1072_199),
	.V (V_1072)
);

VNU_6 #(quan_width) VNU1073 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_1073),
	.C2V_2 (C2V_71_1073),
	.C2V_3 (C2V_93_1073),
	.C2V_4 (C2V_114_1073),
	.C2V_5 (C2V_200_1073),
	.C2V_6 (C2V_205_1073),
	.L (L_1073),
	.V2C_1 (V2C_1073_34),
	.V2C_2 (V2C_1073_71),
	.V2C_3 (V2C_1073_93),
	.V2C_4 (V2C_1073_114),
	.V2C_5 (V2C_1073_200),
	.V2C_6 (V2C_1073_205),
	.V (V_1073)
);

VNU_6 #(quan_width) VNU1074 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_1074),
	.C2V_2 (C2V_77_1074),
	.C2V_3 (C2V_99_1074),
	.C2V_4 (C2V_120_1074),
	.C2V_5 (C2V_206_1074),
	.C2V_6 (C2V_211_1074),
	.L (L_1074),
	.V2C_1 (V2C_1074_40),
	.V2C_2 (V2C_1074_77),
	.V2C_3 (V2C_1074_99),
	.V2C_4 (V2C_1074_120),
	.V2C_5 (V2C_1074_206),
	.V2C_6 (V2C_1074_211),
	.V (V_1074)
);

VNU_6 #(quan_width) VNU1075 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_1075),
	.C2V_2 (C2V_83_1075),
	.C2V_3 (C2V_105_1075),
	.C2V_4 (C2V_126_1075),
	.C2V_5 (C2V_212_1075),
	.C2V_6 (C2V_217_1075),
	.L (L_1075),
	.V2C_1 (V2C_1075_46),
	.V2C_2 (V2C_1075_83),
	.V2C_3 (V2C_1075_105),
	.V2C_4 (V2C_1075_126),
	.V2C_5 (V2C_1075_212),
	.V2C_6 (V2C_1075_217),
	.V (V_1075)
);

VNU_6 #(quan_width) VNU1076 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_1076),
	.C2V_2 (C2V_89_1076),
	.C2V_3 (C2V_111_1076),
	.C2V_4 (C2V_132_1076),
	.C2V_5 (C2V_218_1076),
	.C2V_6 (C2V_223_1076),
	.L (L_1076),
	.V2C_1 (V2C_1076_52),
	.V2C_2 (V2C_1076_89),
	.V2C_3 (V2C_1076_111),
	.V2C_4 (V2C_1076_132),
	.V2C_5 (V2C_1076_218),
	.V2C_6 (V2C_1076_223),
	.V (V_1076)
);

VNU_6 #(quan_width) VNU1077 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_1077),
	.C2V_2 (C2V_95_1077),
	.C2V_3 (C2V_117_1077),
	.C2V_4 (C2V_138_1077),
	.C2V_5 (C2V_224_1077),
	.C2V_6 (C2V_229_1077),
	.L (L_1077),
	.V2C_1 (V2C_1077_58),
	.V2C_2 (V2C_1077_95),
	.V2C_3 (V2C_1077_117),
	.V2C_4 (V2C_1077_138),
	.V2C_5 (V2C_1077_224),
	.V2C_6 (V2C_1077_229),
	.V (V_1077)
);

VNU_6 #(quan_width) VNU1078 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_1078),
	.C2V_2 (C2V_101_1078),
	.C2V_3 (C2V_123_1078),
	.C2V_4 (C2V_144_1078),
	.C2V_5 (C2V_230_1078),
	.C2V_6 (C2V_235_1078),
	.L (L_1078),
	.V2C_1 (V2C_1078_64),
	.V2C_2 (V2C_1078_101),
	.V2C_3 (V2C_1078_123),
	.V2C_4 (V2C_1078_144),
	.V2C_5 (V2C_1078_230),
	.V2C_6 (V2C_1078_235),
	.V (V_1078)
);

VNU_6 #(quan_width) VNU1079 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_1079),
	.C2V_2 (C2V_107_1079),
	.C2V_3 (C2V_129_1079),
	.C2V_4 (C2V_150_1079),
	.C2V_5 (C2V_236_1079),
	.C2V_6 (C2V_241_1079),
	.L (L_1079),
	.V2C_1 (V2C_1079_70),
	.V2C_2 (V2C_1079_107),
	.V2C_3 (V2C_1079_129),
	.V2C_4 (V2C_1079_150),
	.V2C_5 (V2C_1079_236),
	.V2C_6 (V2C_1079_241),
	.V (V_1079)
);

VNU_6 #(quan_width) VNU1080 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_1080),
	.C2V_2 (C2V_113_1080),
	.C2V_3 (C2V_135_1080),
	.C2V_4 (C2V_156_1080),
	.C2V_5 (C2V_242_1080),
	.C2V_6 (C2V_247_1080),
	.L (L_1080),
	.V2C_1 (V2C_1080_76),
	.V2C_2 (V2C_1080_113),
	.V2C_3 (V2C_1080_135),
	.V2C_4 (V2C_1080_156),
	.V2C_5 (V2C_1080_242),
	.V2C_6 (V2C_1080_247),
	.V (V_1080)
);

VNU_6 #(quan_width) VNU1081 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_1081),
	.C2V_2 (C2V_119_1081),
	.C2V_3 (C2V_141_1081),
	.C2V_4 (C2V_162_1081),
	.C2V_5 (C2V_248_1081),
	.C2V_6 (C2V_253_1081),
	.L (L_1081),
	.V2C_1 (V2C_1081_82),
	.V2C_2 (V2C_1081_119),
	.V2C_3 (V2C_1081_141),
	.V2C_4 (V2C_1081_162),
	.V2C_5 (V2C_1081_248),
	.V2C_6 (V2C_1081_253),
	.V (V_1081)
);

VNU_6 #(quan_width) VNU1082 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_1082),
	.C2V_2 (C2V_125_1082),
	.C2V_3 (C2V_147_1082),
	.C2V_4 (C2V_168_1082),
	.C2V_5 (C2V_254_1082),
	.C2V_6 (C2V_259_1082),
	.L (L_1082),
	.V2C_1 (V2C_1082_88),
	.V2C_2 (V2C_1082_125),
	.V2C_3 (V2C_1082_147),
	.V2C_4 (V2C_1082_168),
	.V2C_5 (V2C_1082_254),
	.V2C_6 (V2C_1082_259),
	.V (V_1082)
);

VNU_6 #(quan_width) VNU1083 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_1083),
	.C2V_2 (C2V_131_1083),
	.C2V_3 (C2V_153_1083),
	.C2V_4 (C2V_174_1083),
	.C2V_5 (C2V_260_1083),
	.C2V_6 (C2V_265_1083),
	.L (L_1083),
	.V2C_1 (V2C_1083_94),
	.V2C_2 (V2C_1083_131),
	.V2C_3 (V2C_1083_153),
	.V2C_4 (V2C_1083_174),
	.V2C_5 (V2C_1083_260),
	.V2C_6 (V2C_1083_265),
	.V (V_1083)
);

VNU_6 #(quan_width) VNU1084 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_1084),
	.C2V_2 (C2V_137_1084),
	.C2V_3 (C2V_159_1084),
	.C2V_4 (C2V_180_1084),
	.C2V_5 (C2V_266_1084),
	.C2V_6 (C2V_271_1084),
	.L (L_1084),
	.V2C_1 (V2C_1084_100),
	.V2C_2 (V2C_1084_137),
	.V2C_3 (V2C_1084_159),
	.V2C_4 (V2C_1084_180),
	.V2C_5 (V2C_1084_266),
	.V2C_6 (V2C_1084_271),
	.V (V_1084)
);

VNU_6 #(quan_width) VNU1085 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_1085),
	.C2V_2 (C2V_143_1085),
	.C2V_3 (C2V_165_1085),
	.C2V_4 (C2V_186_1085),
	.C2V_5 (C2V_272_1085),
	.C2V_6 (C2V_277_1085),
	.L (L_1085),
	.V2C_1 (V2C_1085_106),
	.V2C_2 (V2C_1085_143),
	.V2C_3 (V2C_1085_165),
	.V2C_4 (V2C_1085_186),
	.V2C_5 (V2C_1085_272),
	.V2C_6 (V2C_1085_277),
	.V (V_1085)
);

VNU_6 #(quan_width) VNU1086 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_1086),
	.C2V_2 (C2V_149_1086),
	.C2V_3 (C2V_171_1086),
	.C2V_4 (C2V_192_1086),
	.C2V_5 (C2V_278_1086),
	.C2V_6 (C2V_283_1086),
	.L (L_1086),
	.V2C_1 (V2C_1086_112),
	.V2C_2 (V2C_1086_149),
	.V2C_3 (V2C_1086_171),
	.V2C_4 (V2C_1086_192),
	.V2C_5 (V2C_1086_278),
	.V2C_6 (V2C_1086_283),
	.V (V_1086)
);

VNU_6 #(quan_width) VNU1087 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_1087),
	.C2V_2 (C2V_118_1087),
	.C2V_3 (C2V_155_1087),
	.C2V_4 (C2V_177_1087),
	.C2V_5 (C2V_198_1087),
	.C2V_6 (C2V_284_1087),
	.L (L_1087),
	.V2C_1 (V2C_1087_1),
	.V2C_2 (V2C_1087_118),
	.V2C_3 (V2C_1087_155),
	.V2C_4 (V2C_1087_177),
	.V2C_5 (V2C_1087_198),
	.V2C_6 (V2C_1087_284),
	.V (V_1087)
);

VNU_6 #(quan_width) VNU1088 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_1088),
	.C2V_2 (C2V_7_1088),
	.C2V_3 (C2V_124_1088),
	.C2V_4 (C2V_161_1088),
	.C2V_5 (C2V_183_1088),
	.C2V_6 (C2V_204_1088),
	.L (L_1088),
	.V2C_1 (V2C_1088_2),
	.V2C_2 (V2C_1088_7),
	.V2C_3 (V2C_1088_124),
	.V2C_4 (V2C_1088_161),
	.V2C_5 (V2C_1088_183),
	.V2C_6 (V2C_1088_204),
	.V (V_1088)
);

VNU_6 #(quan_width) VNU1089 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_1089),
	.C2V_2 (C2V_13_1089),
	.C2V_3 (C2V_130_1089),
	.C2V_4 (C2V_167_1089),
	.C2V_5 (C2V_189_1089),
	.C2V_6 (C2V_210_1089),
	.L (L_1089),
	.V2C_1 (V2C_1089_8),
	.V2C_2 (V2C_1089_13),
	.V2C_3 (V2C_1089_130),
	.V2C_4 (V2C_1089_167),
	.V2C_5 (V2C_1089_189),
	.V2C_6 (V2C_1089_210),
	.V (V_1089)
);

VNU_6 #(quan_width) VNU1090 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_1090),
	.C2V_2 (C2V_19_1090),
	.C2V_3 (C2V_136_1090),
	.C2V_4 (C2V_173_1090),
	.C2V_5 (C2V_195_1090),
	.C2V_6 (C2V_216_1090),
	.L (L_1090),
	.V2C_1 (V2C_1090_14),
	.V2C_2 (V2C_1090_19),
	.V2C_3 (V2C_1090_136),
	.V2C_4 (V2C_1090_173),
	.V2C_5 (V2C_1090_195),
	.V2C_6 (V2C_1090_216),
	.V (V_1090)
);

VNU_6 #(quan_width) VNU1091 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_1091),
	.C2V_2 (C2V_25_1091),
	.C2V_3 (C2V_142_1091),
	.C2V_4 (C2V_179_1091),
	.C2V_5 (C2V_201_1091),
	.C2V_6 (C2V_222_1091),
	.L (L_1091),
	.V2C_1 (V2C_1091_20),
	.V2C_2 (V2C_1091_25),
	.V2C_3 (V2C_1091_142),
	.V2C_4 (V2C_1091_179),
	.V2C_5 (V2C_1091_201),
	.V2C_6 (V2C_1091_222),
	.V (V_1091)
);

VNU_6 #(quan_width) VNU1092 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_1092),
	.C2V_2 (C2V_31_1092),
	.C2V_3 (C2V_148_1092),
	.C2V_4 (C2V_185_1092),
	.C2V_5 (C2V_207_1092),
	.C2V_6 (C2V_228_1092),
	.L (L_1092),
	.V2C_1 (V2C_1092_26),
	.V2C_2 (V2C_1092_31),
	.V2C_3 (V2C_1092_148),
	.V2C_4 (V2C_1092_185),
	.V2C_5 (V2C_1092_207),
	.V2C_6 (V2C_1092_228),
	.V (V_1092)
);

VNU_6 #(quan_width) VNU1093 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_1093),
	.C2V_2 (C2V_37_1093),
	.C2V_3 (C2V_154_1093),
	.C2V_4 (C2V_191_1093),
	.C2V_5 (C2V_213_1093),
	.C2V_6 (C2V_234_1093),
	.L (L_1093),
	.V2C_1 (V2C_1093_32),
	.V2C_2 (V2C_1093_37),
	.V2C_3 (V2C_1093_154),
	.V2C_4 (V2C_1093_191),
	.V2C_5 (V2C_1093_213),
	.V2C_6 (V2C_1093_234),
	.V (V_1093)
);

VNU_6 #(quan_width) VNU1094 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_1094),
	.C2V_2 (C2V_43_1094),
	.C2V_3 (C2V_160_1094),
	.C2V_4 (C2V_197_1094),
	.C2V_5 (C2V_219_1094),
	.C2V_6 (C2V_240_1094),
	.L (L_1094),
	.V2C_1 (V2C_1094_38),
	.V2C_2 (V2C_1094_43),
	.V2C_3 (V2C_1094_160),
	.V2C_4 (V2C_1094_197),
	.V2C_5 (V2C_1094_219),
	.V2C_6 (V2C_1094_240),
	.V (V_1094)
);

VNU_6 #(quan_width) VNU1095 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_1095),
	.C2V_2 (C2V_49_1095),
	.C2V_3 (C2V_166_1095),
	.C2V_4 (C2V_203_1095),
	.C2V_5 (C2V_225_1095),
	.C2V_6 (C2V_246_1095),
	.L (L_1095),
	.V2C_1 (V2C_1095_44),
	.V2C_2 (V2C_1095_49),
	.V2C_3 (V2C_1095_166),
	.V2C_4 (V2C_1095_203),
	.V2C_5 (V2C_1095_225),
	.V2C_6 (V2C_1095_246),
	.V (V_1095)
);

VNU_6 #(quan_width) VNU1096 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_1096),
	.C2V_2 (C2V_55_1096),
	.C2V_3 (C2V_172_1096),
	.C2V_4 (C2V_209_1096),
	.C2V_5 (C2V_231_1096),
	.C2V_6 (C2V_252_1096),
	.L (L_1096),
	.V2C_1 (V2C_1096_50),
	.V2C_2 (V2C_1096_55),
	.V2C_3 (V2C_1096_172),
	.V2C_4 (V2C_1096_209),
	.V2C_5 (V2C_1096_231),
	.V2C_6 (V2C_1096_252),
	.V (V_1096)
);

VNU_6 #(quan_width) VNU1097 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_1097),
	.C2V_2 (C2V_61_1097),
	.C2V_3 (C2V_178_1097),
	.C2V_4 (C2V_215_1097),
	.C2V_5 (C2V_237_1097),
	.C2V_6 (C2V_258_1097),
	.L (L_1097),
	.V2C_1 (V2C_1097_56),
	.V2C_2 (V2C_1097_61),
	.V2C_3 (V2C_1097_178),
	.V2C_4 (V2C_1097_215),
	.V2C_5 (V2C_1097_237),
	.V2C_6 (V2C_1097_258),
	.V (V_1097)
);

VNU_6 #(quan_width) VNU1098 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_1098),
	.C2V_2 (C2V_67_1098),
	.C2V_3 (C2V_184_1098),
	.C2V_4 (C2V_221_1098),
	.C2V_5 (C2V_243_1098),
	.C2V_6 (C2V_264_1098),
	.L (L_1098),
	.V2C_1 (V2C_1098_62),
	.V2C_2 (V2C_1098_67),
	.V2C_3 (V2C_1098_184),
	.V2C_4 (V2C_1098_221),
	.V2C_5 (V2C_1098_243),
	.V2C_6 (V2C_1098_264),
	.V (V_1098)
);

VNU_6 #(quan_width) VNU1099 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_1099),
	.C2V_2 (C2V_73_1099),
	.C2V_3 (C2V_190_1099),
	.C2V_4 (C2V_227_1099),
	.C2V_5 (C2V_249_1099),
	.C2V_6 (C2V_270_1099),
	.L (L_1099),
	.V2C_1 (V2C_1099_68),
	.V2C_2 (V2C_1099_73),
	.V2C_3 (V2C_1099_190),
	.V2C_4 (V2C_1099_227),
	.V2C_5 (V2C_1099_249),
	.V2C_6 (V2C_1099_270),
	.V (V_1099)
);

VNU_6 #(quan_width) VNU1100 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_1100),
	.C2V_2 (C2V_79_1100),
	.C2V_3 (C2V_196_1100),
	.C2V_4 (C2V_233_1100),
	.C2V_5 (C2V_255_1100),
	.C2V_6 (C2V_276_1100),
	.L (L_1100),
	.V2C_1 (V2C_1100_74),
	.V2C_2 (V2C_1100_79),
	.V2C_3 (V2C_1100_196),
	.V2C_4 (V2C_1100_233),
	.V2C_5 (V2C_1100_255),
	.V2C_6 (V2C_1100_276),
	.V (V_1100)
);

VNU_6 #(quan_width) VNU1101 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_80_1101),
	.C2V_2 (C2V_85_1101),
	.C2V_3 (C2V_202_1101),
	.C2V_4 (C2V_239_1101),
	.C2V_5 (C2V_261_1101),
	.C2V_6 (C2V_282_1101),
	.L (L_1101),
	.V2C_1 (V2C_1101_80),
	.V2C_2 (V2C_1101_85),
	.V2C_3 (V2C_1101_202),
	.V2C_4 (V2C_1101_239),
	.V2C_5 (V2C_1101_261),
	.V2C_6 (V2C_1101_282),
	.V (V_1101)
);

VNU_6 #(quan_width) VNU1102 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_86_1102),
	.C2V_2 (C2V_91_1102),
	.C2V_3 (C2V_208_1102),
	.C2V_4 (C2V_245_1102),
	.C2V_5 (C2V_267_1102),
	.C2V_6 (C2V_288_1102),
	.L (L_1102),
	.V2C_1 (V2C_1102_86),
	.V2C_2 (V2C_1102_91),
	.V2C_3 (V2C_1102_208),
	.V2C_4 (V2C_1102_245),
	.V2C_5 (V2C_1102_267),
	.V2C_6 (V2C_1102_288),
	.V (V_1102)
);

VNU_6 #(quan_width) VNU1103 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_1103),
	.C2V_2 (C2V_92_1103),
	.C2V_3 (C2V_97_1103),
	.C2V_4 (C2V_214_1103),
	.C2V_5 (C2V_251_1103),
	.C2V_6 (C2V_273_1103),
	.L (L_1103),
	.V2C_1 (V2C_1103_6),
	.V2C_2 (V2C_1103_92),
	.V2C_3 (V2C_1103_97),
	.V2C_4 (V2C_1103_214),
	.V2C_5 (V2C_1103_251),
	.V2C_6 (V2C_1103_273),
	.V (V_1103)
);

VNU_6 #(quan_width) VNU1104 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_1104),
	.C2V_2 (C2V_98_1104),
	.C2V_3 (C2V_103_1104),
	.C2V_4 (C2V_220_1104),
	.C2V_5 (C2V_257_1104),
	.C2V_6 (C2V_279_1104),
	.L (L_1104),
	.V2C_1 (V2C_1104_12),
	.V2C_2 (V2C_1104_98),
	.V2C_3 (V2C_1104_103),
	.V2C_4 (V2C_1104_220),
	.V2C_5 (V2C_1104_257),
	.V2C_6 (V2C_1104_279),
	.V (V_1104)
);

VNU_6 #(quan_width) VNU1105 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_1105),
	.C2V_2 (C2V_15_1105),
	.C2V_3 (C2V_43_1105),
	.C2V_4 (C2V_130_1105),
	.C2V_5 (C2V_206_1105),
	.C2V_6 (C2V_263_1105),
	.L (L_1105),
	.V2C_1 (V2C_1105_6),
	.V2C_2 (V2C_1105_15),
	.V2C_3 (V2C_1105_43),
	.V2C_4 (V2C_1105_130),
	.V2C_5 (V2C_1105_206),
	.V2C_6 (V2C_1105_263),
	.V (V_1105)
);

VNU_6 #(quan_width) VNU1106 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_1106),
	.C2V_2 (C2V_21_1106),
	.C2V_3 (C2V_49_1106),
	.C2V_4 (C2V_136_1106),
	.C2V_5 (C2V_212_1106),
	.C2V_6 (C2V_269_1106),
	.L (L_1106),
	.V2C_1 (V2C_1106_12),
	.V2C_2 (V2C_1106_21),
	.V2C_3 (V2C_1106_49),
	.V2C_4 (V2C_1106_136),
	.V2C_5 (V2C_1106_212),
	.V2C_6 (V2C_1106_269),
	.V (V_1106)
);

VNU_6 #(quan_width) VNU1107 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_1107),
	.C2V_2 (C2V_27_1107),
	.C2V_3 (C2V_55_1107),
	.C2V_4 (C2V_142_1107),
	.C2V_5 (C2V_218_1107),
	.C2V_6 (C2V_275_1107),
	.L (L_1107),
	.V2C_1 (V2C_1107_18),
	.V2C_2 (V2C_1107_27),
	.V2C_3 (V2C_1107_55),
	.V2C_4 (V2C_1107_142),
	.V2C_5 (V2C_1107_218),
	.V2C_6 (V2C_1107_275),
	.V (V_1107)
);

VNU_6 #(quan_width) VNU1108 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_1108),
	.C2V_2 (C2V_33_1108),
	.C2V_3 (C2V_61_1108),
	.C2V_4 (C2V_148_1108),
	.C2V_5 (C2V_224_1108),
	.C2V_6 (C2V_281_1108),
	.L (L_1108),
	.V2C_1 (V2C_1108_24),
	.V2C_2 (V2C_1108_33),
	.V2C_3 (V2C_1108_61),
	.V2C_4 (V2C_1108_148),
	.V2C_5 (V2C_1108_224),
	.V2C_6 (V2C_1108_281),
	.V (V_1108)
);

VNU_6 #(quan_width) VNU1109 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_1109),
	.C2V_2 (C2V_39_1109),
	.C2V_3 (C2V_67_1109),
	.C2V_4 (C2V_154_1109),
	.C2V_5 (C2V_230_1109),
	.C2V_6 (C2V_287_1109),
	.L (L_1109),
	.V2C_1 (V2C_1109_30),
	.V2C_2 (V2C_1109_39),
	.V2C_3 (V2C_1109_67),
	.V2C_4 (V2C_1109_154),
	.V2C_5 (V2C_1109_230),
	.V2C_6 (V2C_1109_287),
	.V (V_1109)
);

VNU_6 #(quan_width) VNU1110 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_1110),
	.C2V_2 (C2V_36_1110),
	.C2V_3 (C2V_45_1110),
	.C2V_4 (C2V_73_1110),
	.C2V_5 (C2V_160_1110),
	.C2V_6 (C2V_236_1110),
	.L (L_1110),
	.V2C_1 (V2C_1110_5),
	.V2C_2 (V2C_1110_36),
	.V2C_3 (V2C_1110_45),
	.V2C_4 (V2C_1110_73),
	.V2C_5 (V2C_1110_160),
	.V2C_6 (V2C_1110_236),
	.V (V_1110)
);

VNU_6 #(quan_width) VNU1111 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_1111),
	.C2V_2 (C2V_42_1111),
	.C2V_3 (C2V_51_1111),
	.C2V_4 (C2V_79_1111),
	.C2V_5 (C2V_166_1111),
	.C2V_6 (C2V_242_1111),
	.L (L_1111),
	.V2C_1 (V2C_1111_11),
	.V2C_2 (V2C_1111_42),
	.V2C_3 (V2C_1111_51),
	.V2C_4 (V2C_1111_79),
	.V2C_5 (V2C_1111_166),
	.V2C_6 (V2C_1111_242),
	.V (V_1111)
);

VNU_6 #(quan_width) VNU1112 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_1112),
	.C2V_2 (C2V_48_1112),
	.C2V_3 (C2V_57_1112),
	.C2V_4 (C2V_85_1112),
	.C2V_5 (C2V_172_1112),
	.C2V_6 (C2V_248_1112),
	.L (L_1112),
	.V2C_1 (V2C_1112_17),
	.V2C_2 (V2C_1112_48),
	.V2C_3 (V2C_1112_57),
	.V2C_4 (V2C_1112_85),
	.V2C_5 (V2C_1112_172),
	.V2C_6 (V2C_1112_248),
	.V (V_1112)
);

VNU_6 #(quan_width) VNU1113 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_1113),
	.C2V_2 (C2V_54_1113),
	.C2V_3 (C2V_63_1113),
	.C2V_4 (C2V_91_1113),
	.C2V_5 (C2V_178_1113),
	.C2V_6 (C2V_254_1113),
	.L (L_1113),
	.V2C_1 (V2C_1113_23),
	.V2C_2 (V2C_1113_54),
	.V2C_3 (V2C_1113_63),
	.V2C_4 (V2C_1113_91),
	.V2C_5 (V2C_1113_178),
	.V2C_6 (V2C_1113_254),
	.V (V_1113)
);

VNU_6 #(quan_width) VNU1114 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_1114),
	.C2V_2 (C2V_60_1114),
	.C2V_3 (C2V_69_1114),
	.C2V_4 (C2V_97_1114),
	.C2V_5 (C2V_184_1114),
	.C2V_6 (C2V_260_1114),
	.L (L_1114),
	.V2C_1 (V2C_1114_29),
	.V2C_2 (V2C_1114_60),
	.V2C_3 (V2C_1114_69),
	.V2C_4 (V2C_1114_97),
	.V2C_5 (V2C_1114_184),
	.V2C_6 (V2C_1114_260),
	.V (V_1114)
);

VNU_6 #(quan_width) VNU1115 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_1115),
	.C2V_2 (C2V_66_1115),
	.C2V_3 (C2V_75_1115),
	.C2V_4 (C2V_103_1115),
	.C2V_5 (C2V_190_1115),
	.C2V_6 (C2V_266_1115),
	.L (L_1115),
	.V2C_1 (V2C_1115_35),
	.V2C_2 (V2C_1115_66),
	.V2C_3 (V2C_1115_75),
	.V2C_4 (V2C_1115_103),
	.V2C_5 (V2C_1115_190),
	.V2C_6 (V2C_1115_266),
	.V (V_1115)
);

VNU_6 #(quan_width) VNU1116 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_1116),
	.C2V_2 (C2V_72_1116),
	.C2V_3 (C2V_81_1116),
	.C2V_4 (C2V_109_1116),
	.C2V_5 (C2V_196_1116),
	.C2V_6 (C2V_272_1116),
	.L (L_1116),
	.V2C_1 (V2C_1116_41),
	.V2C_2 (V2C_1116_72),
	.V2C_3 (V2C_1116_81),
	.V2C_4 (V2C_1116_109),
	.V2C_5 (V2C_1116_196),
	.V2C_6 (V2C_1116_272),
	.V (V_1116)
);

VNU_6 #(quan_width) VNU1117 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_1117),
	.C2V_2 (C2V_78_1117),
	.C2V_3 (C2V_87_1117),
	.C2V_4 (C2V_115_1117),
	.C2V_5 (C2V_202_1117),
	.C2V_6 (C2V_278_1117),
	.L (L_1117),
	.V2C_1 (V2C_1117_47),
	.V2C_2 (V2C_1117_78),
	.V2C_3 (V2C_1117_87),
	.V2C_4 (V2C_1117_115),
	.V2C_5 (V2C_1117_202),
	.V2C_6 (V2C_1117_278),
	.V (V_1117)
);

VNU_6 #(quan_width) VNU1118 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_1118),
	.C2V_2 (C2V_84_1118),
	.C2V_3 (C2V_93_1118),
	.C2V_4 (C2V_121_1118),
	.C2V_5 (C2V_208_1118),
	.C2V_6 (C2V_284_1118),
	.L (L_1118),
	.V2C_1 (V2C_1118_53),
	.V2C_2 (V2C_1118_84),
	.V2C_3 (V2C_1118_93),
	.V2C_4 (V2C_1118_121),
	.V2C_5 (V2C_1118_208),
	.V2C_6 (V2C_1118_284),
	.V (V_1118)
);

VNU_6 #(quan_width) VNU1119 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_1119),
	.C2V_2 (C2V_59_1119),
	.C2V_3 (C2V_90_1119),
	.C2V_4 (C2V_99_1119),
	.C2V_5 (C2V_127_1119),
	.C2V_6 (C2V_214_1119),
	.L (L_1119),
	.V2C_1 (V2C_1119_2),
	.V2C_2 (V2C_1119_59),
	.V2C_3 (V2C_1119_90),
	.V2C_4 (V2C_1119_99),
	.V2C_5 (V2C_1119_127),
	.V2C_6 (V2C_1119_214),
	.V (V_1119)
);

VNU_6 #(quan_width) VNU1120 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_1120),
	.C2V_2 (C2V_65_1120),
	.C2V_3 (C2V_96_1120),
	.C2V_4 (C2V_105_1120),
	.C2V_5 (C2V_133_1120),
	.C2V_6 (C2V_220_1120),
	.L (L_1120),
	.V2C_1 (V2C_1120_8),
	.V2C_2 (V2C_1120_65),
	.V2C_3 (V2C_1120_96),
	.V2C_4 (V2C_1120_105),
	.V2C_5 (V2C_1120_133),
	.V2C_6 (V2C_1120_220),
	.V (V_1120)
);

VNU_6 #(quan_width) VNU1121 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_1121),
	.C2V_2 (C2V_71_1121),
	.C2V_3 (C2V_102_1121),
	.C2V_4 (C2V_111_1121),
	.C2V_5 (C2V_139_1121),
	.C2V_6 (C2V_226_1121),
	.L (L_1121),
	.V2C_1 (V2C_1121_14),
	.V2C_2 (V2C_1121_71),
	.V2C_3 (V2C_1121_102),
	.V2C_4 (V2C_1121_111),
	.V2C_5 (V2C_1121_139),
	.V2C_6 (V2C_1121_226),
	.V (V_1121)
);

VNU_6 #(quan_width) VNU1122 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_1122),
	.C2V_2 (C2V_77_1122),
	.C2V_3 (C2V_108_1122),
	.C2V_4 (C2V_117_1122),
	.C2V_5 (C2V_145_1122),
	.C2V_6 (C2V_232_1122),
	.L (L_1122),
	.V2C_1 (V2C_1122_20),
	.V2C_2 (V2C_1122_77),
	.V2C_3 (V2C_1122_108),
	.V2C_4 (V2C_1122_117),
	.V2C_5 (V2C_1122_145),
	.V2C_6 (V2C_1122_232),
	.V (V_1122)
);

VNU_6 #(quan_width) VNU1123 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_1123),
	.C2V_2 (C2V_83_1123),
	.C2V_3 (C2V_114_1123),
	.C2V_4 (C2V_123_1123),
	.C2V_5 (C2V_151_1123),
	.C2V_6 (C2V_238_1123),
	.L (L_1123),
	.V2C_1 (V2C_1123_26),
	.V2C_2 (V2C_1123_83),
	.V2C_3 (V2C_1123_114),
	.V2C_4 (V2C_1123_123),
	.V2C_5 (V2C_1123_151),
	.V2C_6 (V2C_1123_238),
	.V (V_1123)
);

VNU_6 #(quan_width) VNU1124 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_1124),
	.C2V_2 (C2V_89_1124),
	.C2V_3 (C2V_120_1124),
	.C2V_4 (C2V_129_1124),
	.C2V_5 (C2V_157_1124),
	.C2V_6 (C2V_244_1124),
	.L (L_1124),
	.V2C_1 (V2C_1124_32),
	.V2C_2 (V2C_1124_89),
	.V2C_3 (V2C_1124_120),
	.V2C_4 (V2C_1124_129),
	.V2C_5 (V2C_1124_157),
	.V2C_6 (V2C_1124_244),
	.V (V_1124)
);

VNU_6 #(quan_width) VNU1125 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_1125),
	.C2V_2 (C2V_95_1125),
	.C2V_3 (C2V_126_1125),
	.C2V_4 (C2V_135_1125),
	.C2V_5 (C2V_163_1125),
	.C2V_6 (C2V_250_1125),
	.L (L_1125),
	.V2C_1 (V2C_1125_38),
	.V2C_2 (V2C_1125_95),
	.V2C_3 (V2C_1125_126),
	.V2C_4 (V2C_1125_135),
	.V2C_5 (V2C_1125_163),
	.V2C_6 (V2C_1125_250),
	.V (V_1125)
);

VNU_6 #(quan_width) VNU1126 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_1126),
	.C2V_2 (C2V_101_1126),
	.C2V_3 (C2V_132_1126),
	.C2V_4 (C2V_141_1126),
	.C2V_5 (C2V_169_1126),
	.C2V_6 (C2V_256_1126),
	.L (L_1126),
	.V2C_1 (V2C_1126_44),
	.V2C_2 (V2C_1126_101),
	.V2C_3 (V2C_1126_132),
	.V2C_4 (V2C_1126_141),
	.V2C_5 (V2C_1126_169),
	.V2C_6 (V2C_1126_256),
	.V (V_1126)
);

VNU_6 #(quan_width) VNU1127 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_1127),
	.C2V_2 (C2V_107_1127),
	.C2V_3 (C2V_138_1127),
	.C2V_4 (C2V_147_1127),
	.C2V_5 (C2V_175_1127),
	.C2V_6 (C2V_262_1127),
	.L (L_1127),
	.V2C_1 (V2C_1127_50),
	.V2C_2 (V2C_1127_107),
	.V2C_3 (V2C_1127_138),
	.V2C_4 (V2C_1127_147),
	.V2C_5 (V2C_1127_175),
	.V2C_6 (V2C_1127_262),
	.V (V_1127)
);

VNU_6 #(quan_width) VNU1128 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_1128),
	.C2V_2 (C2V_113_1128),
	.C2V_3 (C2V_144_1128),
	.C2V_4 (C2V_153_1128),
	.C2V_5 (C2V_181_1128),
	.C2V_6 (C2V_268_1128),
	.L (L_1128),
	.V2C_1 (V2C_1128_56),
	.V2C_2 (V2C_1128_113),
	.V2C_3 (V2C_1128_144),
	.V2C_4 (V2C_1128_153),
	.V2C_5 (V2C_1128_181),
	.V2C_6 (V2C_1128_268),
	.V (V_1128)
);

VNU_6 #(quan_width) VNU1129 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_1129),
	.C2V_2 (C2V_119_1129),
	.C2V_3 (C2V_150_1129),
	.C2V_4 (C2V_159_1129),
	.C2V_5 (C2V_187_1129),
	.C2V_6 (C2V_274_1129),
	.L (L_1129),
	.V2C_1 (V2C_1129_62),
	.V2C_2 (V2C_1129_119),
	.V2C_3 (V2C_1129_150),
	.V2C_4 (V2C_1129_159),
	.V2C_5 (V2C_1129_187),
	.V2C_6 (V2C_1129_274),
	.V (V_1129)
);

VNU_6 #(quan_width) VNU1130 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_1130),
	.C2V_2 (C2V_125_1130),
	.C2V_3 (C2V_156_1130),
	.C2V_4 (C2V_165_1130),
	.C2V_5 (C2V_193_1130),
	.C2V_6 (C2V_280_1130),
	.L (L_1130),
	.V2C_1 (V2C_1130_68),
	.V2C_2 (V2C_1130_125),
	.V2C_3 (V2C_1130_156),
	.V2C_4 (V2C_1130_165),
	.V2C_5 (V2C_1130_193),
	.V2C_6 (V2C_1130_280),
	.V (V_1130)
);

VNU_6 #(quan_width) VNU1131 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_1131),
	.C2V_2 (C2V_131_1131),
	.C2V_3 (C2V_162_1131),
	.C2V_4 (C2V_171_1131),
	.C2V_5 (C2V_199_1131),
	.C2V_6 (C2V_286_1131),
	.L (L_1131),
	.V2C_1 (V2C_1131_74),
	.V2C_2 (V2C_1131_131),
	.V2C_3 (V2C_1131_162),
	.V2C_4 (V2C_1131_171),
	.V2C_5 (V2C_1131_199),
	.V2C_6 (V2C_1131_286),
	.V (V_1131)
);

VNU_6 #(quan_width) VNU1132 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_1132),
	.C2V_2 (C2V_80_1132),
	.C2V_3 (C2V_137_1132),
	.C2V_4 (C2V_168_1132),
	.C2V_5 (C2V_177_1132),
	.C2V_6 (C2V_205_1132),
	.L (L_1132),
	.V2C_1 (V2C_1132_4),
	.V2C_2 (V2C_1132_80),
	.V2C_3 (V2C_1132_137),
	.V2C_4 (V2C_1132_168),
	.V2C_5 (V2C_1132_177),
	.V2C_6 (V2C_1132_205),
	.V (V_1132)
);

VNU_6 #(quan_width) VNU1133 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_1133),
	.C2V_2 (C2V_86_1133),
	.C2V_3 (C2V_143_1133),
	.C2V_4 (C2V_174_1133),
	.C2V_5 (C2V_183_1133),
	.C2V_6 (C2V_211_1133),
	.L (L_1133),
	.V2C_1 (V2C_1133_10),
	.V2C_2 (V2C_1133_86),
	.V2C_3 (V2C_1133_143),
	.V2C_4 (V2C_1133_174),
	.V2C_5 (V2C_1133_183),
	.V2C_6 (V2C_1133_211),
	.V (V_1133)
);

VNU_6 #(quan_width) VNU1134 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_1134),
	.C2V_2 (C2V_92_1134),
	.C2V_3 (C2V_149_1134),
	.C2V_4 (C2V_180_1134),
	.C2V_5 (C2V_189_1134),
	.C2V_6 (C2V_217_1134),
	.L (L_1134),
	.V2C_1 (V2C_1134_16),
	.V2C_2 (V2C_1134_92),
	.V2C_3 (V2C_1134_149),
	.V2C_4 (V2C_1134_180),
	.V2C_5 (V2C_1134_189),
	.V2C_6 (V2C_1134_217),
	.V (V_1134)
);

VNU_6 #(quan_width) VNU1135 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_1135),
	.C2V_2 (C2V_98_1135),
	.C2V_3 (C2V_155_1135),
	.C2V_4 (C2V_186_1135),
	.C2V_5 (C2V_195_1135),
	.C2V_6 (C2V_223_1135),
	.L (L_1135),
	.V2C_1 (V2C_1135_22),
	.V2C_2 (V2C_1135_98),
	.V2C_3 (V2C_1135_155),
	.V2C_4 (V2C_1135_186),
	.V2C_5 (V2C_1135_195),
	.V2C_6 (V2C_1135_223),
	.V (V_1135)
);

VNU_6 #(quan_width) VNU1136 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_1136),
	.C2V_2 (C2V_104_1136),
	.C2V_3 (C2V_161_1136),
	.C2V_4 (C2V_192_1136),
	.C2V_5 (C2V_201_1136),
	.C2V_6 (C2V_229_1136),
	.L (L_1136),
	.V2C_1 (V2C_1136_28),
	.V2C_2 (V2C_1136_104),
	.V2C_3 (V2C_1136_161),
	.V2C_4 (V2C_1136_192),
	.V2C_5 (V2C_1136_201),
	.V2C_6 (V2C_1136_229),
	.V (V_1136)
);

VNU_6 #(quan_width) VNU1137 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_1137),
	.C2V_2 (C2V_110_1137),
	.C2V_3 (C2V_167_1137),
	.C2V_4 (C2V_198_1137),
	.C2V_5 (C2V_207_1137),
	.C2V_6 (C2V_235_1137),
	.L (L_1137),
	.V2C_1 (V2C_1137_34),
	.V2C_2 (V2C_1137_110),
	.V2C_3 (V2C_1137_167),
	.V2C_4 (V2C_1137_198),
	.V2C_5 (V2C_1137_207),
	.V2C_6 (V2C_1137_235),
	.V (V_1137)
);

VNU_6 #(quan_width) VNU1138 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_1138),
	.C2V_2 (C2V_116_1138),
	.C2V_3 (C2V_173_1138),
	.C2V_4 (C2V_204_1138),
	.C2V_5 (C2V_213_1138),
	.C2V_6 (C2V_241_1138),
	.L (L_1138),
	.V2C_1 (V2C_1138_40),
	.V2C_2 (V2C_1138_116),
	.V2C_3 (V2C_1138_173),
	.V2C_4 (V2C_1138_204),
	.V2C_5 (V2C_1138_213),
	.V2C_6 (V2C_1138_241),
	.V (V_1138)
);

VNU_6 #(quan_width) VNU1139 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_1139),
	.C2V_2 (C2V_122_1139),
	.C2V_3 (C2V_179_1139),
	.C2V_4 (C2V_210_1139),
	.C2V_5 (C2V_219_1139),
	.C2V_6 (C2V_247_1139),
	.L (L_1139),
	.V2C_1 (V2C_1139_46),
	.V2C_2 (V2C_1139_122),
	.V2C_3 (V2C_1139_179),
	.V2C_4 (V2C_1139_210),
	.V2C_5 (V2C_1139_219),
	.V2C_6 (V2C_1139_247),
	.V (V_1139)
);

VNU_6 #(quan_width) VNU1140 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_1140),
	.C2V_2 (C2V_128_1140),
	.C2V_3 (C2V_185_1140),
	.C2V_4 (C2V_216_1140),
	.C2V_5 (C2V_225_1140),
	.C2V_6 (C2V_253_1140),
	.L (L_1140),
	.V2C_1 (V2C_1140_52),
	.V2C_2 (V2C_1140_128),
	.V2C_3 (V2C_1140_185),
	.V2C_4 (V2C_1140_216),
	.V2C_5 (V2C_1140_225),
	.V2C_6 (V2C_1140_253),
	.V (V_1140)
);

VNU_6 #(quan_width) VNU1141 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_1141),
	.C2V_2 (C2V_134_1141),
	.C2V_3 (C2V_191_1141),
	.C2V_4 (C2V_222_1141),
	.C2V_5 (C2V_231_1141),
	.C2V_6 (C2V_259_1141),
	.L (L_1141),
	.V2C_1 (V2C_1141_58),
	.V2C_2 (V2C_1141_134),
	.V2C_3 (V2C_1141_191),
	.V2C_4 (V2C_1141_222),
	.V2C_5 (V2C_1141_231),
	.V2C_6 (V2C_1141_259),
	.V (V_1141)
);

VNU_6 #(quan_width) VNU1142 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_1142),
	.C2V_2 (C2V_140_1142),
	.C2V_3 (C2V_197_1142),
	.C2V_4 (C2V_228_1142),
	.C2V_5 (C2V_237_1142),
	.C2V_6 (C2V_265_1142),
	.L (L_1142),
	.V2C_1 (V2C_1142_64),
	.V2C_2 (V2C_1142_140),
	.V2C_3 (V2C_1142_197),
	.V2C_4 (V2C_1142_228),
	.V2C_5 (V2C_1142_237),
	.V2C_6 (V2C_1142_265),
	.V (V_1142)
);

VNU_6 #(quan_width) VNU1143 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_1143),
	.C2V_2 (C2V_146_1143),
	.C2V_3 (C2V_203_1143),
	.C2V_4 (C2V_234_1143),
	.C2V_5 (C2V_243_1143),
	.C2V_6 (C2V_271_1143),
	.L (L_1143),
	.V2C_1 (V2C_1143_70),
	.V2C_2 (V2C_1143_146),
	.V2C_3 (V2C_1143_203),
	.V2C_4 (V2C_1143_234),
	.V2C_5 (V2C_1143_243),
	.V2C_6 (V2C_1143_271),
	.V (V_1143)
);

VNU_6 #(quan_width) VNU1144 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_1144),
	.C2V_2 (C2V_152_1144),
	.C2V_3 (C2V_209_1144),
	.C2V_4 (C2V_240_1144),
	.C2V_5 (C2V_249_1144),
	.C2V_6 (C2V_277_1144),
	.L (L_1144),
	.V2C_1 (V2C_1144_76),
	.V2C_2 (V2C_1144_152),
	.V2C_3 (V2C_1144_209),
	.V2C_4 (V2C_1144_240),
	.V2C_5 (V2C_1144_249),
	.V2C_6 (V2C_1144_277),
	.V (V_1144)
);

VNU_6 #(quan_width) VNU1145 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_1145),
	.C2V_2 (C2V_158_1145),
	.C2V_3 (C2V_215_1145),
	.C2V_4 (C2V_246_1145),
	.C2V_5 (C2V_255_1145),
	.C2V_6 (C2V_283_1145),
	.L (L_1145),
	.V2C_1 (V2C_1145_82),
	.V2C_2 (V2C_1145_158),
	.V2C_3 (V2C_1145_215),
	.V2C_4 (V2C_1145_246),
	.V2C_5 (V2C_1145_255),
	.V2C_6 (V2C_1145_283),
	.V (V_1145)
);

VNU_6 #(quan_width) VNU1146 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_1146),
	.C2V_2 (C2V_88_1146),
	.C2V_3 (C2V_164_1146),
	.C2V_4 (C2V_221_1146),
	.C2V_5 (C2V_252_1146),
	.C2V_6 (C2V_261_1146),
	.L (L_1146),
	.V2C_1 (V2C_1146_1),
	.V2C_2 (V2C_1146_88),
	.V2C_3 (V2C_1146_164),
	.V2C_4 (V2C_1146_221),
	.V2C_5 (V2C_1146_252),
	.V2C_6 (V2C_1146_261),
	.V (V_1146)
);

VNU_6 #(quan_width) VNU1147 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_1147),
	.C2V_2 (C2V_94_1147),
	.C2V_3 (C2V_170_1147),
	.C2V_4 (C2V_227_1147),
	.C2V_5 (C2V_258_1147),
	.C2V_6 (C2V_267_1147),
	.L (L_1147),
	.V2C_1 (V2C_1147_7),
	.V2C_2 (V2C_1147_94),
	.V2C_3 (V2C_1147_170),
	.V2C_4 (V2C_1147_227),
	.V2C_5 (V2C_1147_258),
	.V2C_6 (V2C_1147_267),
	.V (V_1147)
);

VNU_6 #(quan_width) VNU1148 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_1148),
	.C2V_2 (C2V_100_1148),
	.C2V_3 (C2V_176_1148),
	.C2V_4 (C2V_233_1148),
	.C2V_5 (C2V_264_1148),
	.C2V_6 (C2V_273_1148),
	.L (L_1148),
	.V2C_1 (V2C_1148_13),
	.V2C_2 (V2C_1148_100),
	.V2C_3 (V2C_1148_176),
	.V2C_4 (V2C_1148_233),
	.V2C_5 (V2C_1148_264),
	.V2C_6 (V2C_1148_273),
	.V (V_1148)
);

VNU_6 #(quan_width) VNU1149 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_1149),
	.C2V_2 (C2V_106_1149),
	.C2V_3 (C2V_182_1149),
	.C2V_4 (C2V_239_1149),
	.C2V_5 (C2V_270_1149),
	.C2V_6 (C2V_279_1149),
	.L (L_1149),
	.V2C_1 (V2C_1149_19),
	.V2C_2 (V2C_1149_106),
	.V2C_3 (V2C_1149_182),
	.V2C_4 (V2C_1149_239),
	.V2C_5 (V2C_1149_270),
	.V2C_6 (V2C_1149_279),
	.V (V_1149)
);

VNU_6 #(quan_width) VNU1150 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_1150),
	.C2V_2 (C2V_112_1150),
	.C2V_3 (C2V_188_1150),
	.C2V_4 (C2V_245_1150),
	.C2V_5 (C2V_276_1150),
	.C2V_6 (C2V_285_1150),
	.L (L_1150),
	.V2C_1 (V2C_1150_25),
	.V2C_2 (V2C_1150_112),
	.V2C_3 (V2C_1150_188),
	.V2C_4 (V2C_1150_245),
	.V2C_5 (V2C_1150_276),
	.V2C_6 (V2C_1150_285),
	.V (V_1150)
);

VNU_6 #(quan_width) VNU1151 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_1151),
	.C2V_2 (C2V_31_1151),
	.C2V_3 (C2V_118_1151),
	.C2V_4 (C2V_194_1151),
	.C2V_5 (C2V_251_1151),
	.C2V_6 (C2V_282_1151),
	.L (L_1151),
	.V2C_1 (V2C_1151_3),
	.V2C_2 (V2C_1151_31),
	.V2C_3 (V2C_1151_118),
	.V2C_4 (V2C_1151_194),
	.V2C_5 (V2C_1151_251),
	.V2C_6 (V2C_1151_282),
	.V (V_1151)
);

VNU_6 #(quan_width) VNU1152 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_1152),
	.C2V_2 (C2V_37_1152),
	.C2V_3 (C2V_124_1152),
	.C2V_4 (C2V_200_1152),
	.C2V_5 (C2V_257_1152),
	.C2V_6 (C2V_288_1152),
	.L (L_1152),
	.V2C_1 (V2C_1152_9),
	.V2C_2 (V2C_1152_37),
	.V2C_3 (V2C_1152_124),
	.V2C_4 (V2C_1152_200),
	.V2C_5 (V2C_1152_257),
	.V2C_6 (V2C_1152_288),
	.V (V_1152)
);

VNU_2 #(quan_width) VNU1153 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_1_1153),
	.C2V_2 (C2V_2_1153),
	.L (L_1153),
	.V2C_1 (V2C_1153_1),
	.V2C_2 (V2C_1153_2),
	.V (V_1153)
);

VNU_2 #(quan_width) VNU1154 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_2_1154),
	.C2V_2 (C2V_3_1154),
	.L (L_1154),
	.V2C_1 (V2C_1154_2),
	.V2C_2 (V2C_1154_3),
	.V (V_1154)
);

VNU_2 #(quan_width) VNU1155 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_3_1155),
	.C2V_2 (C2V_4_1155),
	.L (L_1155),
	.V2C_1 (V2C_1155_3),
	.V2C_2 (V2C_1155_4),
	.V (V_1155)
);

VNU_2 #(quan_width) VNU1156 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_4_1156),
	.C2V_2 (C2V_5_1156),
	.L (L_1156),
	.V2C_1 (V2C_1156_4),
	.V2C_2 (V2C_1156_5),
	.V (V_1156)
);

VNU_2 #(quan_width) VNU1157 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_5_1157),
	.C2V_2 (C2V_6_1157),
	.L (L_1157),
	.V2C_1 (V2C_1157_5),
	.V2C_2 (V2C_1157_6),
	.V (V_1157)
);

VNU_2 #(quan_width) VNU1158 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_6_1158),
	.C2V_2 (C2V_7_1158),
	.L (L_1158),
	.V2C_1 (V2C_1158_6),
	.V2C_2 (V2C_1158_7),
	.V (V_1158)
);

VNU_2 #(quan_width) VNU1159 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_7_1159),
	.C2V_2 (C2V_8_1159),
	.L (L_1159),
	.V2C_1 (V2C_1159_7),
	.V2C_2 (V2C_1159_8),
	.V (V_1159)
);

VNU_2 #(quan_width) VNU1160 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_8_1160),
	.C2V_2 (C2V_9_1160),
	.L (L_1160),
	.V2C_1 (V2C_1160_8),
	.V2C_2 (V2C_1160_9),
	.V (V_1160)
);

VNU_2 #(quan_width) VNU1161 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_9_1161),
	.C2V_2 (C2V_10_1161),
	.L (L_1161),
	.V2C_1 (V2C_1161_9),
	.V2C_2 (V2C_1161_10),
	.V (V_1161)
);

VNU_2 #(quan_width) VNU1162 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_10_1162),
	.C2V_2 (C2V_11_1162),
	.L (L_1162),
	.V2C_1 (V2C_1162_10),
	.V2C_2 (V2C_1162_11),
	.V (V_1162)
);

VNU_2 #(quan_width) VNU1163 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_11_1163),
	.C2V_2 (C2V_12_1163),
	.L (L_1163),
	.V2C_1 (V2C_1163_11),
	.V2C_2 (V2C_1163_12),
	.V (V_1163)
);

VNU_2 #(quan_width) VNU1164 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_12_1164),
	.C2V_2 (C2V_13_1164),
	.L (L_1164),
	.V2C_1 (V2C_1164_12),
	.V2C_2 (V2C_1164_13),
	.V (V_1164)
);

VNU_2 #(quan_width) VNU1165 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_13_1165),
	.C2V_2 (C2V_14_1165),
	.L (L_1165),
	.V2C_1 (V2C_1165_13),
	.V2C_2 (V2C_1165_14),
	.V (V_1165)
);

VNU_2 #(quan_width) VNU1166 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_14_1166),
	.C2V_2 (C2V_15_1166),
	.L (L_1166),
	.V2C_1 (V2C_1166_14),
	.V2C_2 (V2C_1166_15),
	.V (V_1166)
);

VNU_2 #(quan_width) VNU1167 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_15_1167),
	.C2V_2 (C2V_16_1167),
	.L (L_1167),
	.V2C_1 (V2C_1167_15),
	.V2C_2 (V2C_1167_16),
	.V (V_1167)
);

VNU_2 #(quan_width) VNU1168 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_16_1168),
	.C2V_2 (C2V_17_1168),
	.L (L_1168),
	.V2C_1 (V2C_1168_16),
	.V2C_2 (V2C_1168_17),
	.V (V_1168)
);

VNU_2 #(quan_width) VNU1169 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_17_1169),
	.C2V_2 (C2V_18_1169),
	.L (L_1169),
	.V2C_1 (V2C_1169_17),
	.V2C_2 (V2C_1169_18),
	.V (V_1169)
);

VNU_2 #(quan_width) VNU1170 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_18_1170),
	.C2V_2 (C2V_19_1170),
	.L (L_1170),
	.V2C_1 (V2C_1170_18),
	.V2C_2 (V2C_1170_19),
	.V (V_1170)
);

VNU_2 #(quan_width) VNU1171 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_19_1171),
	.C2V_2 (C2V_20_1171),
	.L (L_1171),
	.V2C_1 (V2C_1171_19),
	.V2C_2 (V2C_1171_20),
	.V (V_1171)
);

VNU_2 #(quan_width) VNU1172 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_20_1172),
	.C2V_2 (C2V_21_1172),
	.L (L_1172),
	.V2C_1 (V2C_1172_20),
	.V2C_2 (V2C_1172_21),
	.V (V_1172)
);

VNU_2 #(quan_width) VNU1173 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_21_1173),
	.C2V_2 (C2V_22_1173),
	.L (L_1173),
	.V2C_1 (V2C_1173_21),
	.V2C_2 (V2C_1173_22),
	.V (V_1173)
);

VNU_2 #(quan_width) VNU1174 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_22_1174),
	.C2V_2 (C2V_23_1174),
	.L (L_1174),
	.V2C_1 (V2C_1174_22),
	.V2C_2 (V2C_1174_23),
	.V (V_1174)
);

VNU_2 #(quan_width) VNU1175 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_23_1175),
	.C2V_2 (C2V_24_1175),
	.L (L_1175),
	.V2C_1 (V2C_1175_23),
	.V2C_2 (V2C_1175_24),
	.V (V_1175)
);

VNU_2 #(quan_width) VNU1176 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_24_1176),
	.C2V_2 (C2V_25_1176),
	.L (L_1176),
	.V2C_1 (V2C_1176_24),
	.V2C_2 (V2C_1176_25),
	.V (V_1176)
);

VNU_2 #(quan_width) VNU1177 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_25_1177),
	.C2V_2 (C2V_26_1177),
	.L (L_1177),
	.V2C_1 (V2C_1177_25),
	.V2C_2 (V2C_1177_26),
	.V (V_1177)
);

VNU_2 #(quan_width) VNU1178 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_26_1178),
	.C2V_2 (C2V_27_1178),
	.L (L_1178),
	.V2C_1 (V2C_1178_26),
	.V2C_2 (V2C_1178_27),
	.V (V_1178)
);

VNU_2 #(quan_width) VNU1179 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_27_1179),
	.C2V_2 (C2V_28_1179),
	.L (L_1179),
	.V2C_1 (V2C_1179_27),
	.V2C_2 (V2C_1179_28),
	.V (V_1179)
);

VNU_2 #(quan_width) VNU1180 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_28_1180),
	.C2V_2 (C2V_29_1180),
	.L (L_1180),
	.V2C_1 (V2C_1180_28),
	.V2C_2 (V2C_1180_29),
	.V (V_1180)
);

VNU_2 #(quan_width) VNU1181 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_29_1181),
	.C2V_2 (C2V_30_1181),
	.L (L_1181),
	.V2C_1 (V2C_1181_29),
	.V2C_2 (V2C_1181_30),
	.V (V_1181)
);

VNU_2 #(quan_width) VNU1182 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_30_1182),
	.C2V_2 (C2V_31_1182),
	.L (L_1182),
	.V2C_1 (V2C_1182_30),
	.V2C_2 (V2C_1182_31),
	.V (V_1182)
);

VNU_2 #(quan_width) VNU1183 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_31_1183),
	.C2V_2 (C2V_32_1183),
	.L (L_1183),
	.V2C_1 (V2C_1183_31),
	.V2C_2 (V2C_1183_32),
	.V (V_1183)
);

VNU_2 #(quan_width) VNU1184 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_32_1184),
	.C2V_2 (C2V_33_1184),
	.L (L_1184),
	.V2C_1 (V2C_1184_32),
	.V2C_2 (V2C_1184_33),
	.V (V_1184)
);

VNU_2 #(quan_width) VNU1185 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_33_1185),
	.C2V_2 (C2V_34_1185),
	.L (L_1185),
	.V2C_1 (V2C_1185_33),
	.V2C_2 (V2C_1185_34),
	.V (V_1185)
);

VNU_2 #(quan_width) VNU1186 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_34_1186),
	.C2V_2 (C2V_35_1186),
	.L (L_1186),
	.V2C_1 (V2C_1186_34),
	.V2C_2 (V2C_1186_35),
	.V (V_1186)
);

VNU_2 #(quan_width) VNU1187 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_35_1187),
	.C2V_2 (C2V_36_1187),
	.L (L_1187),
	.V2C_1 (V2C_1187_35),
	.V2C_2 (V2C_1187_36),
	.V (V_1187)
);

VNU_2 #(quan_width) VNU1188 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_36_1188),
	.C2V_2 (C2V_37_1188),
	.L (L_1188),
	.V2C_1 (V2C_1188_36),
	.V2C_2 (V2C_1188_37),
	.V (V_1188)
);

VNU_2 #(quan_width) VNU1189 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_37_1189),
	.C2V_2 (C2V_38_1189),
	.L (L_1189),
	.V2C_1 (V2C_1189_37),
	.V2C_2 (V2C_1189_38),
	.V (V_1189)
);

VNU_2 #(quan_width) VNU1190 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_38_1190),
	.C2V_2 (C2V_39_1190),
	.L (L_1190),
	.V2C_1 (V2C_1190_38),
	.V2C_2 (V2C_1190_39),
	.V (V_1190)
);

VNU_2 #(quan_width) VNU1191 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_39_1191),
	.C2V_2 (C2V_40_1191),
	.L (L_1191),
	.V2C_1 (V2C_1191_39),
	.V2C_2 (V2C_1191_40),
	.V (V_1191)
);

VNU_2 #(quan_width) VNU1192 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_40_1192),
	.C2V_2 (C2V_41_1192),
	.L (L_1192),
	.V2C_1 (V2C_1192_40),
	.V2C_2 (V2C_1192_41),
	.V (V_1192)
);

VNU_2 #(quan_width) VNU1193 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_41_1193),
	.C2V_2 (C2V_42_1193),
	.L (L_1193),
	.V2C_1 (V2C_1193_41),
	.V2C_2 (V2C_1193_42),
	.V (V_1193)
);

VNU_2 #(quan_width) VNU1194 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_42_1194),
	.C2V_2 (C2V_43_1194),
	.L (L_1194),
	.V2C_1 (V2C_1194_42),
	.V2C_2 (V2C_1194_43),
	.V (V_1194)
);

VNU_2 #(quan_width) VNU1195 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_43_1195),
	.C2V_2 (C2V_44_1195),
	.L (L_1195),
	.V2C_1 (V2C_1195_43),
	.V2C_2 (V2C_1195_44),
	.V (V_1195)
);

VNU_2 #(quan_width) VNU1196 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_44_1196),
	.C2V_2 (C2V_45_1196),
	.L (L_1196),
	.V2C_1 (V2C_1196_44),
	.V2C_2 (V2C_1196_45),
	.V (V_1196)
);

VNU_2 #(quan_width) VNU1197 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_45_1197),
	.C2V_2 (C2V_46_1197),
	.L (L_1197),
	.V2C_1 (V2C_1197_45),
	.V2C_2 (V2C_1197_46),
	.V (V_1197)
);

VNU_2 #(quan_width) VNU1198 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_46_1198),
	.C2V_2 (C2V_47_1198),
	.L (L_1198),
	.V2C_1 (V2C_1198_46),
	.V2C_2 (V2C_1198_47),
	.V (V_1198)
);

VNU_2 #(quan_width) VNU1199 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_47_1199),
	.C2V_2 (C2V_48_1199),
	.L (L_1199),
	.V2C_1 (V2C_1199_47),
	.V2C_2 (V2C_1199_48),
	.V (V_1199)
);

VNU_2 #(quan_width) VNU1200 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_48_1200),
	.C2V_2 (C2V_49_1200),
	.L (L_1200),
	.V2C_1 (V2C_1200_48),
	.V2C_2 (V2C_1200_49),
	.V (V_1200)
);

VNU_2 #(quan_width) VNU1201 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_49_1201),
	.C2V_2 (C2V_50_1201),
	.L (L_1201),
	.V2C_1 (V2C_1201_49),
	.V2C_2 (V2C_1201_50),
	.V (V_1201)
);

VNU_2 #(quan_width) VNU1202 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_50_1202),
	.C2V_2 (C2V_51_1202),
	.L (L_1202),
	.V2C_1 (V2C_1202_50),
	.V2C_2 (V2C_1202_51),
	.V (V_1202)
);

VNU_2 #(quan_width) VNU1203 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_51_1203),
	.C2V_2 (C2V_52_1203),
	.L (L_1203),
	.V2C_1 (V2C_1203_51),
	.V2C_2 (V2C_1203_52),
	.V (V_1203)
);

VNU_2 #(quan_width) VNU1204 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_52_1204),
	.C2V_2 (C2V_53_1204),
	.L (L_1204),
	.V2C_1 (V2C_1204_52),
	.V2C_2 (V2C_1204_53),
	.V (V_1204)
);

VNU_2 #(quan_width) VNU1205 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_53_1205),
	.C2V_2 (C2V_54_1205),
	.L (L_1205),
	.V2C_1 (V2C_1205_53),
	.V2C_2 (V2C_1205_54),
	.V (V_1205)
);

VNU_2 #(quan_width) VNU1206 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_54_1206),
	.C2V_2 (C2V_55_1206),
	.L (L_1206),
	.V2C_1 (V2C_1206_54),
	.V2C_2 (V2C_1206_55),
	.V (V_1206)
);

VNU_2 #(quan_width) VNU1207 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_55_1207),
	.C2V_2 (C2V_56_1207),
	.L (L_1207),
	.V2C_1 (V2C_1207_55),
	.V2C_2 (V2C_1207_56),
	.V (V_1207)
);

VNU_2 #(quan_width) VNU1208 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_56_1208),
	.C2V_2 (C2V_57_1208),
	.L (L_1208),
	.V2C_1 (V2C_1208_56),
	.V2C_2 (V2C_1208_57),
	.V (V_1208)
);

VNU_2 #(quan_width) VNU1209 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_57_1209),
	.C2V_2 (C2V_58_1209),
	.L (L_1209),
	.V2C_1 (V2C_1209_57),
	.V2C_2 (V2C_1209_58),
	.V (V_1209)
);

VNU_2 #(quan_width) VNU1210 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_58_1210),
	.C2V_2 (C2V_59_1210),
	.L (L_1210),
	.V2C_1 (V2C_1210_58),
	.V2C_2 (V2C_1210_59),
	.V (V_1210)
);

VNU_2 #(quan_width) VNU1211 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_59_1211),
	.C2V_2 (C2V_60_1211),
	.L (L_1211),
	.V2C_1 (V2C_1211_59),
	.V2C_2 (V2C_1211_60),
	.V (V_1211)
);

VNU_2 #(quan_width) VNU1212 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_60_1212),
	.C2V_2 (C2V_61_1212),
	.L (L_1212),
	.V2C_1 (V2C_1212_60),
	.V2C_2 (V2C_1212_61),
	.V (V_1212)
);

VNU_2 #(quan_width) VNU1213 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_61_1213),
	.C2V_2 (C2V_62_1213),
	.L (L_1213),
	.V2C_1 (V2C_1213_61),
	.V2C_2 (V2C_1213_62),
	.V (V_1213)
);

VNU_2 #(quan_width) VNU1214 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_62_1214),
	.C2V_2 (C2V_63_1214),
	.L (L_1214),
	.V2C_1 (V2C_1214_62),
	.V2C_2 (V2C_1214_63),
	.V (V_1214)
);

VNU_2 #(quan_width) VNU1215 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_63_1215),
	.C2V_2 (C2V_64_1215),
	.L (L_1215),
	.V2C_1 (V2C_1215_63),
	.V2C_2 (V2C_1215_64),
	.V (V_1215)
);

VNU_2 #(quan_width) VNU1216 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_64_1216),
	.C2V_2 (C2V_65_1216),
	.L (L_1216),
	.V2C_1 (V2C_1216_64),
	.V2C_2 (V2C_1216_65),
	.V (V_1216)
);

VNU_2 #(quan_width) VNU1217 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_65_1217),
	.C2V_2 (C2V_66_1217),
	.L (L_1217),
	.V2C_1 (V2C_1217_65),
	.V2C_2 (V2C_1217_66),
	.V (V_1217)
);

VNU_2 #(quan_width) VNU1218 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_66_1218),
	.C2V_2 (C2V_67_1218),
	.L (L_1218),
	.V2C_1 (V2C_1218_66),
	.V2C_2 (V2C_1218_67),
	.V (V_1218)
);

VNU_2 #(quan_width) VNU1219 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_67_1219),
	.C2V_2 (C2V_68_1219),
	.L (L_1219),
	.V2C_1 (V2C_1219_67),
	.V2C_2 (V2C_1219_68),
	.V (V_1219)
);

VNU_2 #(quan_width) VNU1220 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_68_1220),
	.C2V_2 (C2V_69_1220),
	.L (L_1220),
	.V2C_1 (V2C_1220_68),
	.V2C_2 (V2C_1220_69),
	.V (V_1220)
);

VNU_2 #(quan_width) VNU1221 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_69_1221),
	.C2V_2 (C2V_70_1221),
	.L (L_1221),
	.V2C_1 (V2C_1221_69),
	.V2C_2 (V2C_1221_70),
	.V (V_1221)
);

VNU_2 #(quan_width) VNU1222 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_70_1222),
	.C2V_2 (C2V_71_1222),
	.L (L_1222),
	.V2C_1 (V2C_1222_70),
	.V2C_2 (V2C_1222_71),
	.V (V_1222)
);

VNU_2 #(quan_width) VNU1223 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_71_1223),
	.C2V_2 (C2V_72_1223),
	.L (L_1223),
	.V2C_1 (V2C_1223_71),
	.V2C_2 (V2C_1223_72),
	.V (V_1223)
);

VNU_2 #(quan_width) VNU1224 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_72_1224),
	.C2V_2 (C2V_73_1224),
	.L (L_1224),
	.V2C_1 (V2C_1224_72),
	.V2C_2 (V2C_1224_73),
	.V (V_1224)
);

VNU_2 #(quan_width) VNU1225 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_73_1225),
	.C2V_2 (C2V_74_1225),
	.L (L_1225),
	.V2C_1 (V2C_1225_73),
	.V2C_2 (V2C_1225_74),
	.V (V_1225)
);

VNU_2 #(quan_width) VNU1226 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_74_1226),
	.C2V_2 (C2V_75_1226),
	.L (L_1226),
	.V2C_1 (V2C_1226_74),
	.V2C_2 (V2C_1226_75),
	.V (V_1226)
);

VNU_2 #(quan_width) VNU1227 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_75_1227),
	.C2V_2 (C2V_76_1227),
	.L (L_1227),
	.V2C_1 (V2C_1227_75),
	.V2C_2 (V2C_1227_76),
	.V (V_1227)
);

VNU_2 #(quan_width) VNU1228 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_76_1228),
	.C2V_2 (C2V_77_1228),
	.L (L_1228),
	.V2C_1 (V2C_1228_76),
	.V2C_2 (V2C_1228_77),
	.V (V_1228)
);

VNU_2 #(quan_width) VNU1229 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_77_1229),
	.C2V_2 (C2V_78_1229),
	.L (L_1229),
	.V2C_1 (V2C_1229_77),
	.V2C_2 (V2C_1229_78),
	.V (V_1229)
);

VNU_2 #(quan_width) VNU1230 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_78_1230),
	.C2V_2 (C2V_79_1230),
	.L (L_1230),
	.V2C_1 (V2C_1230_78),
	.V2C_2 (V2C_1230_79),
	.V (V_1230)
);

VNU_2 #(quan_width) VNU1231 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_79_1231),
	.C2V_2 (C2V_80_1231),
	.L (L_1231),
	.V2C_1 (V2C_1231_79),
	.V2C_2 (V2C_1231_80),
	.V (V_1231)
);

VNU_2 #(quan_width) VNU1232 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_80_1232),
	.C2V_2 (C2V_81_1232),
	.L (L_1232),
	.V2C_1 (V2C_1232_80),
	.V2C_2 (V2C_1232_81),
	.V (V_1232)
);

VNU_2 #(quan_width) VNU1233 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_81_1233),
	.C2V_2 (C2V_82_1233),
	.L (L_1233),
	.V2C_1 (V2C_1233_81),
	.V2C_2 (V2C_1233_82),
	.V (V_1233)
);

VNU_2 #(quan_width) VNU1234 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_82_1234),
	.C2V_2 (C2V_83_1234),
	.L (L_1234),
	.V2C_1 (V2C_1234_82),
	.V2C_2 (V2C_1234_83),
	.V (V_1234)
);

VNU_2 #(quan_width) VNU1235 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_83_1235),
	.C2V_2 (C2V_84_1235),
	.L (L_1235),
	.V2C_1 (V2C_1235_83),
	.V2C_2 (V2C_1235_84),
	.V (V_1235)
);

VNU_2 #(quan_width) VNU1236 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_84_1236),
	.C2V_2 (C2V_85_1236),
	.L (L_1236),
	.V2C_1 (V2C_1236_84),
	.V2C_2 (V2C_1236_85),
	.V (V_1236)
);

VNU_2 #(quan_width) VNU1237 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_85_1237),
	.C2V_2 (C2V_86_1237),
	.L (L_1237),
	.V2C_1 (V2C_1237_85),
	.V2C_2 (V2C_1237_86),
	.V (V_1237)
);

VNU_2 #(quan_width) VNU1238 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_86_1238),
	.C2V_2 (C2V_87_1238),
	.L (L_1238),
	.V2C_1 (V2C_1238_86),
	.V2C_2 (V2C_1238_87),
	.V (V_1238)
);

VNU_2 #(quan_width) VNU1239 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_87_1239),
	.C2V_2 (C2V_88_1239),
	.L (L_1239),
	.V2C_1 (V2C_1239_87),
	.V2C_2 (V2C_1239_88),
	.V (V_1239)
);

VNU_2 #(quan_width) VNU1240 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_88_1240),
	.C2V_2 (C2V_89_1240),
	.L (L_1240),
	.V2C_1 (V2C_1240_88),
	.V2C_2 (V2C_1240_89),
	.V (V_1240)
);

VNU_2 #(quan_width) VNU1241 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_89_1241),
	.C2V_2 (C2V_90_1241),
	.L (L_1241),
	.V2C_1 (V2C_1241_89),
	.V2C_2 (V2C_1241_90),
	.V (V_1241)
);

VNU_2 #(quan_width) VNU1242 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_90_1242),
	.C2V_2 (C2V_91_1242),
	.L (L_1242),
	.V2C_1 (V2C_1242_90),
	.V2C_2 (V2C_1242_91),
	.V (V_1242)
);

VNU_2 #(quan_width) VNU1243 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_91_1243),
	.C2V_2 (C2V_92_1243),
	.L (L_1243),
	.V2C_1 (V2C_1243_91),
	.V2C_2 (V2C_1243_92),
	.V (V_1243)
);

VNU_2 #(quan_width) VNU1244 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_92_1244),
	.C2V_2 (C2V_93_1244),
	.L (L_1244),
	.V2C_1 (V2C_1244_92),
	.V2C_2 (V2C_1244_93),
	.V (V_1244)
);

VNU_2 #(quan_width) VNU1245 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_93_1245),
	.C2V_2 (C2V_94_1245),
	.L (L_1245),
	.V2C_1 (V2C_1245_93),
	.V2C_2 (V2C_1245_94),
	.V (V_1245)
);

VNU_2 #(quan_width) VNU1246 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_94_1246),
	.C2V_2 (C2V_95_1246),
	.L (L_1246),
	.V2C_1 (V2C_1246_94),
	.V2C_2 (V2C_1246_95),
	.V (V_1246)
);

VNU_2 #(quan_width) VNU1247 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_95_1247),
	.C2V_2 (C2V_96_1247),
	.L (L_1247),
	.V2C_1 (V2C_1247_95),
	.V2C_2 (V2C_1247_96),
	.V (V_1247)
);

VNU_2 #(quan_width) VNU1248 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_96_1248),
	.C2V_2 (C2V_97_1248),
	.L (L_1248),
	.V2C_1 (V2C_1248_96),
	.V2C_2 (V2C_1248_97),
	.V (V_1248)
);

VNU_2 #(quan_width) VNU1249 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_97_1249),
	.C2V_2 (C2V_98_1249),
	.L (L_1249),
	.V2C_1 (V2C_1249_97),
	.V2C_2 (V2C_1249_98),
	.V (V_1249)
);

VNU_2 #(quan_width) VNU1250 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_98_1250),
	.C2V_2 (C2V_99_1250),
	.L (L_1250),
	.V2C_1 (V2C_1250_98),
	.V2C_2 (V2C_1250_99),
	.V (V_1250)
);

VNU_2 #(quan_width) VNU1251 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_99_1251),
	.C2V_2 (C2V_100_1251),
	.L (L_1251),
	.V2C_1 (V2C_1251_99),
	.V2C_2 (V2C_1251_100),
	.V (V_1251)
);

VNU_2 #(quan_width) VNU1252 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_100_1252),
	.C2V_2 (C2V_101_1252),
	.L (L_1252),
	.V2C_1 (V2C_1252_100),
	.V2C_2 (V2C_1252_101),
	.V (V_1252)
);

VNU_2 #(quan_width) VNU1253 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_101_1253),
	.C2V_2 (C2V_102_1253),
	.L (L_1253),
	.V2C_1 (V2C_1253_101),
	.V2C_2 (V2C_1253_102),
	.V (V_1253)
);

VNU_2 #(quan_width) VNU1254 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_102_1254),
	.C2V_2 (C2V_103_1254),
	.L (L_1254),
	.V2C_1 (V2C_1254_102),
	.V2C_2 (V2C_1254_103),
	.V (V_1254)
);

VNU_2 #(quan_width) VNU1255 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_103_1255),
	.C2V_2 (C2V_104_1255),
	.L (L_1255),
	.V2C_1 (V2C_1255_103),
	.V2C_2 (V2C_1255_104),
	.V (V_1255)
);

VNU_2 #(quan_width) VNU1256 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_104_1256),
	.C2V_2 (C2V_105_1256),
	.L (L_1256),
	.V2C_1 (V2C_1256_104),
	.V2C_2 (V2C_1256_105),
	.V (V_1256)
);

VNU_2 #(quan_width) VNU1257 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_105_1257),
	.C2V_2 (C2V_106_1257),
	.L (L_1257),
	.V2C_1 (V2C_1257_105),
	.V2C_2 (V2C_1257_106),
	.V (V_1257)
);

VNU_2 #(quan_width) VNU1258 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_106_1258),
	.C2V_2 (C2V_107_1258),
	.L (L_1258),
	.V2C_1 (V2C_1258_106),
	.V2C_2 (V2C_1258_107),
	.V (V_1258)
);

VNU_2 #(quan_width) VNU1259 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_107_1259),
	.C2V_2 (C2V_108_1259),
	.L (L_1259),
	.V2C_1 (V2C_1259_107),
	.V2C_2 (V2C_1259_108),
	.V (V_1259)
);

VNU_2 #(quan_width) VNU1260 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_108_1260),
	.C2V_2 (C2V_109_1260),
	.L (L_1260),
	.V2C_1 (V2C_1260_108),
	.V2C_2 (V2C_1260_109),
	.V (V_1260)
);

VNU_2 #(quan_width) VNU1261 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_109_1261),
	.C2V_2 (C2V_110_1261),
	.L (L_1261),
	.V2C_1 (V2C_1261_109),
	.V2C_2 (V2C_1261_110),
	.V (V_1261)
);

VNU_2 #(quan_width) VNU1262 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_110_1262),
	.C2V_2 (C2V_111_1262),
	.L (L_1262),
	.V2C_1 (V2C_1262_110),
	.V2C_2 (V2C_1262_111),
	.V (V_1262)
);

VNU_2 #(quan_width) VNU1263 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_111_1263),
	.C2V_2 (C2V_112_1263),
	.L (L_1263),
	.V2C_1 (V2C_1263_111),
	.V2C_2 (V2C_1263_112),
	.V (V_1263)
);

VNU_2 #(quan_width) VNU1264 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_112_1264),
	.C2V_2 (C2V_113_1264),
	.L (L_1264),
	.V2C_1 (V2C_1264_112),
	.V2C_2 (V2C_1264_113),
	.V (V_1264)
);

VNU_2 #(quan_width) VNU1265 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_113_1265),
	.C2V_2 (C2V_114_1265),
	.L (L_1265),
	.V2C_1 (V2C_1265_113),
	.V2C_2 (V2C_1265_114),
	.V (V_1265)
);

VNU_2 #(quan_width) VNU1266 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_114_1266),
	.C2V_2 (C2V_115_1266),
	.L (L_1266),
	.V2C_1 (V2C_1266_114),
	.V2C_2 (V2C_1266_115),
	.V (V_1266)
);

VNU_2 #(quan_width) VNU1267 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_115_1267),
	.C2V_2 (C2V_116_1267),
	.L (L_1267),
	.V2C_1 (V2C_1267_115),
	.V2C_2 (V2C_1267_116),
	.V (V_1267)
);

VNU_2 #(quan_width) VNU1268 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_116_1268),
	.C2V_2 (C2V_117_1268),
	.L (L_1268),
	.V2C_1 (V2C_1268_116),
	.V2C_2 (V2C_1268_117),
	.V (V_1268)
);

VNU_2 #(quan_width) VNU1269 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_117_1269),
	.C2V_2 (C2V_118_1269),
	.L (L_1269),
	.V2C_1 (V2C_1269_117),
	.V2C_2 (V2C_1269_118),
	.V (V_1269)
);

VNU_2 #(quan_width) VNU1270 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_118_1270),
	.C2V_2 (C2V_119_1270),
	.L (L_1270),
	.V2C_1 (V2C_1270_118),
	.V2C_2 (V2C_1270_119),
	.V (V_1270)
);

VNU_2 #(quan_width) VNU1271 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_119_1271),
	.C2V_2 (C2V_120_1271),
	.L (L_1271),
	.V2C_1 (V2C_1271_119),
	.V2C_2 (V2C_1271_120),
	.V (V_1271)
);

VNU_2 #(quan_width) VNU1272 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_120_1272),
	.C2V_2 (C2V_121_1272),
	.L (L_1272),
	.V2C_1 (V2C_1272_120),
	.V2C_2 (V2C_1272_121),
	.V (V_1272)
);

VNU_2 #(quan_width) VNU1273 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_121_1273),
	.C2V_2 (C2V_122_1273),
	.L (L_1273),
	.V2C_1 (V2C_1273_121),
	.V2C_2 (V2C_1273_122),
	.V (V_1273)
);

VNU_2 #(quan_width) VNU1274 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_122_1274),
	.C2V_2 (C2V_123_1274),
	.L (L_1274),
	.V2C_1 (V2C_1274_122),
	.V2C_2 (V2C_1274_123),
	.V (V_1274)
);

VNU_2 #(quan_width) VNU1275 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_123_1275),
	.C2V_2 (C2V_124_1275),
	.L (L_1275),
	.V2C_1 (V2C_1275_123),
	.V2C_2 (V2C_1275_124),
	.V (V_1275)
);

VNU_2 #(quan_width) VNU1276 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_124_1276),
	.C2V_2 (C2V_125_1276),
	.L (L_1276),
	.V2C_1 (V2C_1276_124),
	.V2C_2 (V2C_1276_125),
	.V (V_1276)
);

VNU_2 #(quan_width) VNU1277 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_125_1277),
	.C2V_2 (C2V_126_1277),
	.L (L_1277),
	.V2C_1 (V2C_1277_125),
	.V2C_2 (V2C_1277_126),
	.V (V_1277)
);

VNU_2 #(quan_width) VNU1278 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_126_1278),
	.C2V_2 (C2V_127_1278),
	.L (L_1278),
	.V2C_1 (V2C_1278_126),
	.V2C_2 (V2C_1278_127),
	.V (V_1278)
);

VNU_2 #(quan_width) VNU1279 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_127_1279),
	.C2V_2 (C2V_128_1279),
	.L (L_1279),
	.V2C_1 (V2C_1279_127),
	.V2C_2 (V2C_1279_128),
	.V (V_1279)
);

VNU_2 #(quan_width) VNU1280 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_128_1280),
	.C2V_2 (C2V_129_1280),
	.L (L_1280),
	.V2C_1 (V2C_1280_128),
	.V2C_2 (V2C_1280_129),
	.V (V_1280)
);

VNU_2 #(quan_width) VNU1281 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_129_1281),
	.C2V_2 (C2V_130_1281),
	.L (L_1281),
	.V2C_1 (V2C_1281_129),
	.V2C_2 (V2C_1281_130),
	.V (V_1281)
);

VNU_2 #(quan_width) VNU1282 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_130_1282),
	.C2V_2 (C2V_131_1282),
	.L (L_1282),
	.V2C_1 (V2C_1282_130),
	.V2C_2 (V2C_1282_131),
	.V (V_1282)
);

VNU_2 #(quan_width) VNU1283 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_131_1283),
	.C2V_2 (C2V_132_1283),
	.L (L_1283),
	.V2C_1 (V2C_1283_131),
	.V2C_2 (V2C_1283_132),
	.V (V_1283)
);

VNU_2 #(quan_width) VNU1284 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_132_1284),
	.C2V_2 (C2V_133_1284),
	.L (L_1284),
	.V2C_1 (V2C_1284_132),
	.V2C_2 (V2C_1284_133),
	.V (V_1284)
);

VNU_2 #(quan_width) VNU1285 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_133_1285),
	.C2V_2 (C2V_134_1285),
	.L (L_1285),
	.V2C_1 (V2C_1285_133),
	.V2C_2 (V2C_1285_134),
	.V (V_1285)
);

VNU_2 #(quan_width) VNU1286 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_134_1286),
	.C2V_2 (C2V_135_1286),
	.L (L_1286),
	.V2C_1 (V2C_1286_134),
	.V2C_2 (V2C_1286_135),
	.V (V_1286)
);

VNU_2 #(quan_width) VNU1287 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_135_1287),
	.C2V_2 (C2V_136_1287),
	.L (L_1287),
	.V2C_1 (V2C_1287_135),
	.V2C_2 (V2C_1287_136),
	.V (V_1287)
);

VNU_2 #(quan_width) VNU1288 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_136_1288),
	.C2V_2 (C2V_137_1288),
	.L (L_1288),
	.V2C_1 (V2C_1288_136),
	.V2C_2 (V2C_1288_137),
	.V (V_1288)
);

VNU_2 #(quan_width) VNU1289 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_137_1289),
	.C2V_2 (C2V_138_1289),
	.L (L_1289),
	.V2C_1 (V2C_1289_137),
	.V2C_2 (V2C_1289_138),
	.V (V_1289)
);

VNU_2 #(quan_width) VNU1290 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_138_1290),
	.C2V_2 (C2V_139_1290),
	.L (L_1290),
	.V2C_1 (V2C_1290_138),
	.V2C_2 (V2C_1290_139),
	.V (V_1290)
);

VNU_2 #(quan_width) VNU1291 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_139_1291),
	.C2V_2 (C2V_140_1291),
	.L (L_1291),
	.V2C_1 (V2C_1291_139),
	.V2C_2 (V2C_1291_140),
	.V (V_1291)
);

VNU_2 #(quan_width) VNU1292 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_140_1292),
	.C2V_2 (C2V_141_1292),
	.L (L_1292),
	.V2C_1 (V2C_1292_140),
	.V2C_2 (V2C_1292_141),
	.V (V_1292)
);

VNU_2 #(quan_width) VNU1293 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_141_1293),
	.C2V_2 (C2V_142_1293),
	.L (L_1293),
	.V2C_1 (V2C_1293_141),
	.V2C_2 (V2C_1293_142),
	.V (V_1293)
);

VNU_2 #(quan_width) VNU1294 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_142_1294),
	.C2V_2 (C2V_143_1294),
	.L (L_1294),
	.V2C_1 (V2C_1294_142),
	.V2C_2 (V2C_1294_143),
	.V (V_1294)
);

VNU_2 #(quan_width) VNU1295 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_143_1295),
	.C2V_2 (C2V_144_1295),
	.L (L_1295),
	.V2C_1 (V2C_1295_143),
	.V2C_2 (V2C_1295_144),
	.V (V_1295)
);

VNU_2 #(quan_width) VNU1296 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_144_1296),
	.C2V_2 (C2V_145_1296),
	.L (L_1296),
	.V2C_1 (V2C_1296_144),
	.V2C_2 (V2C_1296_145),
	.V (V_1296)
);

VNU_2 #(quan_width) VNU1297 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_145_1297),
	.C2V_2 (C2V_146_1297),
	.L (L_1297),
	.V2C_1 (V2C_1297_145),
	.V2C_2 (V2C_1297_146),
	.V (V_1297)
);

VNU_2 #(quan_width) VNU1298 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_146_1298),
	.C2V_2 (C2V_147_1298),
	.L (L_1298),
	.V2C_1 (V2C_1298_146),
	.V2C_2 (V2C_1298_147),
	.V (V_1298)
);

VNU_2 #(quan_width) VNU1299 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_147_1299),
	.C2V_2 (C2V_148_1299),
	.L (L_1299),
	.V2C_1 (V2C_1299_147),
	.V2C_2 (V2C_1299_148),
	.V (V_1299)
);

VNU_2 #(quan_width) VNU1300 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_148_1300),
	.C2V_2 (C2V_149_1300),
	.L (L_1300),
	.V2C_1 (V2C_1300_148),
	.V2C_2 (V2C_1300_149),
	.V (V_1300)
);

VNU_2 #(quan_width) VNU1301 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_149_1301),
	.C2V_2 (C2V_150_1301),
	.L (L_1301),
	.V2C_1 (V2C_1301_149),
	.V2C_2 (V2C_1301_150),
	.V (V_1301)
);

VNU_2 #(quan_width) VNU1302 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_150_1302),
	.C2V_2 (C2V_151_1302),
	.L (L_1302),
	.V2C_1 (V2C_1302_150),
	.V2C_2 (V2C_1302_151),
	.V (V_1302)
);

VNU_2 #(quan_width) VNU1303 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_151_1303),
	.C2V_2 (C2V_152_1303),
	.L (L_1303),
	.V2C_1 (V2C_1303_151),
	.V2C_2 (V2C_1303_152),
	.V (V_1303)
);

VNU_2 #(quan_width) VNU1304 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_152_1304),
	.C2V_2 (C2V_153_1304),
	.L (L_1304),
	.V2C_1 (V2C_1304_152),
	.V2C_2 (V2C_1304_153),
	.V (V_1304)
);

VNU_2 #(quan_width) VNU1305 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_153_1305),
	.C2V_2 (C2V_154_1305),
	.L (L_1305),
	.V2C_1 (V2C_1305_153),
	.V2C_2 (V2C_1305_154),
	.V (V_1305)
);

VNU_2 #(quan_width) VNU1306 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_154_1306),
	.C2V_2 (C2V_155_1306),
	.L (L_1306),
	.V2C_1 (V2C_1306_154),
	.V2C_2 (V2C_1306_155),
	.V (V_1306)
);

VNU_2 #(quan_width) VNU1307 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_155_1307),
	.C2V_2 (C2V_156_1307),
	.L (L_1307),
	.V2C_1 (V2C_1307_155),
	.V2C_2 (V2C_1307_156),
	.V (V_1307)
);

VNU_2 #(quan_width) VNU1308 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_156_1308),
	.C2V_2 (C2V_157_1308),
	.L (L_1308),
	.V2C_1 (V2C_1308_156),
	.V2C_2 (V2C_1308_157),
	.V (V_1308)
);

VNU_2 #(quan_width) VNU1309 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_157_1309),
	.C2V_2 (C2V_158_1309),
	.L (L_1309),
	.V2C_1 (V2C_1309_157),
	.V2C_2 (V2C_1309_158),
	.V (V_1309)
);

VNU_2 #(quan_width) VNU1310 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_158_1310),
	.C2V_2 (C2V_159_1310),
	.L (L_1310),
	.V2C_1 (V2C_1310_158),
	.V2C_2 (V2C_1310_159),
	.V (V_1310)
);

VNU_2 #(quan_width) VNU1311 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_159_1311),
	.C2V_2 (C2V_160_1311),
	.L (L_1311),
	.V2C_1 (V2C_1311_159),
	.V2C_2 (V2C_1311_160),
	.V (V_1311)
);

VNU_2 #(quan_width) VNU1312 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_160_1312),
	.C2V_2 (C2V_161_1312),
	.L (L_1312),
	.V2C_1 (V2C_1312_160),
	.V2C_2 (V2C_1312_161),
	.V (V_1312)
);

VNU_2 #(quan_width) VNU1313 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_161_1313),
	.C2V_2 (C2V_162_1313),
	.L (L_1313),
	.V2C_1 (V2C_1313_161),
	.V2C_2 (V2C_1313_162),
	.V (V_1313)
);

VNU_2 #(quan_width) VNU1314 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_162_1314),
	.C2V_2 (C2V_163_1314),
	.L (L_1314),
	.V2C_1 (V2C_1314_162),
	.V2C_2 (V2C_1314_163),
	.V (V_1314)
);

VNU_2 #(quan_width) VNU1315 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_163_1315),
	.C2V_2 (C2V_164_1315),
	.L (L_1315),
	.V2C_1 (V2C_1315_163),
	.V2C_2 (V2C_1315_164),
	.V (V_1315)
);

VNU_2 #(quan_width) VNU1316 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_164_1316),
	.C2V_2 (C2V_165_1316),
	.L (L_1316),
	.V2C_1 (V2C_1316_164),
	.V2C_2 (V2C_1316_165),
	.V (V_1316)
);

VNU_2 #(quan_width) VNU1317 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_165_1317),
	.C2V_2 (C2V_166_1317),
	.L (L_1317),
	.V2C_1 (V2C_1317_165),
	.V2C_2 (V2C_1317_166),
	.V (V_1317)
);

VNU_2 #(quan_width) VNU1318 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_166_1318),
	.C2V_2 (C2V_167_1318),
	.L (L_1318),
	.V2C_1 (V2C_1318_166),
	.V2C_2 (V2C_1318_167),
	.V (V_1318)
);

VNU_2 #(quan_width) VNU1319 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_167_1319),
	.C2V_2 (C2V_168_1319),
	.L (L_1319),
	.V2C_1 (V2C_1319_167),
	.V2C_2 (V2C_1319_168),
	.V (V_1319)
);

VNU_2 #(quan_width) VNU1320 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_168_1320),
	.C2V_2 (C2V_169_1320),
	.L (L_1320),
	.V2C_1 (V2C_1320_168),
	.V2C_2 (V2C_1320_169),
	.V (V_1320)
);

VNU_2 #(quan_width) VNU1321 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_169_1321),
	.C2V_2 (C2V_170_1321),
	.L (L_1321),
	.V2C_1 (V2C_1321_169),
	.V2C_2 (V2C_1321_170),
	.V (V_1321)
);

VNU_2 #(quan_width) VNU1322 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_170_1322),
	.C2V_2 (C2V_171_1322),
	.L (L_1322),
	.V2C_1 (V2C_1322_170),
	.V2C_2 (V2C_1322_171),
	.V (V_1322)
);

VNU_2 #(quan_width) VNU1323 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_171_1323),
	.C2V_2 (C2V_172_1323),
	.L (L_1323),
	.V2C_1 (V2C_1323_171),
	.V2C_2 (V2C_1323_172),
	.V (V_1323)
);

VNU_2 #(quan_width) VNU1324 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_172_1324),
	.C2V_2 (C2V_173_1324),
	.L (L_1324),
	.V2C_1 (V2C_1324_172),
	.V2C_2 (V2C_1324_173),
	.V (V_1324)
);

VNU_2 #(quan_width) VNU1325 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_173_1325),
	.C2V_2 (C2V_174_1325),
	.L (L_1325),
	.V2C_1 (V2C_1325_173),
	.V2C_2 (V2C_1325_174),
	.V (V_1325)
);

VNU_2 #(quan_width) VNU1326 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_174_1326),
	.C2V_2 (C2V_175_1326),
	.L (L_1326),
	.V2C_1 (V2C_1326_174),
	.V2C_2 (V2C_1326_175),
	.V (V_1326)
);

VNU_2 #(quan_width) VNU1327 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_175_1327),
	.C2V_2 (C2V_176_1327),
	.L (L_1327),
	.V2C_1 (V2C_1327_175),
	.V2C_2 (V2C_1327_176),
	.V (V_1327)
);

VNU_2 #(quan_width) VNU1328 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_176_1328),
	.C2V_2 (C2V_177_1328),
	.L (L_1328),
	.V2C_1 (V2C_1328_176),
	.V2C_2 (V2C_1328_177),
	.V (V_1328)
);

VNU_2 #(quan_width) VNU1329 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_177_1329),
	.C2V_2 (C2V_178_1329),
	.L (L_1329),
	.V2C_1 (V2C_1329_177),
	.V2C_2 (V2C_1329_178),
	.V (V_1329)
);

VNU_2 #(quan_width) VNU1330 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_178_1330),
	.C2V_2 (C2V_179_1330),
	.L (L_1330),
	.V2C_1 (V2C_1330_178),
	.V2C_2 (V2C_1330_179),
	.V (V_1330)
);

VNU_2 #(quan_width) VNU1331 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_179_1331),
	.C2V_2 (C2V_180_1331),
	.L (L_1331),
	.V2C_1 (V2C_1331_179),
	.V2C_2 (V2C_1331_180),
	.V (V_1331)
);

VNU_2 #(quan_width) VNU1332 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_180_1332),
	.C2V_2 (C2V_181_1332),
	.L (L_1332),
	.V2C_1 (V2C_1332_180),
	.V2C_2 (V2C_1332_181),
	.V (V_1332)
);

VNU_2 #(quan_width) VNU1333 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_181_1333),
	.C2V_2 (C2V_182_1333),
	.L (L_1333),
	.V2C_1 (V2C_1333_181),
	.V2C_2 (V2C_1333_182),
	.V (V_1333)
);

VNU_2 #(quan_width) VNU1334 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_182_1334),
	.C2V_2 (C2V_183_1334),
	.L (L_1334),
	.V2C_1 (V2C_1334_182),
	.V2C_2 (V2C_1334_183),
	.V (V_1334)
);

VNU_2 #(quan_width) VNU1335 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_183_1335),
	.C2V_2 (C2V_184_1335),
	.L (L_1335),
	.V2C_1 (V2C_1335_183),
	.V2C_2 (V2C_1335_184),
	.V (V_1335)
);

VNU_2 #(quan_width) VNU1336 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_184_1336),
	.C2V_2 (C2V_185_1336),
	.L (L_1336),
	.V2C_1 (V2C_1336_184),
	.V2C_2 (V2C_1336_185),
	.V (V_1336)
);

VNU_2 #(quan_width) VNU1337 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_185_1337),
	.C2V_2 (C2V_186_1337),
	.L (L_1337),
	.V2C_1 (V2C_1337_185),
	.V2C_2 (V2C_1337_186),
	.V (V_1337)
);

VNU_2 #(quan_width) VNU1338 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_186_1338),
	.C2V_2 (C2V_187_1338),
	.L (L_1338),
	.V2C_1 (V2C_1338_186),
	.V2C_2 (V2C_1338_187),
	.V (V_1338)
);

VNU_2 #(quan_width) VNU1339 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_187_1339),
	.C2V_2 (C2V_188_1339),
	.L (L_1339),
	.V2C_1 (V2C_1339_187),
	.V2C_2 (V2C_1339_188),
	.V (V_1339)
);

VNU_2 #(quan_width) VNU1340 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_188_1340),
	.C2V_2 (C2V_189_1340),
	.L (L_1340),
	.V2C_1 (V2C_1340_188),
	.V2C_2 (V2C_1340_189),
	.V (V_1340)
);

VNU_2 #(quan_width) VNU1341 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_189_1341),
	.C2V_2 (C2V_190_1341),
	.L (L_1341),
	.V2C_1 (V2C_1341_189),
	.V2C_2 (V2C_1341_190),
	.V (V_1341)
);

VNU_2 #(quan_width) VNU1342 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_190_1342),
	.C2V_2 (C2V_191_1342),
	.L (L_1342),
	.V2C_1 (V2C_1342_190),
	.V2C_2 (V2C_1342_191),
	.V (V_1342)
);

VNU_2 #(quan_width) VNU1343 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_191_1343),
	.C2V_2 (C2V_192_1343),
	.L (L_1343),
	.V2C_1 (V2C_1343_191),
	.V2C_2 (V2C_1343_192),
	.V (V_1343)
);

VNU_2 #(quan_width) VNU1344 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_192_1344),
	.C2V_2 (C2V_193_1344),
	.L (L_1344),
	.V2C_1 (V2C_1344_192),
	.V2C_2 (V2C_1344_193),
	.V (V_1344)
);

VNU_2 #(quan_width) VNU1345 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_193_1345),
	.C2V_2 (C2V_194_1345),
	.L (L_1345),
	.V2C_1 (V2C_1345_193),
	.V2C_2 (V2C_1345_194),
	.V (V_1345)
);

VNU_2 #(quan_width) VNU1346 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_194_1346),
	.C2V_2 (C2V_195_1346),
	.L (L_1346),
	.V2C_1 (V2C_1346_194),
	.V2C_2 (V2C_1346_195),
	.V (V_1346)
);

VNU_2 #(quan_width) VNU1347 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_195_1347),
	.C2V_2 (C2V_196_1347),
	.L (L_1347),
	.V2C_1 (V2C_1347_195),
	.V2C_2 (V2C_1347_196),
	.V (V_1347)
);

VNU_2 #(quan_width) VNU1348 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_196_1348),
	.C2V_2 (C2V_197_1348),
	.L (L_1348),
	.V2C_1 (V2C_1348_196),
	.V2C_2 (V2C_1348_197),
	.V (V_1348)
);

VNU_2 #(quan_width) VNU1349 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_197_1349),
	.C2V_2 (C2V_198_1349),
	.L (L_1349),
	.V2C_1 (V2C_1349_197),
	.V2C_2 (V2C_1349_198),
	.V (V_1349)
);

VNU_2 #(quan_width) VNU1350 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_198_1350),
	.C2V_2 (C2V_199_1350),
	.L (L_1350),
	.V2C_1 (V2C_1350_198),
	.V2C_2 (V2C_1350_199),
	.V (V_1350)
);

VNU_2 #(quan_width) VNU1351 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_199_1351),
	.C2V_2 (C2V_200_1351),
	.L (L_1351),
	.V2C_1 (V2C_1351_199),
	.V2C_2 (V2C_1351_200),
	.V (V_1351)
);

VNU_2 #(quan_width) VNU1352 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_200_1352),
	.C2V_2 (C2V_201_1352),
	.L (L_1352),
	.V2C_1 (V2C_1352_200),
	.V2C_2 (V2C_1352_201),
	.V (V_1352)
);

VNU_2 #(quan_width) VNU1353 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_201_1353),
	.C2V_2 (C2V_202_1353),
	.L (L_1353),
	.V2C_1 (V2C_1353_201),
	.V2C_2 (V2C_1353_202),
	.V (V_1353)
);

VNU_2 #(quan_width) VNU1354 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_202_1354),
	.C2V_2 (C2V_203_1354),
	.L (L_1354),
	.V2C_1 (V2C_1354_202),
	.V2C_2 (V2C_1354_203),
	.V (V_1354)
);

VNU_2 #(quan_width) VNU1355 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_203_1355),
	.C2V_2 (C2V_204_1355),
	.L (L_1355),
	.V2C_1 (V2C_1355_203),
	.V2C_2 (V2C_1355_204),
	.V (V_1355)
);

VNU_2 #(quan_width) VNU1356 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_204_1356),
	.C2V_2 (C2V_205_1356),
	.L (L_1356),
	.V2C_1 (V2C_1356_204),
	.V2C_2 (V2C_1356_205),
	.V (V_1356)
);

VNU_2 #(quan_width) VNU1357 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_205_1357),
	.C2V_2 (C2V_206_1357),
	.L (L_1357),
	.V2C_1 (V2C_1357_205),
	.V2C_2 (V2C_1357_206),
	.V (V_1357)
);

VNU_2 #(quan_width) VNU1358 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_206_1358),
	.C2V_2 (C2V_207_1358),
	.L (L_1358),
	.V2C_1 (V2C_1358_206),
	.V2C_2 (V2C_1358_207),
	.V (V_1358)
);

VNU_2 #(quan_width) VNU1359 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_207_1359),
	.C2V_2 (C2V_208_1359),
	.L (L_1359),
	.V2C_1 (V2C_1359_207),
	.V2C_2 (V2C_1359_208),
	.V (V_1359)
);

VNU_2 #(quan_width) VNU1360 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_208_1360),
	.C2V_2 (C2V_209_1360),
	.L (L_1360),
	.V2C_1 (V2C_1360_208),
	.V2C_2 (V2C_1360_209),
	.V (V_1360)
);

VNU_2 #(quan_width) VNU1361 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_209_1361),
	.C2V_2 (C2V_210_1361),
	.L (L_1361),
	.V2C_1 (V2C_1361_209),
	.V2C_2 (V2C_1361_210),
	.V (V_1361)
);

VNU_2 #(quan_width) VNU1362 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_210_1362),
	.C2V_2 (C2V_211_1362),
	.L (L_1362),
	.V2C_1 (V2C_1362_210),
	.V2C_2 (V2C_1362_211),
	.V (V_1362)
);

VNU_2 #(quan_width) VNU1363 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_211_1363),
	.C2V_2 (C2V_212_1363),
	.L (L_1363),
	.V2C_1 (V2C_1363_211),
	.V2C_2 (V2C_1363_212),
	.V (V_1363)
);

VNU_2 #(quan_width) VNU1364 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_212_1364),
	.C2V_2 (C2V_213_1364),
	.L (L_1364),
	.V2C_1 (V2C_1364_212),
	.V2C_2 (V2C_1364_213),
	.V (V_1364)
);

VNU_2 #(quan_width) VNU1365 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_213_1365),
	.C2V_2 (C2V_214_1365),
	.L (L_1365),
	.V2C_1 (V2C_1365_213),
	.V2C_2 (V2C_1365_214),
	.V (V_1365)
);

VNU_2 #(quan_width) VNU1366 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_214_1366),
	.C2V_2 (C2V_215_1366),
	.L (L_1366),
	.V2C_1 (V2C_1366_214),
	.V2C_2 (V2C_1366_215),
	.V (V_1366)
);

VNU_2 #(quan_width) VNU1367 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_215_1367),
	.C2V_2 (C2V_216_1367),
	.L (L_1367),
	.V2C_1 (V2C_1367_215),
	.V2C_2 (V2C_1367_216),
	.V (V_1367)
);

VNU_2 #(quan_width) VNU1368 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_216_1368),
	.C2V_2 (C2V_217_1368),
	.L (L_1368),
	.V2C_1 (V2C_1368_216),
	.V2C_2 (V2C_1368_217),
	.V (V_1368)
);

VNU_2 #(quan_width) VNU1369 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_217_1369),
	.C2V_2 (C2V_218_1369),
	.L (L_1369),
	.V2C_1 (V2C_1369_217),
	.V2C_2 (V2C_1369_218),
	.V (V_1369)
);

VNU_2 #(quan_width) VNU1370 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_218_1370),
	.C2V_2 (C2V_219_1370),
	.L (L_1370),
	.V2C_1 (V2C_1370_218),
	.V2C_2 (V2C_1370_219),
	.V (V_1370)
);

VNU_2 #(quan_width) VNU1371 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_219_1371),
	.C2V_2 (C2V_220_1371),
	.L (L_1371),
	.V2C_1 (V2C_1371_219),
	.V2C_2 (V2C_1371_220),
	.V (V_1371)
);

VNU_2 #(quan_width) VNU1372 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_220_1372),
	.C2V_2 (C2V_221_1372),
	.L (L_1372),
	.V2C_1 (V2C_1372_220),
	.V2C_2 (V2C_1372_221),
	.V (V_1372)
);

VNU_2 #(quan_width) VNU1373 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_221_1373),
	.C2V_2 (C2V_222_1373),
	.L (L_1373),
	.V2C_1 (V2C_1373_221),
	.V2C_2 (V2C_1373_222),
	.V (V_1373)
);

VNU_2 #(quan_width) VNU1374 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_222_1374),
	.C2V_2 (C2V_223_1374),
	.L (L_1374),
	.V2C_1 (V2C_1374_222),
	.V2C_2 (V2C_1374_223),
	.V (V_1374)
);

VNU_2 #(quan_width) VNU1375 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_223_1375),
	.C2V_2 (C2V_224_1375),
	.L (L_1375),
	.V2C_1 (V2C_1375_223),
	.V2C_2 (V2C_1375_224),
	.V (V_1375)
);

VNU_2 #(quan_width) VNU1376 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_224_1376),
	.C2V_2 (C2V_225_1376),
	.L (L_1376),
	.V2C_1 (V2C_1376_224),
	.V2C_2 (V2C_1376_225),
	.V (V_1376)
);

VNU_2 #(quan_width) VNU1377 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_225_1377),
	.C2V_2 (C2V_226_1377),
	.L (L_1377),
	.V2C_1 (V2C_1377_225),
	.V2C_2 (V2C_1377_226),
	.V (V_1377)
);

VNU_2 #(quan_width) VNU1378 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_226_1378),
	.C2V_2 (C2V_227_1378),
	.L (L_1378),
	.V2C_1 (V2C_1378_226),
	.V2C_2 (V2C_1378_227),
	.V (V_1378)
);

VNU_2 #(quan_width) VNU1379 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_227_1379),
	.C2V_2 (C2V_228_1379),
	.L (L_1379),
	.V2C_1 (V2C_1379_227),
	.V2C_2 (V2C_1379_228),
	.V (V_1379)
);

VNU_2 #(quan_width) VNU1380 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_228_1380),
	.C2V_2 (C2V_229_1380),
	.L (L_1380),
	.V2C_1 (V2C_1380_228),
	.V2C_2 (V2C_1380_229),
	.V (V_1380)
);

VNU_2 #(quan_width) VNU1381 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_229_1381),
	.C2V_2 (C2V_230_1381),
	.L (L_1381),
	.V2C_1 (V2C_1381_229),
	.V2C_2 (V2C_1381_230),
	.V (V_1381)
);

VNU_2 #(quan_width) VNU1382 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_230_1382),
	.C2V_2 (C2V_231_1382),
	.L (L_1382),
	.V2C_1 (V2C_1382_230),
	.V2C_2 (V2C_1382_231),
	.V (V_1382)
);

VNU_2 #(quan_width) VNU1383 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_231_1383),
	.C2V_2 (C2V_232_1383),
	.L (L_1383),
	.V2C_1 (V2C_1383_231),
	.V2C_2 (V2C_1383_232),
	.V (V_1383)
);

VNU_2 #(quan_width) VNU1384 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_232_1384),
	.C2V_2 (C2V_233_1384),
	.L (L_1384),
	.V2C_1 (V2C_1384_232),
	.V2C_2 (V2C_1384_233),
	.V (V_1384)
);

VNU_2 #(quan_width) VNU1385 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_233_1385),
	.C2V_2 (C2V_234_1385),
	.L (L_1385),
	.V2C_1 (V2C_1385_233),
	.V2C_2 (V2C_1385_234),
	.V (V_1385)
);

VNU_2 #(quan_width) VNU1386 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_234_1386),
	.C2V_2 (C2V_235_1386),
	.L (L_1386),
	.V2C_1 (V2C_1386_234),
	.V2C_2 (V2C_1386_235),
	.V (V_1386)
);

VNU_2 #(quan_width) VNU1387 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_235_1387),
	.C2V_2 (C2V_236_1387),
	.L (L_1387),
	.V2C_1 (V2C_1387_235),
	.V2C_2 (V2C_1387_236),
	.V (V_1387)
);

VNU_2 #(quan_width) VNU1388 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_236_1388),
	.C2V_2 (C2V_237_1388),
	.L (L_1388),
	.V2C_1 (V2C_1388_236),
	.V2C_2 (V2C_1388_237),
	.V (V_1388)
);

VNU_2 #(quan_width) VNU1389 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_237_1389),
	.C2V_2 (C2V_238_1389),
	.L (L_1389),
	.V2C_1 (V2C_1389_237),
	.V2C_2 (V2C_1389_238),
	.V (V_1389)
);

VNU_2 #(quan_width) VNU1390 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_238_1390),
	.C2V_2 (C2V_239_1390),
	.L (L_1390),
	.V2C_1 (V2C_1390_238),
	.V2C_2 (V2C_1390_239),
	.V (V_1390)
);

VNU_2 #(quan_width) VNU1391 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_239_1391),
	.C2V_2 (C2V_240_1391),
	.L (L_1391),
	.V2C_1 (V2C_1391_239),
	.V2C_2 (V2C_1391_240),
	.V (V_1391)
);

VNU_2 #(quan_width) VNU1392 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_240_1392),
	.C2V_2 (C2V_241_1392),
	.L (L_1392),
	.V2C_1 (V2C_1392_240),
	.V2C_2 (V2C_1392_241),
	.V (V_1392)
);

VNU_2 #(quan_width) VNU1393 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_241_1393),
	.C2V_2 (C2V_242_1393),
	.L (L_1393),
	.V2C_1 (V2C_1393_241),
	.V2C_2 (V2C_1393_242),
	.V (V_1393)
);

VNU_2 #(quan_width) VNU1394 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_242_1394),
	.C2V_2 (C2V_243_1394),
	.L (L_1394),
	.V2C_1 (V2C_1394_242),
	.V2C_2 (V2C_1394_243),
	.V (V_1394)
);

VNU_2 #(quan_width) VNU1395 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_243_1395),
	.C2V_2 (C2V_244_1395),
	.L (L_1395),
	.V2C_1 (V2C_1395_243),
	.V2C_2 (V2C_1395_244),
	.V (V_1395)
);

VNU_2 #(quan_width) VNU1396 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_244_1396),
	.C2V_2 (C2V_245_1396),
	.L (L_1396),
	.V2C_1 (V2C_1396_244),
	.V2C_2 (V2C_1396_245),
	.V (V_1396)
);

VNU_2 #(quan_width) VNU1397 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_245_1397),
	.C2V_2 (C2V_246_1397),
	.L (L_1397),
	.V2C_1 (V2C_1397_245),
	.V2C_2 (V2C_1397_246),
	.V (V_1397)
);

VNU_2 #(quan_width) VNU1398 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_246_1398),
	.C2V_2 (C2V_247_1398),
	.L (L_1398),
	.V2C_1 (V2C_1398_246),
	.V2C_2 (V2C_1398_247),
	.V (V_1398)
);

VNU_2 #(quan_width) VNU1399 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_247_1399),
	.C2V_2 (C2V_248_1399),
	.L (L_1399),
	.V2C_1 (V2C_1399_247),
	.V2C_2 (V2C_1399_248),
	.V (V_1399)
);

VNU_2 #(quan_width) VNU1400 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_248_1400),
	.C2V_2 (C2V_249_1400),
	.L (L_1400),
	.V2C_1 (V2C_1400_248),
	.V2C_2 (V2C_1400_249),
	.V (V_1400)
);

VNU_2 #(quan_width) VNU1401 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_249_1401),
	.C2V_2 (C2V_250_1401),
	.L (L_1401),
	.V2C_1 (V2C_1401_249),
	.V2C_2 (V2C_1401_250),
	.V (V_1401)
);

VNU_2 #(quan_width) VNU1402 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_250_1402),
	.C2V_2 (C2V_251_1402),
	.L (L_1402),
	.V2C_1 (V2C_1402_250),
	.V2C_2 (V2C_1402_251),
	.V (V_1402)
);

VNU_2 #(quan_width) VNU1403 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_251_1403),
	.C2V_2 (C2V_252_1403),
	.L (L_1403),
	.V2C_1 (V2C_1403_251),
	.V2C_2 (V2C_1403_252),
	.V (V_1403)
);

VNU_2 #(quan_width) VNU1404 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_252_1404),
	.C2V_2 (C2V_253_1404),
	.L (L_1404),
	.V2C_1 (V2C_1404_252),
	.V2C_2 (V2C_1404_253),
	.V (V_1404)
);

VNU_2 #(quan_width) VNU1405 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_253_1405),
	.C2V_2 (C2V_254_1405),
	.L (L_1405),
	.V2C_1 (V2C_1405_253),
	.V2C_2 (V2C_1405_254),
	.V (V_1405)
);

VNU_2 #(quan_width) VNU1406 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_254_1406),
	.C2V_2 (C2V_255_1406),
	.L (L_1406),
	.V2C_1 (V2C_1406_254),
	.V2C_2 (V2C_1406_255),
	.V (V_1406)
);

VNU_2 #(quan_width) VNU1407 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_255_1407),
	.C2V_2 (C2V_256_1407),
	.L (L_1407),
	.V2C_1 (V2C_1407_255),
	.V2C_2 (V2C_1407_256),
	.V (V_1407)
);

VNU_2 #(quan_width) VNU1408 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_256_1408),
	.C2V_2 (C2V_257_1408),
	.L (L_1408),
	.V2C_1 (V2C_1408_256),
	.V2C_2 (V2C_1408_257),
	.V (V_1408)
);

VNU_2 #(quan_width) VNU1409 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_257_1409),
	.C2V_2 (C2V_258_1409),
	.L (L_1409),
	.V2C_1 (V2C_1409_257),
	.V2C_2 (V2C_1409_258),
	.V (V_1409)
);

VNU_2 #(quan_width) VNU1410 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_258_1410),
	.C2V_2 (C2V_259_1410),
	.L (L_1410),
	.V2C_1 (V2C_1410_258),
	.V2C_2 (V2C_1410_259),
	.V (V_1410)
);

VNU_2 #(quan_width) VNU1411 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_259_1411),
	.C2V_2 (C2V_260_1411),
	.L (L_1411),
	.V2C_1 (V2C_1411_259),
	.V2C_2 (V2C_1411_260),
	.V (V_1411)
);

VNU_2 #(quan_width) VNU1412 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_260_1412),
	.C2V_2 (C2V_261_1412),
	.L (L_1412),
	.V2C_1 (V2C_1412_260),
	.V2C_2 (V2C_1412_261),
	.V (V_1412)
);

VNU_2 #(quan_width) VNU1413 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_261_1413),
	.C2V_2 (C2V_262_1413),
	.L (L_1413),
	.V2C_1 (V2C_1413_261),
	.V2C_2 (V2C_1413_262),
	.V (V_1413)
);

VNU_2 #(quan_width) VNU1414 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_262_1414),
	.C2V_2 (C2V_263_1414),
	.L (L_1414),
	.V2C_1 (V2C_1414_262),
	.V2C_2 (V2C_1414_263),
	.V (V_1414)
);

VNU_2 #(quan_width) VNU1415 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_263_1415),
	.C2V_2 (C2V_264_1415),
	.L (L_1415),
	.V2C_1 (V2C_1415_263),
	.V2C_2 (V2C_1415_264),
	.V (V_1415)
);

VNU_2 #(quan_width) VNU1416 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_264_1416),
	.C2V_2 (C2V_265_1416),
	.L (L_1416),
	.V2C_1 (V2C_1416_264),
	.V2C_2 (V2C_1416_265),
	.V (V_1416)
);

VNU_2 #(quan_width) VNU1417 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_265_1417),
	.C2V_2 (C2V_266_1417),
	.L (L_1417),
	.V2C_1 (V2C_1417_265),
	.V2C_2 (V2C_1417_266),
	.V (V_1417)
);

VNU_2 #(quan_width) VNU1418 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_266_1418),
	.C2V_2 (C2V_267_1418),
	.L (L_1418),
	.V2C_1 (V2C_1418_266),
	.V2C_2 (V2C_1418_267),
	.V (V_1418)
);

VNU_2 #(quan_width) VNU1419 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_267_1419),
	.C2V_2 (C2V_268_1419),
	.L (L_1419),
	.V2C_1 (V2C_1419_267),
	.V2C_2 (V2C_1419_268),
	.V (V_1419)
);

VNU_2 #(quan_width) VNU1420 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_268_1420),
	.C2V_2 (C2V_269_1420),
	.L (L_1420),
	.V2C_1 (V2C_1420_268),
	.V2C_2 (V2C_1420_269),
	.V (V_1420)
);

VNU_2 #(quan_width) VNU1421 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_269_1421),
	.C2V_2 (C2V_270_1421),
	.L (L_1421),
	.V2C_1 (V2C_1421_269),
	.V2C_2 (V2C_1421_270),
	.V (V_1421)
);

VNU_2 #(quan_width) VNU1422 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_270_1422),
	.C2V_2 (C2V_271_1422),
	.L (L_1422),
	.V2C_1 (V2C_1422_270),
	.V2C_2 (V2C_1422_271),
	.V (V_1422)
);

VNU_2 #(quan_width) VNU1423 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_271_1423),
	.C2V_2 (C2V_272_1423),
	.L (L_1423),
	.V2C_1 (V2C_1423_271),
	.V2C_2 (V2C_1423_272),
	.V (V_1423)
);

VNU_2 #(quan_width) VNU1424 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_272_1424),
	.C2V_2 (C2V_273_1424),
	.L (L_1424),
	.V2C_1 (V2C_1424_272),
	.V2C_2 (V2C_1424_273),
	.V (V_1424)
);

VNU_2 #(quan_width) VNU1425 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_273_1425),
	.C2V_2 (C2V_274_1425),
	.L (L_1425),
	.V2C_1 (V2C_1425_273),
	.V2C_2 (V2C_1425_274),
	.V (V_1425)
);

VNU_2 #(quan_width) VNU1426 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_274_1426),
	.C2V_2 (C2V_275_1426),
	.L (L_1426),
	.V2C_1 (V2C_1426_274),
	.V2C_2 (V2C_1426_275),
	.V (V_1426)
);

VNU_2 #(quan_width) VNU1427 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_275_1427),
	.C2V_2 (C2V_276_1427),
	.L (L_1427),
	.V2C_1 (V2C_1427_275),
	.V2C_2 (V2C_1427_276),
	.V (V_1427)
);

VNU_2 #(quan_width) VNU1428 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_276_1428),
	.C2V_2 (C2V_277_1428),
	.L (L_1428),
	.V2C_1 (V2C_1428_276),
	.V2C_2 (V2C_1428_277),
	.V (V_1428)
);

VNU_2 #(quan_width) VNU1429 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_277_1429),
	.C2V_2 (C2V_278_1429),
	.L (L_1429),
	.V2C_1 (V2C_1429_277),
	.V2C_2 (V2C_1429_278),
	.V (V_1429)
);

VNU_2 #(quan_width) VNU1430 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_278_1430),
	.C2V_2 (C2V_279_1430),
	.L (L_1430),
	.V2C_1 (V2C_1430_278),
	.V2C_2 (V2C_1430_279),
	.V (V_1430)
);

VNU_2 #(quan_width) VNU1431 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_279_1431),
	.C2V_2 (C2V_280_1431),
	.L (L_1431),
	.V2C_1 (V2C_1431_279),
	.V2C_2 (V2C_1431_280),
	.V (V_1431)
);

VNU_2 #(quan_width) VNU1432 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_280_1432),
	.C2V_2 (C2V_281_1432),
	.L (L_1432),
	.V2C_1 (V2C_1432_280),
	.V2C_2 (V2C_1432_281),
	.V (V_1432)
);

VNU_2 #(quan_width) VNU1433 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_281_1433),
	.C2V_2 (C2V_282_1433),
	.L (L_1433),
	.V2C_1 (V2C_1433_281),
	.V2C_2 (V2C_1433_282),
	.V (V_1433)
);

VNU_2 #(quan_width) VNU1434 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_282_1434),
	.C2V_2 (C2V_283_1434),
	.L (L_1434),
	.V2C_1 (V2C_1434_282),
	.V2C_2 (V2C_1434_283),
	.V (V_1434)
);

VNU_2 #(quan_width) VNU1435 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_283_1435),
	.C2V_2 (C2V_284_1435),
	.L (L_1435),
	.V2C_1 (V2C_1435_283),
	.V2C_2 (V2C_1435_284),
	.V (V_1435)
);

VNU_2 #(quan_width) VNU1436 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_284_1436),
	.C2V_2 (C2V_285_1436),
	.L (L_1436),
	.V2C_1 (V2C_1436_284),
	.V2C_2 (V2C_1436_285),
	.V (V_1436)
);

VNU_2 #(quan_width) VNU1437 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_285_1437),
	.C2V_2 (C2V_286_1437),
	.L (L_1437),
	.V2C_1 (V2C_1437_285),
	.V2C_2 (V2C_1437_286),
	.V (V_1437)
);

VNU_2 #(quan_width) VNU1438 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_286_1438),
	.C2V_2 (C2V_287_1438),
	.L (L_1438),
	.V2C_1 (V2C_1438_286),
	.V2C_2 (V2C_1438_287),
	.V (V_1438)
);

VNU_2 #(quan_width) VNU1439 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_287_1439),
	.C2V_2 (C2V_288_1439),
	.L (L_1439),
	.V2C_1 (V2C_1439_287),
	.V2C_2 (V2C_1439_288),
	.V (V_1439)
);

VNU_1 #(quan_width) VNU1440 (
	.clk (clk),
	.rst (rst),
	.cnt (cnt),
	.init_cnt (8'd11),
	.C2V_1 (C2V_288_1440),
	.L (L_1440),
	.V2C_1 (V2C_1440_288),
	.V (V_1440)
);

endmodule